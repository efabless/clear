* NGSPICE file created from top_left_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

.subckt top_left_tile VGND VPWR ccff_head ccff_head_0 ccff_tail ccff_tail_0 chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[20] chanx_right_in[21] chanx_right_in[22] chanx_right_in[23]
+ chanx_right_in[24] chanx_right_in[25] chanx_right_in[26] chanx_right_in[27] chanx_right_in[28]
+ chanx_right_in[29] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[20] chanx_right_out[21]
+ chanx_right_out[22] chanx_right_out[23] chanx_right_out[24] chanx_right_out[25]
+ chanx_right_out[26] chanx_right_out[27] chanx_right_out[28] chanx_right_out[29]
+ chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6]
+ chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_bottom_in_0[0] chany_bottom_in_0[10]
+ chany_bottom_in_0[11] chany_bottom_in_0[12] chany_bottom_in_0[13] chany_bottom_in_0[14]
+ chany_bottom_in_0[15] chany_bottom_in_0[16] chany_bottom_in_0[17] chany_bottom_in_0[18]
+ chany_bottom_in_0[19] chany_bottom_in_0[1] chany_bottom_in_0[20] chany_bottom_in_0[21]
+ chany_bottom_in_0[22] chany_bottom_in_0[23] chany_bottom_in_0[24] chany_bottom_in_0[25]
+ chany_bottom_in_0[26] chany_bottom_in_0[27] chany_bottom_in_0[28] chany_bottom_in_0[29]
+ chany_bottom_in_0[2] chany_bottom_in_0[3] chany_bottom_in_0[4] chany_bottom_in_0[5]
+ chany_bottom_in_0[6] chany_bottom_in_0[7] chany_bottom_in_0[8] chany_bottom_in_0[9]
+ chany_bottom_out_0[0] chany_bottom_out_0[10] chany_bottom_out_0[11] chany_bottom_out_0[12]
+ chany_bottom_out_0[13] chany_bottom_out_0[14] chany_bottom_out_0[15] chany_bottom_out_0[16]
+ chany_bottom_out_0[17] chany_bottom_out_0[18] chany_bottom_out_0[19] chany_bottom_out_0[1]
+ chany_bottom_out_0[20] chany_bottom_out_0[21] chany_bottom_out_0[22] chany_bottom_out_0[23]
+ chany_bottom_out_0[24] chany_bottom_out_0[25] chany_bottom_out_0[26] chany_bottom_out_0[27]
+ chany_bottom_out_0[28] chany_bottom_out_0[29] chany_bottom_out_0[2] chany_bottom_out_0[3]
+ chany_bottom_out_0[4] chany_bottom_out_0[5] chany_bottom_out_0[6] chany_bottom_out_0[7]
+ chany_bottom_out_0[8] chany_bottom_out_0[9] gfpga_pad_io_soc_dir[0] gfpga_pad_io_soc_dir[1]
+ gfpga_pad_io_soc_dir[2] gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0] gfpga_pad_io_soc_in[1]
+ gfpga_pad_io_soc_in[2] gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0] gfpga_pad_io_soc_out[1]
+ gfpga_pad_io_soc_out[2] gfpga_pad_io_soc_out[3] isol_n prog_clk prog_reset reset
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
+ right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_ right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_ right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ right_width_0_height_0_subtile_0__pin_inpad_0_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ right_width_0_height_0_subtile_2__pin_inpad_0_ right_width_0_height_0_subtile_3__pin_inpad_0_
+ test_enable
XFILLER_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold3_A prog_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0 sb_0__8_.mux_bottom_track_31.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_6.mux_l1_in_0_ net80 net77 sb_0__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_ net58 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__S sb_0__8_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_131_ sb_0__8_.mux_right_track_4.out VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input55_A chany_bottom_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_58.mux_l1_in_0_ net76 net72 sb_0__8_.mem_right_track_58.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_0_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__8_.mem_bottom_track_31.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_33.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_10_0_prog_clk cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
+ net204 VGND VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_ net7 net41 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_14.mux_l1_in_1__167 VGND VGND VPWR VPWR net167 sb_0__8_.mux_right_track_14.mux_l1_in_1__167/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_114_ sb_0__8_.mux_right_track_38.out VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input18_A chanx_right_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_44.mux_l1_in_1__184 VGND VGND VPWR VPWR net184 sb_0__8_.mux_right_track_44.mux_l1_in_1__184/LO
+ sky130_fd_sc_hd__conb_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__8_.mem_right_track_32.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_34.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A0 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput97 net97 VGND VGND VPWR VPWR chanx_right_out[22] sky130_fd_sc_hd__buf_12
XANTENNA_output124_A net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput86 net86 VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A1 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_ cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_6_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_130_ sb_0__8_.mux_right_track_6.out VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_0__A0 right_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input48_A chany_bottom_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__135__A net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_ sb_0__8_.mux_bottom_track_13.out
+ net48 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_bottom_track_47.mux_l1_in_0__A0 right_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_113_ sb_0__8_.mux_right_track_40.out VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_right_track_16.mux_l2_in_0_ sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_16.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A0 sb_0__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_2_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput98 net98 VGND VGND VPWR VPWR chanx_right_out[23] sky130_fd_sc_hd__buf_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput87 net87 VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_12
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input30_A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__143__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_16.mux_l1_in_1_ net168 net62 sb_0__8_.mem_right_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input78_A right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_right_track_56.mux_l1_in_0__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__8_.mem_bottom_track_51.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfrtp_2
XFILLER_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_4.mux_l2_in_1__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_8_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__151__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_ sb_0__8_.mux_bottom_track_7.out
+ net51 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__8_.mem_right_track_52.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_52.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_70_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_112_ sb_0__8_.mux_right_track_42.out VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input60_A chany_bottom_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_bottom_track_13.mux_l1_in_0__A0 right_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold10 ccff_head_0 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__8_.mem_right_track_0.mem_out\[1\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_43_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_bottom_track_31.mux_l2_in_0__154 VGND VGND VPWR VPWR net154 sb_0__8_.mux_bottom_track_31.mux_l2_in_0__154/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_20.out sky130_fd_sc_hd__clkbuf_1
Xoutput99 net99 VGND VGND VPWR VPWR chanx_right_out[24] sky130_fd_sc_hd__buf_12
XFILLER_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput88 net88 VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_12
XANTENNA_input23_A chanx_right_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_16.mux_l1_in_0_ net75 net79 sb_0__8_.mem_right_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__D cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_28.mux_l2_in_0_ sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__8_.mem_bottom_track_49.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_51.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__8_.mux_right_track_30.mux_l2_in_0_ sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_30.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA__154__A sb_0__8_.mux_bottom_track_19.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_14.out sky130_fd_sc_hd__clkbuf_1
XFILLER_27_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_92_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_22.mux_l1_in_0__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__149__A sb_0__8_.mux_bottom_track_29.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_13.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_1__S sb_0__8_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_28.mux_l1_in_1_ net175 net39 sb_0__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_4_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk sb_0__8_.mem_right_track_20.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_13.mux_l2_in_0_ net200 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_13.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mux_right_track_30.mux_l1_in_1_ net176 net40 sb_0__8_.mem_right_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_2_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ sb_0__8_.mux_bottom_track_1.out
+ net54 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__8_.mem_right_track_50.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_111_ sb_0__8_.mux_right_track_44.out VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input53_A chany_bottom_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 net208 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__8_.mem_right_track_0.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_43_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__157__A sb_0__8_.mux_bottom_track_13.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_10.mux_l2_in_1__165 VGND VGND VPWR VPWR net165 sb_0__8_.mux_right_track_10.mux_l2_in_1__165/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__195 VGND VGND VPWR VPWR net195
+ cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__195/LO sky130_fd_sc_hd__conb_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput89 net89 VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_12
XANTENNA_input16_A chanx_right_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__8_.mem_right_track_58.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input8_A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_30.mux_l1_in_1__176 VGND VGND VPWR VPWR net176 sb_0__8_.mux_right_track_30.mux_l1_in_1__176/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_45_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output122_A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_42.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_42.out sky130_fd_sc_hd__clkbuf_1
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_3_0_prog_clk sb_0__8_.mem_right_track_6.mem_out\[1\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_28.mux_l1_in_0_ net73 net77 sb_0__8_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_0__8_.mem_right_track_18.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mux_right_track_2.mux_l3_in_0_ sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sb_0__8_.mem_right_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_36.out sky130_fd_sc_hd__clkbuf_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_30.mux_l1_in_0_ net74 net78 sb_0__8_.mem_right_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_42.mux_l2_in_0_ net183 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_42.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_35.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_5_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_110_ sb_0__8_.mux_right_track_46.out VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_bottom_track_5.mux_l2_in_0_ net160 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_5.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A0 net13 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input46_A chany_bottom_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_2.mux_l2_in_1_ net170 net55 sb_0__8_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_52_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_13.mux_l1_in_0_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ net30 sb_0__8_.mem_bottom_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold12 ccff_head VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net211
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ net209 net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk sb_0__8_.mem_right_track_26.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_26.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_56.mux_l2_in_0__190 VGND VGND VPWR VPWR net190 sb_0__8_.mux_right_track_56.mux_l2_in_0__190/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_3.out sky130_fd_sc_hd__clkbuf_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_0__8_.mem_right_track_56.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_58.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0__S cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_95_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_1__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_0__8_.mem_right_track_6.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input76_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_2.ccff_tail net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_45.mux_l2_in_0__157 VGND VGND VPWR VPWR net157 sb_0__8_.mux_bottom_track_45.mux_l2_in_0__157/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_58.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_58.out sky130_fd_sc_hd__clkbuf_1
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input39_A chany_bottom_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_169_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
Xsb_0__8_.mux_right_track_26.mux_l2_in_0__174 VGND VGND VPWR VPWR net174 sb_0__8_.mux_right_track_26.mux_l2_in_0__174/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_2.mux_l2_in_0_ sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_37_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__S cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold13 net210 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_0__8_.mem_right_track_24.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_26.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__8_.mux_right_track_42.mux_l1_in_0_ net47 net72 sb_0__8_.mem_right_track_42.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_54.mux_l2_in_0_ net189 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_54.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1 sb_0__8_.mux_bottom_track_49.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_bottom_track_5.mux_l1_in_0_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ net26 sb_0__8_.mem_bottom_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mux_right_track_2.mux_l1_in_1_ net75 net72 sb_0__8_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_6.mux_l2_in_1__192 VGND VGND VPWR VPWR net192 sb_0__8_.mux_right_track_6.mux_l2_in_1__192/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input21_A chanx_right_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_13_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__8_.mem_right_track_4.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input69_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__8_.mem_bottom_track_3.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_12.mux_l1_in_1__166 VGND VGND VPWR VPWR net166 sb_0__8_.mux_right_track_12.mux_l1_in_1__166/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__D sb_0__8_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_ net195 sb_0__8_.mux_bottom_track_51.out
+ cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_168_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_1__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input51_A chany_bottom_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_ net15 net34 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mux_right_track_2.mux_l1_in_0_ net69 net78 sb_0__8_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cby_0__8_.cby_0__1_.mem_right_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input14_A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_54.mux_l1_in_0_ net53 net70 sb_0__8_.mem_right_track_54.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_94_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_ cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A0 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__8_.mem_bottom_track_1.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__8_.mux_right_track_38.mux_l2_in_0__180 VGND VGND VPWR VPWR net180 sb_0__8_.mux_right_track_38.mux_l2_in_0__180/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net65 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__8_.mem_right_track_44.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_49.mux_l2_in_0_ net159 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_49.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_51.mux_l2_in_0_ net161 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ net81 VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_ net57 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_167_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__D cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1__S cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_bottom_track_19.mux_l1_in_0__A0 right_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__8_.mem_bottom_track_9.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_input44_A chany_bottom_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_4_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__8_.mem_bottom_track_11.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_ net8 net40 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_0__8_.mem_right_track_12.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output113_A net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_12.mux_l2_in_0_ sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__8_.mem_bottom_track_49.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_49.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__8_.mem_right_track_42.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input74_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net82 net67 VGND VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_ cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0 sb_0__8_.mux_bottom_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_166_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_12.mux_l1_in_1_ net166 net60 sb_0__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_49.mux_l1_in_0_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ net20 sb_0__8_.mem_bottom_track_49.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__8_.mem_bottom_track_7.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input37_A chany_bottom_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_149_ sb_0__8_.mux_bottom_track_29.out VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
Xsb_0__8_.mux_bottom_track_51.mux_l1_in_0_ right_width_0_height_0_subtile_3__pin_inpad_0_
+ net21 sb_0__8_.mem_bottom_track_51.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__8_.mem_bottom_track_11.ccff_head
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_ sb_0__8_.mux_bottom_track_15.out
+ net47 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A0 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_36.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_42.mux_l2_in_0__183 VGND VGND VPWR VPWR net183 sb_0__8_.mux_right_track_42.mux_l2_in_0__183/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__8_.mem_bottom_track_17.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_17.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_0__8_.mem_right_track_10.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_91_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_bottom_track_35.mux_l1_in_0__A0 right_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__8_.mem_bottom_track_47.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_49.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input67_A isol_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A0 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A1 net50 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__S cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_165_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__8_.mem_right_track_18.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_18.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_92_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_12.mux_l1_in_0_ net73 net77 sb_0__8_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mux_bottom_track_17.mux_l2_in_0__202 VGND VGND VPWR VPWR net202 sb_0__8_.mux_bottom_track_17.mux_l2_in_0__202/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail net67 VGND
+ VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A0 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_24.mux_l2_in_0_ net173 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_24.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_148_ sb_0__8_.mux_bottom_track_31.out VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_ sb_0__8_.mux_bottom_track_9.out
+ net50 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__8_.mux_bottom_track_3.mux_l1_in_0__A0 right_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_0_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_10_0_prog_clk cby_0__8_.cby_0__1_.ccff_tail net204 VGND VGND VPWR VPWR
+ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__8_.mem_bottom_track_15.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_17.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__S cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_bottom_track_3.mux_l2_in_0__153 VGND VGND VPWR VPWR net153 sb_0__8_.mux_bottom_track_3.mux_l2_in_0__153/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_91_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input12_A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input4_A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_164_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_0__8_.mem_right_track_16.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_18.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_92_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_5_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_147_ sb_0__8_.mux_bottom_track_33.out VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_ sb_0__8_.mux_bottom_track_3.out
+ net53 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_32.out sky130_fd_sc_hd__clkbuf_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__8_.mem_right_track_30.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_30.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A0 right_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input42_A chany_bottom_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_1__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_31.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_24.mux_l1_in_0_ net37 net71 sb_0__8_.mem_right_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_3_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__8_.mux_right_track_36.mux_l2_in_0_ net179 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_36.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_26.out sky130_fd_sc_hd__clkbuf_1
XFILLER_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0 sb_0__8_.mux_bottom_track_19.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_bottom_track_1.mux_l2_in_0_ sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_19.mux_l2_in_0_ net151 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_19.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0 net15 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output111_A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_19.out sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_1.mux_l1_in_1_ net198 right_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_0__8_.mem_bottom_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input72_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_163_ sb_0__8_.mux_bottom_track_1.out VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_24.mux_l2_in_0__173 VGND VGND VPWR VPWR net173 sb_0__8_.mux_right_track_24.mux_l2_in_0__173/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_146_ sb_0__8_.mux_bottom_track_35.out VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1__D sb_0__8_.mem_right_track_58.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__8_.mem_bottom_track_35.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_35.ccff_tail sky130_fd_sc_hd__dfrtp_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__8_.mem_right_track_28.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_30.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input35_A chany_bottom_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_129_ sb_0__8_.mux_right_track_8.out VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput80 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND
+ VPWR VPWR net80 sky130_fd_sc_hd__buf_2
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_54.out sky130_fd_sc_hd__clkbuf_1
XFILLER_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_11.mux_l2_in_0__199 VGND VGND VPWR VPWR net199 sb_0__8_.mux_bottom_track_11.mux_l2_in_0__199/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__8_.mux_right_track_8.mux_l3_in_0_ sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X sb_0__8_.mem_right_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk sb_0__8_.mem_right_track_36.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_48.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__8_.mux_right_track_36.mux_l1_in_0_ net43 net69 sb_0__8_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_73_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1 net34 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_48.mux_l2_in_0_ sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_48.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_57_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_47.out sky130_fd_sc_hd__clkbuf_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__S sb_0__8_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_50.mux_l2_in_0_ net187 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_50.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mux_bottom_track_1.mux_l1_in_0_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ net14 sb_0__8_.mem_bottom_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_1__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_162_ sb_0__8_.mux_bottom_track_3.out VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_8.mux_l2_in_1_ net193 net58 sb_0__8_.mem_right_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_input65_A gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_bottom_track_19.mux_l1_in_0_ right_width_0_height_0_subtile_3__pin_inpad_0_
+ net4 sb_0__8_.mem_bottom_track_19.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 net215 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_48.mux_l1_in_1_ net186 net50 sb_0__8_.mem_right_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A0 sb_0__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_bottom_track_33.mux_l2_in_0_ net155 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_33.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_145_ net13 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__8_.mem_bottom_track_33.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_35.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_4.mux_l2_in_1__181 VGND VGND VPWR VPWR net181 sb_0__8_.mux_right_track_4.mux_l2_in_1__181/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input28_A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_128_ sb_0__8_.mux_right_track_10.out VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput70 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND VGND VPWR
+ VPWR net70 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_9.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_0__8_.mem_right_track_34.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_14_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input10_A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_8.mux_l2_in_0_ sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_161_ sb_0__8_.mux_bottom_track_5.out VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input58_A chany_bottom_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__136__A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 net213 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
Xsb_0__8_.mux_right_track_48.mux_l1_in_0_ net75 net79 sb_0__8_.mem_right_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_144_ net15 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_50.mux_l1_in_0_ net51 net80 sb_0__8_.mem_right_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_65_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_8.mux_l1_in_1_ net75 net72 sb_0__8_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_ net196 net22 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_127_ sb_0__8_.mux_right_track_12.out VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput71 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND VGND VPWR
+ VPWR net71 sky130_fd_sc_hd__clkbuf_4
Xinput60 chany_bottom_in_0[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_33.mux_l1_in_0_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ net11 sb_0__8_.mem_bottom_track_33.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input40_A chany_bottom_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_bottom_track_45.mux_l2_in_0_ net157 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_45.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__144__A net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_ net16 net62 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_2_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_0__8_.cby_0__1_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__139__A sb_0__8_.mux_bottom_track_49.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_2_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A0 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_ cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
X_160_ sb_0__8_.mux_bottom_track_7.out VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__152__A net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput3 chanx_right_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input70_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_143_ net16 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_ net56 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_8.mux_l1_in_0_ net69 net78 sb_0__8_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_2_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_15_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_126_ sb_0__8_.mux_right_track_14.out VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__8_.mem_right_track_54.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_54.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput72 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND VGND VPWR
+ VPWR net72 sky130_fd_sc_hd__buf_2
Xinput61 chany_bottom_in_0[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput50 chany_bottom_in_0[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_44_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mux_bottom_track_9.mux_l1_in_0__A0 right_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input33_A chany_bottom_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_40.mux_l2_in_0__182 VGND VGND VPWR VPWR net182 sb_0__8_.mux_right_track_40.mux_l2_in_0__182/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_ sb_0__8_.mux_bottom_track_29.out
+ net39 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_2_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__160__A sb_0__8_.mux_bottom_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_109_ sb_0__8_.mux_right_track_48.out VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__8_.mem_right_track_2.mem_out\[1\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_bottom_track_49.mux_l1_in_0__A0 right_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__S sb_0__8_.mem_right_track_58.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A0 sb_0__8_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_45.mux_l1_in_0_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ net18 sb_0__8_.mem_bottom_track_45.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0 net7 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput4 chanx_right_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_15.mux_l2_in_0__201 VGND VGND VPWR VPWR net201 sb_0__8_.mux_bottom_track_15.mux_l2_in_0__201/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_142_ net17 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input63_A gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk sb_0__8_.mem_right_track_22.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_22.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__163__A sb_0__8_.mux_bottom_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_ cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_bottom_track_1.mux_l1_in_1__198 VGND VGND VPWR VPWR net198 sb_0__8_.mux_bottom_track_1.mux_l1_in_1__198/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_125_ sb_0__8_.mux_right_track_16.out VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__8_.mem_right_track_52.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_54.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__158__A sb_0__8_.mux_bottom_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput73 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND VGND VPWR
+ VPWR net73 sky130_fd_sc_hd__buf_2
Xinput62 chany_bottom_in_0[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput40 chany_bottom_in_0[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput51 chany_bottom_in_0[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mux_right_track_6.mux_l2_in_1__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input26_A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_ sb_0__8_.mux_bottom_track_17.out
+ net46 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
X_108_ sb_0__8_.mux_right_track_50.out VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__8_.mem_right_track_2.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_34_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_bottom_track_19.mux_l2_in_0__151 VGND VGND VPWR VPWR net151 sb_0__8_.mux_bottom_track_19.mux_l2_in_0__151/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mux_right_track_18.mux_l2_in_0_ net169 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_18.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_bottom_track_15.mux_l1_in_0__A0 right_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_20.mux_l2_in_0_ net171 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_20.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_2_0_prog_clk sb_0__8_.mem_right_track_8.mem_out\[1\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 chanx_right_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_141_ sb_0__8_.mux_bottom_track_45.out VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input56_A chany_bottom_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_0__8_.mem_right_track_20.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_22.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput150 net150 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__buf_12
XANTENNA_sb_0__8_.mux_right_track_24.mux_l1_in_0__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_124_ sb_0__8_.mux_right_track_18.out VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_10_0_prog_clk cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
+ net204 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput63 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
Xinput74 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND VGND VPWR
+ VPWR net74 sky130_fd_sc_hd__buf_2
XFILLER_88_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput30 chanx_right_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput41 chany_bottom_in_0[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
Xinput52 chany_bottom_in_0[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input19_A chanx_right_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_ sb_0__8_.mux_bottom_track_11.out
+ net49 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_107_ sb_0__8_.mux_right_track_52.out VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_0__8_.mem_right_track_0.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_1.ccff_tail net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_34_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__8_.mem_right_track_28.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1__S cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_0__8_.mem_right_track_8.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_22.mux_l2_in_0__172 VGND VGND VPWR VPWR net172 sb_0__8_.mux_right_track_22.mux_l2_in_0__172/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__8_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_22.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__8_.mux_right_track_18.mux_l1_in_0_ net34 net80 sb_0__8_.mem_right_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_1_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_5_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput6 chanx_right_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_20.mux_l1_in_0_ net35 net69 sb_0__8_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_32.mux_l2_in_0_ sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_32.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_140_ sb_0__8_.mux_bottom_track_47.out VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input49_A chany_bottom_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_16.out sky130_fd_sc_hd__clkbuf_1
XFILLER_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput140 net140 VGND VGND VPWR VPWR chany_bottom_out_0[7] sky130_fd_sc_hd__buf_12
XANTENNA_sb_0__8_.mux_bottom_track_31.mux_l1_in_0__A0 right_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_70_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_123_ sb_0__8_.mux_right_track_20.out VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_6_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput20 chanx_right_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 chanx_right_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_15.out sky130_fd_sc_hd__clkbuf_1
Xinput64 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
Xinput75 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND VGND VPWR
+ VPWR net75 sky130_fd_sc_hd__buf_2
XFILLER_88_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_15.mux_l2_in_0_ net201 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_15.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xinput42 chany_bottom_in_0[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
Xinput53 chany_bottom_in_0[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__8_.mux_right_track_32.mux_l1_in_1_ net177 net41 sb_0__8_.mem_right_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_12_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_ sb_0__8_.mux_bottom_track_5.out
+ net52 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_106_ sb_0__8_.mux_right_track_54.out VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__8_.mem_right_track_26.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_14_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_84_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0 net16 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input31_A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input79_A right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__8_.mem_right_track_40.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_40.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net63 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mux_right_track_40.mux_l1_in_0__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_50.out sky130_fd_sc_hd__clkbuf_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_0__8_.mem_right_track_6.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_77_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput7 chanx_right_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__D sb_0__8_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__8_.mem_bottom_track_5.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput130 net130 VGND VGND VPWR VPWR chany_bottom_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput141 net141 VGND VGND VPWR VPWR chany_bottom_out_0[8] sky130_fd_sc_hd__buf_12
XFILLER_55_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input61_A chany_bottom_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_122_ sb_0__8_.mux_right_track_22.out VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_4.mux_l3_in_0_ sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sb_0__8_.mem_right_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xinput21 chanx_right_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xinput10 chanx_right_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput32 chanx_right_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput54 chany_bottom_in_0[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 chany_bottom_in_0[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput65 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
Xinput76 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND VGND VPWR
+ VPWR net76 sky130_fd_sc_hd__clkbuf_2
Xsb_0__8_.mux_right_track_32.mux_l1_in_0_ net75 net79 sb_0__8_.mem_right_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_38.out sky130_fd_sc_hd__clkbuf_1
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_44.mux_l2_in_0_ sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_105_ sb_0__8_.mux_right_track_56.out VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mux_bottom_track_7.mux_l2_in_0_ sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_bottom_track_7.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_right_track_4.mux_l2_in_1_ net181 net56 sb_0__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input24_A chanx_right_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_bottom_track_15.mux_l1_in_0_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ net31 sb_0__8_.mem_bottom_track_15.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__196 VGND VGND VPWR VPWR net196
+ cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__196/LO sky130_fd_sc_hd__conb_1
XFILLER_16_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_44.mux_l1_in_1_ net184 net48 sb_0__8_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__8_.mem_bottom_track_45.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_0__8_.mem_right_track_38.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_40.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_bottom_track_7.mux_l1_in_1_ net162 right_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_0__8_.mem_bottom_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__A1 net22 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_5.out sky130_fd_sc_hd__clkbuf_1
XFILLER_76_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 chanx_right_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net66 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__8_.mem_bottom_track_3.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__8_.mem_right_track_46.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_46.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__S cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput142 net142 VGND VGND VPWR VPWR chany_bottom_out_0[9] sky130_fd_sc_hd__buf_12
Xoutput120 net120 VGND VGND VPWR VPWR chany_bottom_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chany_bottom_out_0[26] sky130_fd_sc_hd__buf_12
XFILLER_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_right_track_2.mux_l2_in_1__170 VGND VGND VPWR VPWR net170 sb_0__8_.mux_right_track_2.mux_l2_in_1__170/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_121_ sb_0__8_.mux_right_track_24.out VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input54_A chany_bottom_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput77 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND
+ VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xinput66 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
Xinput22 chanx_right_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
Xinput11 chanx_right_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput44 chany_bottom_in_0[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput33 chany_bottom_in_0[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput55 chany_bottom_in_0[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_10_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_104_ sb_0__8_.mux_right_track_58.out VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_4.mux_l2_in_0_ sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__8_.mem_bottom_track_13.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input17_A chanx_right_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_right_track_44.mux_l1_in_0_ net73 net77 sb_0__8_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input9_A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__8_.mem_bottom_track_35.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__8_.mux_right_track_56.mux_l2_in_0_ net190 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_56.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_7.mux_l1_in_0_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ net27 sb_0__8_.mem_bottom_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_4.mux_l1_in_1_ net76 net73 sb_0__8_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 chanx_right_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
Xsb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__8_.mem_right_track_14.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_15_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__8_.mem_right_track_44.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_46.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xoutput143 net143 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
Xoutput121 net121 VGND VGND VPWR VPWR chany_bottom_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput110 net110 VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_12
Xoutput132 net132 VGND VGND VPWR VPWR chany_bottom_out_0[27] sky130_fd_sc_hd__buf_12
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_0_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_120_ sb_0__8_.mux_right_track_26.out VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input47_A chany_bottom_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput78 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND
+ VPWR VPWR net78 sky130_fd_sc_hd__buf_2
Xinput67 isol_n VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 chanx_right_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xinput12 chanx_right_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput45 chany_bottom_in_0[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput56 chany_bottom_in_0[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 chany_bottom_in_0[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_ net197 net23 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__8_.mem_bottom_track_11.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_90_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 net205 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_13_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_ net17 net61 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_4.mux_l1_in_0_ net70 net79 sb_0__8_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cby_0__8_.cby_0__1_.ccff_tail
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input77_A right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__8_.mem_bottom_track_19.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_19.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__8_.mux_bottom_track_13.mux_l2_in_0__200 VGND VGND VPWR VPWR net200 sb_0__8_.mux_bottom_track_13.mux_l2_in_0__200/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_0__8_.mem_right_track_12.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_56.mux_l1_in_0_ net54 net71 sb_0__8_.mem_right_track_56.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__S cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_54.mux_l2_in_0__189 VGND VGND VPWR VPWR net189 sb_0__8_.mux_right_track_54.mux_l2_in_0__189/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput144 net144 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_ cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xoutput100 net100 VGND VGND VPWR VPWR chanx_right_out[25] sky130_fd_sc_hd__buf_12
Xoutput122 net122 VGND VGND VPWR VPWR chany_bottom_out_0[18] sky130_fd_sc_hd__buf_12
Xoutput111 net111 VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_12
Xoutput133 net133 VGND VGND VPWR VPWR chany_bottom_out_0[28] sky130_fd_sc_hd__buf_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 chanx_right_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XFILLER_61_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput79 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND
+ VPWR VPWR net79 sky130_fd_sc_hd__buf_2
Xinput24 chanx_right_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput35 chany_bottom_in_0[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
Xinput46 chany_bottom_in_0[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput68 net206 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
Xinput57 chany_bottom_in_0[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_ net55 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_bottom_track_29.mux_l1_in_0__A0 right_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_1__A1 right_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A0 sb_0__8_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2 net207 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_16
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0 net8 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_ sb_0__8_.mux_bottom_track_31.out
+ net38 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input22_A chanx_right_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_0__8_.mem_bottom_track_17.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_19.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2__A0 net57 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_right_track_38.mux_l1_in_0__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput145 net145 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
Xoutput101 net101 VGND VGND VPWR VPWR chanx_right_out[26] sky130_fd_sc_hd__buf_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xoutput123 net123 VGND VGND VPWR VPWR chany_bottom_out_0[19] sky130_fd_sc_hd__buf_12
Xoutput134 net134 VGND VGND VPWR VPWR chany_bottom_out_0[29] sky130_fd_sc_hd__buf_12
Xoutput112 net112 VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_12
XANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__8_.mem_bottom_track_31.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_31.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput25 chanx_right_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 chanx_right_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput36 chany_bottom_in_0[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput69 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND VGND VPWR
+ VPWR net69 sky130_fd_sc_hd__clkbuf_4
Xsb_0__8_.mux_right_track_14.mux_l2_in_0_ sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_14.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xinput58 chany_bottom_in_0[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
Xinput47 chany_bottom_in_0[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input52_A chany_bottom_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_ cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_0__8_.mux_right_track_14.mux_l1_in_1_ net167 net61 sb_0__8_.mem_right_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__8_.mem_right_track_32.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_32.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xhold3 prog_reset VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_ sb_0__8_.mux_bottom_track_19.out
+ net45 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input15_A chanx_right_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input7_A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_20.mux_l2_in_0__171 VGND VGND VPWR VPWR net171 sb_0__8_.mux_right_track_20.mux_l2_in_0__171/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_bottom_track_5.mux_l1_in_0__A0 right_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A0 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_bottom_track_45.mux_l1_in_0__A0 right_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput146 net146 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
Xoutput102 net102 VGND VGND VPWR VPWR chanx_right_out[27] sky130_fd_sc_hd__buf_12
Xoutput113 net113 VGND VGND VPWR VPWR chany_bottom_out_0[0] sky130_fd_sc_hd__buf_12
Xoutput124 net124 VGND VGND VPWR VPWR chany_bottom_out_0[1] sky130_fd_sc_hd__buf_12
Xoutput135 net135 VGND VGND VPWR VPWR chany_bottom_out_0[2] sky130_fd_sc_hd__buf_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__8_.mem_bottom_track_29.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_31.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput15 chanx_right_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 chanx_right_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput59 chany_bottom_in_0[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
Xinput37 chany_bottom_in_0[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput48 chany_bottom_in_0[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input45_A chany_bottom_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_9.mux_l2_in_0__163 VGND VGND VPWR VPWR net163 sb_0__8_.mux_bottom_track_9.mux_l2_in_0__163/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_40_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_14.mux_l1_in_0_ net74 net78 sb_0__8_.mem_right_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mux_right_track_36.mux_l2_in_0__179 VGND VGND VPWR VPWR net179 sb_0__8_.mux_right_track_36.mux_l2_in_0__179/LO
+ sky130_fd_sc_hd__conb_1
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__194 VGND VGND VPWR VPWR net194
+ cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__194/LO sky130_fd_sc_hd__conb_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 net203 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__8_.mem_right_track_30.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_32.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_90_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_26.mux_l2_in_0_ net174 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_26.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__8_.mux_right_track_54.mux_l1_in_0__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_ sb_0__8_.mux_bottom_track_7.out
+ net51 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A0 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_11.out sky130_fd_sc_hd__clkbuf_1
XFILLER_85_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_2.mux_l2_in_1__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_2_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_48.mux_l1_in_1__186 VGND VGND VPWR VPWR net186 sb_0__8_.mux_right_track_48.mux_l1_in_1__186/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__8_.mux_bottom_track_11.mux_l2_in_0_ net199 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_11.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_12_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__8_.mem_right_track_38.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_38.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input75_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput103 net103 VGND VGND VPWR VPWR chanx_right_out[28] sky130_fd_sc_hd__buf_12
Xoutput125 net125 VGND VGND VPWR VPWR chany_bottom_out_0[20] sky130_fd_sc_hd__buf_12
Xoutput114 net114 VGND VGND VPWR VPWR chany_bottom_out_0[10] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__buf_12
Xoutput136 net136 VGND VGND VPWR VPWR chany_bottom_out_0[3] sky130_fd_sc_hd__buf_12
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_bottom_track_11.mux_l1_in_0__A0 right_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput16 chanx_right_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
Xinput27 chanx_right_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput49 chany_bottom_in_0[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xinput38 chany_bottom_in_0[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0 net17 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input38_A chany_bottom_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_159_ sb_0__8_.mux_bottom_track_9.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_7_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_40.out sky130_fd_sc_hd__clkbuf_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold5 net68 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_ sb_0__8_.mux_bottom_track_1.out
+ net54 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__8_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_34.out sky130_fd_sc_hd__clkbuf_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input20_A chanx_right_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_right_track_26.mux_l1_in_0_ net38 net72 sb_0__8_.mem_right_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_0.mux_l3_in_0_ sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_0__8_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_38.mux_l2_in_0_ net180 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_38.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__142__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_33.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_0__8_.mem_right_track_36.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_38.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mux_right_track_40.mux_l2_in_0_ net182 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_40.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input68_A net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
XANTENNA__137__A net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput148 net148 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__buf_12
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput104 net104 VGND VGND VPWR VPWR chanx_right_out[29] sky130_fd_sc_hd__buf_12
Xoutput115 net115 VGND VGND VPWR VPWR chany_bottom_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput137 net137 VGND VGND VPWR VPWR chany_bottom_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chany_bottom_out_0[21] sky130_fd_sc_hd__buf_12
XFILLER_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_bottom_track_3.mux_l2_in_0_ net153 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_3.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_0.mux_l2_in_1_ net164 net44 sb_0__8_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput17 chanx_right_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
Xinput28 chanx_right_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xsb_0__8_.mux_bottom_track_11.mux_l1_in_0_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ net29 sb_0__8_.mem_bottom_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xinput39 chany_bottom_in_0[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__8_.mem_right_track_50.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_50.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_1.out sky130_fd_sc_hd__clkbuf_2
XFILLER_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_8.out sky130_fd_sc_hd__clkbuf_1
X_158_ sb_0__8_.mux_bottom_track_11.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__150__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_1__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_bottom_track_51.mux_l2_in_0__161 VGND VGND VPWR VPWR net161 sb_0__8_.mux_bottom_track_51.mux_l2_in_0__161/LO
+ sky130_fd_sc_hd__conb_1
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input50_A chany_bottom_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold6 net212 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1 net23 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__145__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A0 sb_0__8_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A0 sb_0__8_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input13_A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_10_0_prog_clk cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
+ net204 VGND VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_bottom_track_35.mux_l2_in_0__156 VGND VGND VPWR VPWR net156 sb_0__8_.mux_bottom_track_35.mux_l2_in_0__156/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input5_A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_56.out sky130_fd_sc_hd__clkbuf_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_18.mux_l2_in_0__169 VGND VGND VPWR VPWR net169 sb_0__8_.mux_right_track_18.mux_l2_in_0__169/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput149 net149 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__buf_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput116 net116 VGND VGND VPWR VPWR chany_bottom_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput138 net138 VGND VGND VPWR VPWR chany_bottom_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput127 net127 VGND VGND VPWR VPWR chany_bottom_out_0[22] sky130_fd_sc_hd__buf_12
Xoutput105 net105 VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_12
XANTENNA__153__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_0.mux_l2_in_0_ sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_36_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input80_A right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_right_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_38.mux_l1_in_0_ net45 net70 sb_0__8_.mem_right_track_38.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xinput29 chanx_right_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__8_.mem_right_track_48.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_50.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_93_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__148__A sb_0__8_.mux_bottom_track_31.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail net67 VGND
+ VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_0__S sb_0__8_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_right_track_40.mux_l1_in_0_ net46 net71 sb_0__8_.mem_right_track_40.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_95_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_52.mux_l2_in_0_ net188 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_52.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_bottom_track_3.mux_l1_in_0_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ net25 sb_0__8_.mem_bottom_track_3.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_157_ sb_0__8_.mux_bottom_track_13.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_49.out sky130_fd_sc_hd__clkbuf_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_0.mux_l1_in_1_ net74 net71 sb_0__8_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_1__A1 right_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input43_A chany_bottom_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold7 net2 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_1__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__161__A sb_0__8_.mux_bottom_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_9_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_11_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_bottom_track_35.mux_l2_in_0_ net156 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_35.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__8_.mem_right_track_56.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_56.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_88_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_1__S sb_0__8_.mem_right_track_58.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__156__A sb_0__8_.mux_bottom_track_15.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_0__8_.mem_right_track_4.mem_out\[1\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_52.mux_l2_in_0__188 VGND VGND VPWR VPWR net188 sb_0__8_.mux_right_track_52.mux_l2_in_0__188/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output112_A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_bottom_track_7.mux_l1_in_1__162 VGND VGND VPWR VPWR net162 sb_0__8_.mux_bottom_track_7.mux_l1_in_1__162/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput128 net128 VGND VGND VPWR VPWR chany_bottom_out_0[23] sky130_fd_sc_hd__buf_12
Xoutput117 net117 VGND VGND VPWR VPWR chany_bottom_out_0[13] sky130_fd_sc_hd__buf_12
Xoutput139 net139 VGND VGND VPWR VPWR chany_bottom_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput106 net106 VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_12
XFILLER_70_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\] net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_right_track_34.mux_l1_in_1__178 VGND VGND VPWR VPWR net178 sb_0__8_.mux_right_track_34.mux_l1_in_1__178/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput19 chanx_right_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input73_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_11_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_156_ sb_0__8_.mux_bottom_track_15.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__159__A sb_0__8_.mux_bottom_track_9.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_0.mux_l1_in_0_ net80 net77 sb_0__8_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk sb_0__8_.mem_right_track_24.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_24.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail net67 VGND
+ VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold8 net214 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input36_A chany_bottom_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_139_ sb_0__8_.mux_bottom_track_49.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_10.mux_l3_in_0_ sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_0__8_.mem_right_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__8_.mem_right_track_54.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_56.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__8_.mux_right_track_52.mux_l1_in_0_ net52 net69 sb_0__8_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__8_.mem_right_track_4.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_bottom_track_35.mux_l1_in_0_ right_width_0_height_0_subtile_3__pin_inpad_0_
+ net12 sb_0__8_.mem_bottom_track_35.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_10.mux_l2_in_1_ net165 net59 sb_0__8_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_bottom_track_47.mux_l2_in_0_ net158 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_47.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput107 net107 VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_12
Xoutput118 net118 VGND VGND VPWR VPWR chany_bottom_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput129 net129 VGND VGND VPWR VPWR chany_bottom_out_0[24] sky130_fd_sc_hd__buf_12
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ cby_0__8_.cby_0__1_.mem_right_ipin_0.ccff_tail net204 VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_1__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input66_A gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_155_ sb_0__8_.mux_bottom_track_17.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__8_.mem_bottom_track_29.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk sb_0__8_.mem_right_track_22.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_24.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A0 sb_0__8_.mux_bottom_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold9 net1 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input29_A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_138_ sb_0__8_.mux_bottom_track_51.out VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__S cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_49.mux_l2_in_0__159 VGND VGND VPWR VPWR net159 sb_0__8_.mux_bottom_track_49.mux_l2_in_0__159/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output135_A net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0 net56 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_26.mux_l1_in_0__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__8_.mem_right_track_2.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_10.mux_l2_in_0_ sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mux_right_track_8.mux_l2_in_1__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input11_A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__8_.mem_bottom_track_1.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput119 net119 VGND VGND VPWR VPWR chany_bottom_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput108 net108 VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_12
XANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput90 net90 VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_12
XFILLER_55_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input3_A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_171_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
Xsb_0__8_.mux_right_track_10.mux_l1_in_1_ net76 net73 sb_0__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_89_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input59_A chany_bottom_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_bottom_track_17.mux_l1_in_0__A0 right_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_bottom_track_47.mux_l1_in_0_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ net19 sb_0__8_.mem_bottom_track_47.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_154_ sb_0__8_.mux_bottom_track_19.out VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__8_.mem_bottom_track_19.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_83_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_137_ net22 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_16.mux_l1_in_1__168 VGND VGND VPWR VPWR net168 sb_0__8_.mux_right_track_16.mux_l1_in_1__168/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input41_A chany_bottom_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__8_.mux_right_track_26.mux_l1_in_0__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_8_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_46.mux_l1_in_1__185 VGND VGND VPWR VPWR net185 sb_0__8_.mux_right_track_46.mux_l1_in_1__185/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_2_0_prog_clk sb_0__8_.mem_right_track_10.mem_out\[1\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput109 net109 VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_12
Xsb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__8_.mem_bottom_track_1.ccff_head
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xoutput91 net91 VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_12
XFILLER_63_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net64 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__8_.mem_right_track_42.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_42.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_170_ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_29.mux_l2_in_0__152 VGND VGND VPWR VPWR net152 sb_0__8_.mux_bottom_track_29.mux_l2_in_0__152/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__8_.mux_right_track_10.mux_l1_in_0_ net70 net79 sb_0__8_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_22.mux_l2_in_0_ net172 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_right_track_22.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hold12_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_153_ net5 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input71_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__8_.mem_bottom_track_7.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_10_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_136_ net23 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0__S cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input34_A chany_bottom_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_119_ sb_0__8_.mux_right_track_28.out VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_bottom_track_33.mux_l1_in_0__A0 right_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A0 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_0__8_.mem_right_track_10.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput81 net81 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
Xoutput92 net92 VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_12
Xsb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__8_.mem_bottom_track_47.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_47.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__8_.mem_right_track_40.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_42.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__8_.mux_right_track_0.mux_l2_in_1__164 VGND VGND VPWR VPWR net164 sb_0__8_.mux_right_track_0.mux_l2_in_1__164/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_54_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_3_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_30.out sky130_fd_sc_hd__clkbuf_1
XFILLER_3_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__S cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_152_ net6 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input64_A gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
+ clknet_4_10_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_0__A0 right_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__8_.mem_bottom_track_5.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__8_.mem_right_track_48.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_48.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_74_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_22.mux_l1_in_0_ net36 net70 sb_0__8_.mem_right_track_22.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
X_135_ net24 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xsb_0__8_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_24.out sky130_fd_sc_hd__clkbuf_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_34.mux_l2_in_0_ sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_34.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__8_.mux_right_track_58.mux_l1_in_1__191 VGND VGND VPWR VPWR net191 sb_0__8_.mux_right_track_58.mux_l1_in_1__191/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input27_A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_118_ sb_0__8_.mux_right_track_30.out VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_8_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_18.out sky130_fd_sc_hd__clkbuf_1
XFILLER_84_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__8_.mux_bottom_track_17.mux_l2_in_0_ net202 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_17.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mux_right_track_34.mux_l1_in_1_ net178 net42 sb_0__8_.mem_right_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__8_.mem_bottom_track_15.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_15.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_bottom_track_33.mux_l2_in_0__155 VGND VGND VPWR VPWR net155 sb_0__8_.mux_bottom_track_33.mux_l2_in_0__155/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_0__8_.mem_right_track_10.ccff_head
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_17.out sky130_fd_sc_hd__clkbuf_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput82 net82 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
XANTENNA_hold5_A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput93 net93 VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_12
Xsb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__8_.mem_bottom_track_45.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_47.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__8_.mem_right_track_16.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_16.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_151_ net7 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input57_A chany_bottom_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_28.mux_l1_in_1__175 VGND VGND VPWR VPWR net175 sb_0__8_.mux_right_track_28.mux_l1_in_1__175/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_1__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A0 sb_0__8_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__S cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__8_.mem_right_track_46.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_48.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_134_ net3 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
XFILLER_23_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_51.out sky130_fd_sc_hd__clkbuf_1
XFILLER_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0 sb_0__8_.mux_bottom_track_15.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
+ clknet_4_10_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_117_ sb_0__8_.mux_right_track_32.out VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__8_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_46.out sky130_fd_sc_hd__clkbuf_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__8_.mux_right_track_6.mux_l3_in_0_ sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_0__8_.mem_right_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_34.mux_l1_in_0_ net76 net80 sb_0__8_.mem_right_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_75_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_45.out sky130_fd_sc_hd__clkbuf_1
XFILLER_90_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__8_.mem_bottom_track_13.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__8_.mux_right_track_46.mux_l2_in_0_ sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_46.ccff_tail
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_right_track_50.mux_l2_in_0__187 VGND VGND VPWR VPWR net187 sb_0__8_.mux_right_track_50.mux_l2_in_0__187/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_bottom_track_9.mux_l2_in_0_ net163 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_11.ccff_head VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput94 net94 VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_12
Xoutput83 net83 VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_12
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_0__8_.mux_right_track_6.mux_l2_in_1_ net192 net57 sb_0__8_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_bottom_track_17.mux_l1_in_0_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ net32 sb_0__8_.mem_bottom_track_17.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_7_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__S cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__8_.mux_right_track_32.mux_l1_in_1__177 VGND VGND VPWR VPWR net177 sb_0__8_.mux_right_track_32.mux_l1_in_1__177/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_29.mux_l2_in_0_ net152 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_29.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mux_right_track_46.mux_l1_in_1_ net185 net49 sb_0__8_.mem_right_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_95_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__8_.mux_bottom_track_31.mux_l2_in_0_ net154 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__8_.mem_bottom_track_31.ccff_tail VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_0__8_.mem_right_track_14.ccff_tail
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_16.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_150_ net8 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold10_A ccff_head_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_133_ sb_0__8_.mux_right_track_0.out VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__110__A sb_0__8_.mux_right_track_46.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_7.out sky130_fd_sc_hd__clkbuf_2
XFILLER_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_116_ sb_0__8_.mux_right_track_34.out VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
+ clknet_4_10_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input32_A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_12_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__197 VGND VGND VPWR VPWR net197
+ cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__197/LO sky130_fd_sc_hd__conb_1
XFILLER_1_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_1__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput95 net95 VGND VGND VPWR VPWR chanx_right_out[20] sky130_fd_sc_hd__buf_12
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput84 net84 VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_12
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__8_.mux_right_track_52.mux_l2_in_0__A0 net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_6.mux_l2_in_0_ sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_46.mux_l1_in_0_ net74 net78 sb_0__8_.mem_right_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_9_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__8_.mux_right_track_58.mux_l2_in_0_ sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_0_X sb_0__8_.mem_bottom_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mux_bottom_track_9.mux_l1_in_0_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ net28 sb_0__8_.mem_bottom_track_9.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_ net194 sb_0__8_.mux_bottom_track_49.out
+ cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__8_.mux_right_track_6.mux_l1_in_1_ net74 net71 sb_0__8_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_5.mux_l2_in_0__160 VGND VGND VPWR VPWR net160 sb_0__8_.mux_bottom_track_5.mux_l2_in_0__160/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_29.mux_l1_in_0_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ net9 sb_0__8_.mem_bottom_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_132_ sb_0__8_.mux_right_track_2.out VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input62_A chany_bottom_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_31.mux_l1_in_0_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ net10 sb_0__8_.mem_bottom_track_31.mem_out\[0\] VGND VGND VPWR VPWR sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__8_.mux_right_track_58.mux_l1_in_1_ net191 net33 sb_0__8_.mem_right_track_58.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_73_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__8_.mem_bottom_track_33.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_bottom_track_33.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__8_.mux_bottom_track_47.mux_l2_in_0__158 VGND VGND VPWR VPWR net158 sb_0__8_.mux_bottom_track_47.mux_l2_in_0__158/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_ net13 net35 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ sb_0__8_.mux_right_track_36.out VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net204 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_ cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_0__8_.cby_0__1_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input25_A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net204 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__8_.mem_right_track_34.mem_out\[0\]
+ net204 VGND VGND VPWR VPWR sb_0__8_.mem_right_track_34.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput96 net96 VGND VGND VPWR VPWR chanx_right_out[21] sky130_fd_sc_hd__buf_12
Xoutput85 net85 VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_12
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__8_.mux_right_track_8.mux_l2_in_1__193 VGND VGND VPWR VPWR net193 sb_0__8_.mux_right_track_8.mux_l2_in_1__193/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
+ clknet_4_10_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_ cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
.ends

