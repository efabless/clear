magic
tech sky130A
magscale 1 2
timestamp 1656943068
<< viali >>
rect 5181 14569 5215 14603
rect 4997 14229 5031 14263
rect 4169 14025 4203 14059
rect 4537 14025 4571 14059
rect 4997 14025 5031 14059
rect 5457 14025 5491 14059
rect 10333 14025 10367 14059
rect 14657 14025 14691 14059
rect 13093 13957 13127 13991
rect 14289 13957 14323 13991
rect 14381 13957 14415 13991
rect 15301 13957 15335 13991
rect 16221 13957 16255 13991
rect 5365 13889 5399 13923
rect 5825 13889 5859 13923
rect 10517 13889 10551 13923
rect 10885 13889 10919 13923
rect 12817 13889 12851 13923
rect 15025 13889 15059 13923
rect 16681 13889 16715 13923
rect 17049 13889 17083 13923
rect 4629 13821 4663 13855
rect 4721 13821 4755 13855
rect 5641 13821 5675 13855
rect 6101 13821 6135 13855
rect 6653 13821 6687 13855
rect 11253 13821 11287 13855
rect 13737 13821 13771 13855
rect 15209 13821 15243 13855
rect 16313 13821 16347 13855
rect 14841 13753 14875 13787
rect 16865 13753 16899 13787
rect 6469 13685 6503 13719
rect 2789 13481 2823 13515
rect 3617 13481 3651 13515
rect 6285 13481 6319 13515
rect 13415 13481 13449 13515
rect 2973 13345 3007 13379
rect 5181 13345 5215 13379
rect 5917 13345 5951 13379
rect 6561 13345 6595 13379
rect 3249 13277 3283 13311
rect 5733 13277 5767 13311
rect 13344 13277 13378 13311
rect 3893 13209 3927 13243
rect 4445 13209 4479 13243
rect 4905 13209 4939 13243
rect 6745 13209 6779 13243
rect 3157 13141 3191 13175
rect 4077 13141 4111 13175
rect 4537 13141 4571 13175
rect 4997 13141 5031 13175
rect 5365 13141 5399 13175
rect 5825 13141 5859 13175
rect 6653 13141 6687 13175
rect 7113 13141 7147 13175
rect 15209 13141 15243 13175
rect 4537 12937 4571 12971
rect 4629 12937 4663 12971
rect 5733 12937 5767 12971
rect 6193 12937 6227 12971
rect 7021 12937 7055 12971
rect 13461 12937 13495 12971
rect 14197 12937 14231 12971
rect 2145 12869 2179 12903
rect 5365 12869 5399 12903
rect 5181 12801 5215 12835
rect 5825 12801 5859 12835
rect 6561 12801 6595 12835
rect 7389 12801 7423 12835
rect 7481 12801 7515 12835
rect 8125 12801 8159 12835
rect 13369 12801 13403 12835
rect 13921 12801 13955 12835
rect 4721 12733 4755 12767
rect 5641 12733 5675 12767
rect 7665 12733 7699 12767
rect 13645 12733 13679 12767
rect 2605 12665 2639 12699
rect 2513 12597 2547 12631
rect 4169 12597 4203 12631
rect 6377 12597 6411 12631
rect 6929 12597 6963 12631
rect 7941 12597 7975 12631
rect 9689 12597 9723 12631
rect 13001 12597 13035 12631
rect 11805 12393 11839 12427
rect 14933 12325 14967 12359
rect 2237 12257 2271 12291
rect 3433 12257 3467 12291
rect 4445 12257 4479 12291
rect 4813 12257 4847 12291
rect 6009 12257 6043 12291
rect 7021 12257 7055 12291
rect 7849 12257 7883 12291
rect 9505 12257 9539 12291
rect 10241 12257 10275 12291
rect 10425 12257 10459 12291
rect 12541 12257 12575 12291
rect 12909 12257 12943 12291
rect 13645 12257 13679 12291
rect 14565 12257 14599 12291
rect 14749 12257 14783 12291
rect 17785 12257 17819 12291
rect 1961 12189 1995 12223
rect 3249 12189 3283 12223
rect 4905 12189 4939 12223
rect 5917 12189 5951 12223
rect 6837 12189 6871 12223
rect 10609 12189 10643 12223
rect 12449 12189 12483 12223
rect 13185 12189 13219 12223
rect 17693 12189 17727 12223
rect 18061 12189 18095 12223
rect 2329 12121 2363 12155
rect 6285 12121 6319 12155
rect 8309 12121 8343 12155
rect 13093 12121 13127 12155
rect 1777 12053 1811 12087
rect 2421 12053 2455 12087
rect 2789 12053 2823 12087
rect 2881 12053 2915 12087
rect 3341 12053 3375 12087
rect 3801 12053 3835 12087
rect 4169 12053 4203 12087
rect 4261 12053 4295 12087
rect 4997 12053 5031 12087
rect 5365 12053 5399 12087
rect 5457 12053 5491 12087
rect 5825 12053 5859 12087
rect 6469 12053 6503 12087
rect 6929 12053 6963 12087
rect 7297 12053 7331 12087
rect 7665 12053 7699 12087
rect 7757 12053 7791 12087
rect 8125 12053 8159 12087
rect 8953 12053 8987 12087
rect 9321 12053 9355 12087
rect 9413 12053 9447 12087
rect 9781 12053 9815 12087
rect 10149 12053 10183 12087
rect 11989 12053 12023 12087
rect 12357 12053 12391 12087
rect 13553 12053 13587 12087
rect 14105 12053 14139 12087
rect 14473 12053 14507 12087
rect 17049 12053 17083 12087
rect 17233 12053 17267 12087
rect 17601 12053 17635 12087
rect 18245 12053 18279 12087
rect 2513 11849 2547 11883
rect 2605 11849 2639 11883
rect 3065 11849 3099 11883
rect 4077 11849 4111 11883
rect 4997 11849 5031 11883
rect 5457 11849 5491 11883
rect 5549 11849 5583 11883
rect 6009 11849 6043 11883
rect 6929 11849 6963 11883
rect 7297 11849 7331 11883
rect 7757 11849 7791 11883
rect 8125 11849 8159 11883
rect 8953 11849 8987 11883
rect 9413 11849 9447 11883
rect 10793 11849 10827 11883
rect 12909 11849 12943 11883
rect 17141 11849 17175 11883
rect 17693 11849 17727 11883
rect 17969 11849 18003 11883
rect 2053 11781 2087 11815
rect 6469 11781 6503 11815
rect 9045 11781 9079 11815
rect 9873 11781 9907 11815
rect 18061 11781 18095 11815
rect 1685 11713 1719 11747
rect 2145 11713 2179 11747
rect 2973 11713 3007 11747
rect 3433 11713 3467 11747
rect 3985 11713 4019 11747
rect 4445 11713 4479 11747
rect 8217 11713 8251 11747
rect 10241 11713 10275 11747
rect 10701 11713 10735 11747
rect 11897 11713 11931 11747
rect 13461 11713 13495 11747
rect 15301 11713 15335 11747
rect 17049 11713 17083 11747
rect 1961 11645 1995 11679
rect 3249 11645 3283 11679
rect 4537 11645 4571 11679
rect 4721 11645 4755 11679
rect 5365 11645 5399 11679
rect 6837 11645 6871 11679
rect 7389 11645 7423 11679
rect 7481 11645 7515 11679
rect 8309 11645 8343 11679
rect 9137 11645 9171 11679
rect 10885 11645 10919 11679
rect 11989 11645 12023 11679
rect 12081 11645 12115 11679
rect 13553 11645 13587 11679
rect 13645 11645 13679 11679
rect 15071 11645 15105 11679
rect 15209 11645 15243 11679
rect 17233 11645 17267 11679
rect 12449 11577 12483 11611
rect 15853 11577 15887 11611
rect 16681 11577 16715 11611
rect 1501 11509 1535 11543
rect 3801 11509 3835 11543
rect 5917 11509 5951 11543
rect 8585 11509 8619 11543
rect 10333 11509 10367 11543
rect 11253 11509 11287 11543
rect 11529 11509 11563 11543
rect 13093 11509 13127 11543
rect 13921 11509 13955 11543
rect 14749 11509 14783 11543
rect 15669 11509 15703 11543
rect 18337 11509 18371 11543
rect 1685 11305 1719 11339
rect 2605 11305 2639 11339
rect 4537 11305 4571 11339
rect 8953 11305 8987 11339
rect 14933 11305 14967 11339
rect 17049 11305 17083 11339
rect 18061 11305 18095 11339
rect 2145 11237 2179 11271
rect 3433 11237 3467 11271
rect 5549 11237 5583 11271
rect 6377 11237 6411 11271
rect 8033 11237 8067 11271
rect 9321 11237 9355 11271
rect 10149 11237 10183 11271
rect 10977 11237 11011 11271
rect 14105 11237 14139 11271
rect 16497 11237 16531 11271
rect 18429 11237 18463 11271
rect 2789 11169 2823 11203
rect 3985 11169 4019 11203
rect 4721 11169 4755 11203
rect 4905 11169 4939 11203
rect 6193 11169 6227 11203
rect 6837 11169 6871 11203
rect 6929 11169 6963 11203
rect 7757 11169 7791 11203
rect 8493 11169 8527 11203
rect 8585 11169 8619 11203
rect 9781 11169 9815 11203
rect 9965 11169 9999 11203
rect 10609 11169 10643 11203
rect 10793 11169 10827 11203
rect 11529 11169 11563 11203
rect 12909 11169 12943 11203
rect 13001 11169 13035 11203
rect 14657 11169 14691 11203
rect 15761 11169 15795 11203
rect 17509 11169 17543 11203
rect 17601 11169 17635 11203
rect 1961 11101 1995 11135
rect 2329 11101 2363 11135
rect 3065 11101 3099 11135
rect 4077 11101 4111 11135
rect 4997 11101 5031 11135
rect 5917 11101 5951 11135
rect 6745 11101 6779 11135
rect 9689 11101 9723 11135
rect 10517 11101 10551 11135
rect 13093 11101 13127 11135
rect 13921 11101 13955 11135
rect 14473 11101 14507 11135
rect 16037 11101 16071 11135
rect 16681 11101 16715 11135
rect 17877 11101 17911 11135
rect 18245 11101 18279 11135
rect 2973 11033 3007 11067
rect 6009 11033 6043 11067
rect 7665 11033 7699 11067
rect 9137 11033 9171 11067
rect 11437 11033 11471 11067
rect 14565 11033 14599 11067
rect 15577 11033 15611 11067
rect 1501 10965 1535 10999
rect 4169 10965 4203 10999
rect 5365 10965 5399 10999
rect 7205 10965 7239 10999
rect 7573 10965 7607 10999
rect 8401 10965 8435 10999
rect 11345 10965 11379 10999
rect 11805 10965 11839 10999
rect 13461 10965 13495 10999
rect 15117 10965 15151 10999
rect 15485 10965 15519 10999
rect 16221 10965 16255 10999
rect 17417 10965 17451 10999
rect 2513 10761 2547 10795
rect 2697 10761 2731 10795
rect 3157 10761 3191 10795
rect 4261 10761 4295 10795
rect 5273 10761 5307 10795
rect 6101 10761 6135 10795
rect 7757 10761 7791 10795
rect 8125 10761 8159 10795
rect 8493 10761 8527 10795
rect 8953 10761 8987 10795
rect 9413 10761 9447 10795
rect 10241 10761 10275 10795
rect 10609 10761 10643 10795
rect 10885 10761 10919 10795
rect 11253 10761 11287 10795
rect 11897 10761 11931 10795
rect 12909 10761 12943 10795
rect 13277 10761 13311 10795
rect 13737 10761 13771 10795
rect 14473 10761 14507 10795
rect 15301 10761 15335 10795
rect 15761 10761 15795 10795
rect 16681 10761 16715 10795
rect 17049 10761 17083 10795
rect 17509 10761 17543 10795
rect 1593 10693 1627 10727
rect 2053 10693 2087 10727
rect 3617 10693 3651 10727
rect 4629 10693 4663 10727
rect 14381 10693 14415 10727
rect 15209 10693 15243 10727
rect 18429 10693 18463 10727
rect 3065 10625 3099 10659
rect 4721 10625 4755 10659
rect 6009 10625 6043 10659
rect 6745 10625 6779 10659
rect 7665 10625 7699 10659
rect 9321 10625 9355 10659
rect 10149 10625 10183 10659
rect 13369 10625 13403 10659
rect 16129 10625 16163 10659
rect 17877 10625 17911 10659
rect 18245 10625 18279 10659
rect 1777 10557 1811 10591
rect 1961 10557 1995 10591
rect 3341 10557 3375 10591
rect 4169 10557 4203 10591
rect 4813 10557 4847 10591
rect 5181 10557 5215 10591
rect 6837 10557 6871 10591
rect 6929 10557 6963 10591
rect 7849 10557 7883 10591
rect 8585 10557 8619 10591
rect 8677 10557 8711 10591
rect 9505 10557 9539 10591
rect 10333 10557 10367 10591
rect 11989 10557 12023 10591
rect 12173 10557 12207 10591
rect 13553 10557 13587 10591
rect 14565 10557 14599 10591
rect 15393 10557 15427 10591
rect 16221 10557 16255 10591
rect 16313 10557 16347 10591
rect 17141 10557 17175 10591
rect 17233 10557 17267 10591
rect 6377 10489 6411 10523
rect 12449 10489 12483 10523
rect 18061 10489 18095 10523
rect 2421 10421 2455 10455
rect 5549 10421 5583 10455
rect 7297 10421 7331 10455
rect 9781 10421 9815 10455
rect 11529 10421 11563 10455
rect 12633 10421 12667 10455
rect 14013 10421 14047 10455
rect 14841 10421 14875 10455
rect 2237 10217 2271 10251
rect 2605 10217 2639 10251
rect 3985 10217 4019 10251
rect 7665 10217 7699 10251
rect 10149 10217 10183 10251
rect 17325 10217 17359 10251
rect 4813 10149 4847 10183
rect 7481 10149 7515 10183
rect 17693 10149 17727 10183
rect 3801 10081 3835 10115
rect 4537 10081 4571 10115
rect 5273 10081 5307 10115
rect 5457 10081 5491 10115
rect 6285 10081 6319 10115
rect 7113 10081 7147 10115
rect 8217 10081 8251 10115
rect 9505 10081 9539 10115
rect 9965 10081 9999 10115
rect 10517 10081 10551 10115
rect 10609 10081 10643 10115
rect 11713 10081 11747 10115
rect 12725 10081 12759 10115
rect 13461 10081 13495 10115
rect 14657 10081 14691 10115
rect 15485 10081 15519 10115
rect 16313 10081 16347 10115
rect 16589 10081 16623 10115
rect 17049 10081 17083 10115
rect 2053 10013 2087 10047
rect 4353 10013 4387 10047
rect 5181 10013 5215 10047
rect 6009 10013 6043 10047
rect 6837 10013 6871 10047
rect 8493 10013 8527 10047
rect 9413 10013 9447 10047
rect 10701 10013 10735 10047
rect 13277 10013 13311 10047
rect 14473 10013 14507 10047
rect 17509 10013 17543 10047
rect 17877 10013 17911 10047
rect 18245 10013 18279 10047
rect 4445 9945 4479 9979
rect 6101 9945 6135 9979
rect 8033 9945 8067 9979
rect 11529 9945 11563 9979
rect 12449 9945 12483 9979
rect 16221 9945 16255 9979
rect 1869 9877 1903 9911
rect 5641 9877 5675 9911
rect 6469 9877 6503 9911
rect 6929 9877 6963 9911
rect 7389 9877 7423 9911
rect 8125 9877 8159 9911
rect 8677 9877 8711 9911
rect 8953 9877 8987 9911
rect 9321 9877 9355 9911
rect 11069 9877 11103 9911
rect 11161 9877 11195 9911
rect 11621 9877 11655 9911
rect 12081 9877 12115 9911
rect 12541 9877 12575 9911
rect 12909 9877 12943 9911
rect 13369 9877 13403 9911
rect 14105 9877 14139 9911
rect 14565 9877 14599 9911
rect 14933 9877 14967 9911
rect 15301 9877 15335 9911
rect 15393 9877 15427 9911
rect 15761 9877 15795 9911
rect 16129 9877 16163 9911
rect 16865 9877 16899 9911
rect 18061 9877 18095 9911
rect 18429 9877 18463 9911
rect 2237 9673 2271 9707
rect 4353 9673 4387 9707
rect 5641 9673 5675 9707
rect 6101 9673 6135 9707
rect 6837 9673 6871 9707
rect 7941 9673 7975 9707
rect 8309 9673 8343 9707
rect 9873 9673 9907 9707
rect 11161 9673 11195 9707
rect 11897 9673 11931 9707
rect 12357 9673 12391 9707
rect 13185 9673 13219 9707
rect 13553 9673 13587 9707
rect 14841 9673 14875 9707
rect 15209 9673 15243 9707
rect 16681 9673 16715 9707
rect 17877 9673 17911 9707
rect 18337 9673 18371 9707
rect 3525 9605 3559 9639
rect 6745 9605 6779 9639
rect 9137 9605 9171 9639
rect 11345 9605 11379 9639
rect 11989 9605 12023 9639
rect 14381 9605 14415 9639
rect 15945 9605 15979 9639
rect 16037 9605 16071 9639
rect 17049 9605 17083 9639
rect 2789 9537 2823 9571
rect 4445 9537 4479 9571
rect 5089 9537 5123 9571
rect 5549 9537 5583 9571
rect 7665 9537 7699 9571
rect 7849 9537 7883 9571
rect 8401 9537 8435 9571
rect 9965 9537 9999 9571
rect 10793 9537 10827 9571
rect 12725 9537 12759 9571
rect 12817 9537 12851 9571
rect 1961 9469 1995 9503
rect 2145 9469 2179 9503
rect 3617 9469 3651 9503
rect 3801 9469 3835 9503
rect 4537 9469 4571 9503
rect 5825 9469 5859 9503
rect 6929 9469 6963 9503
rect 8585 9469 8619 9503
rect 9229 9469 9263 9503
rect 9413 9469 9447 9503
rect 9781 9469 9815 9503
rect 10609 9469 10643 9503
rect 10701 9469 10735 9503
rect 12081 9469 12115 9503
rect 12909 9469 12943 9503
rect 13645 9469 13679 9503
rect 13737 9469 13771 9503
rect 14105 9469 14139 9503
rect 14289 9469 14323 9503
rect 15301 9469 15335 9503
rect 15393 9469 15427 9503
rect 15761 9469 15795 9503
rect 17141 9469 17175 9503
rect 17325 9469 17359 9503
rect 17969 9469 18003 9503
rect 18061 9469 18095 9503
rect 2605 9401 2639 9435
rect 2973 9401 3007 9435
rect 3985 9401 4019 9435
rect 4813 9401 4847 9435
rect 7389 9401 7423 9435
rect 10333 9401 10367 9435
rect 11529 9401 11563 9435
rect 14749 9401 14783 9435
rect 3157 9333 3191 9367
rect 5181 9333 5215 9367
rect 6377 9333 6411 9367
rect 7205 9333 7239 9367
rect 8769 9333 8803 9367
rect 16405 9333 16439 9367
rect 17509 9333 17543 9367
rect 1961 9129 1995 9163
rect 3157 9129 3191 9163
rect 8953 9129 8987 9163
rect 10517 9129 10551 9163
rect 11621 9129 11655 9163
rect 14197 9129 14231 9163
rect 15393 9129 15427 9163
rect 17049 9129 17083 9163
rect 17417 9129 17451 9163
rect 7941 9061 7975 9095
rect 9873 9061 9907 9095
rect 12449 9061 12483 9095
rect 14381 9061 14415 9095
rect 2421 8993 2455 9027
rect 2605 8993 2639 9027
rect 4445 8993 4479 9027
rect 5181 8993 5215 9027
rect 5549 8993 5583 9027
rect 8125 8993 8159 9027
rect 8309 8993 8343 9027
rect 9505 8993 9539 9027
rect 11161 8993 11195 9027
rect 11345 8993 11379 9027
rect 11989 8993 12023 9027
rect 14657 8993 14691 9027
rect 15853 8993 15887 9027
rect 15945 8993 15979 9027
rect 16773 8993 16807 9027
rect 17969 8993 18003 9027
rect 1501 8925 1535 8959
rect 1869 8925 1903 8959
rect 3617 8925 3651 8959
rect 4261 8925 4295 8959
rect 6561 8925 6595 8959
rect 6817 8925 6851 8959
rect 8401 8925 8435 8959
rect 10149 8925 10183 8959
rect 11069 8925 11103 8959
rect 14933 8925 14967 8959
rect 16589 8925 16623 8959
rect 17785 8925 17819 8959
rect 18245 8925 18279 8959
rect 3433 8857 3467 8891
rect 4169 8857 4203 8891
rect 5825 8857 5859 8891
rect 9413 8857 9447 8891
rect 13737 8857 13771 8891
rect 17233 8857 17267 8891
rect 1685 8789 1719 8823
rect 2329 8789 2363 8823
rect 2881 8789 2915 8823
rect 3801 8789 3835 8823
rect 4629 8789 4663 8823
rect 4997 8789 5031 8823
rect 5089 8789 5123 8823
rect 5733 8789 5767 8823
rect 6193 8789 6227 8823
rect 6469 8789 6503 8823
rect 8769 8789 8803 8823
rect 9321 8789 9355 8823
rect 10057 8789 10091 8823
rect 10701 8789 10735 8823
rect 13001 8789 13035 8823
rect 13277 8789 13311 8823
rect 13921 8789 13955 8823
rect 14841 8789 14875 8823
rect 15301 8789 15335 8823
rect 15761 8789 15795 8823
rect 16221 8789 16255 8823
rect 16681 8789 16715 8823
rect 17877 8789 17911 8823
rect 18429 8789 18463 8823
rect 2053 8585 2087 8619
rect 3249 8585 3283 8619
rect 4445 8585 4479 8619
rect 6377 8585 6411 8619
rect 6837 8585 6871 8619
rect 8585 8585 8619 8619
rect 10517 8585 10551 8619
rect 11621 8585 11655 8619
rect 14841 8585 14875 8619
rect 16681 8585 16715 8619
rect 1685 8517 1719 8551
rect 2513 8517 2547 8551
rect 3341 8517 3375 8551
rect 7450 8517 7484 8551
rect 8861 8517 8895 8551
rect 9382 8517 9416 8551
rect 12756 8517 12790 8551
rect 17693 8517 17727 8551
rect 1869 8449 1903 8483
rect 2421 8449 2455 8483
rect 4353 8449 4387 8483
rect 4813 8449 4847 8483
rect 5080 8449 5114 8483
rect 6745 8449 6779 8483
rect 7205 8449 7239 8483
rect 13728 8449 13762 8483
rect 16046 8449 16080 8483
rect 17049 8449 17083 8483
rect 17877 8449 17911 8483
rect 18245 8449 18279 8483
rect 2697 8381 2731 8415
rect 3433 8381 3467 8415
rect 3893 8381 3927 8415
rect 4629 8381 4663 8415
rect 6929 8381 6963 8415
rect 9137 8381 9171 8415
rect 13001 8381 13035 8415
rect 13369 8381 13403 8415
rect 13461 8381 13495 8415
rect 16313 8381 16347 8415
rect 16405 8381 16439 8415
rect 17141 8381 17175 8415
rect 17233 8381 17267 8415
rect 2881 8313 2915 8347
rect 3985 8313 4019 8347
rect 6193 8313 6227 8347
rect 14933 8313 14967 8347
rect 17509 8313 17543 8347
rect 18061 8313 18095 8347
rect 18429 8313 18463 8347
rect 8953 8245 8987 8279
rect 10701 8245 10735 8279
rect 11253 8245 11287 8279
rect 2237 8041 2271 8075
rect 2605 8041 2639 8075
rect 4721 8041 4755 8075
rect 5549 8041 5583 8075
rect 7297 8041 7331 8075
rect 9597 8041 9631 8075
rect 12725 8041 12759 8075
rect 15577 8041 15611 8075
rect 17049 8041 17083 8075
rect 18245 8041 18279 8075
rect 2697 7973 2731 8007
rect 18061 7973 18095 8007
rect 1685 7905 1719 7939
rect 3525 7905 3559 7939
rect 4169 7905 4203 7939
rect 4997 7905 5031 7939
rect 5089 7905 5123 7939
rect 17601 7905 17635 7939
rect 1501 7837 1535 7871
rect 2053 7837 2087 7871
rect 2421 7837 2455 7871
rect 4353 7837 4387 7871
rect 5917 7837 5951 7871
rect 6184 7837 6218 7871
rect 8769 7837 8803 7871
rect 8953 7837 8987 7871
rect 10710 7837 10744 7871
rect 10977 7837 11011 7871
rect 11161 7837 11195 7871
rect 11345 7837 11379 7871
rect 11601 7837 11635 7871
rect 13829 7837 13863 7871
rect 15485 7837 15519 7871
rect 16957 7837 16991 7871
rect 17417 7837 17451 7871
rect 17877 7837 17911 7871
rect 5181 7769 5215 7803
rect 8524 7769 8558 7803
rect 15218 7769 15252 7803
rect 16712 7769 16746 7803
rect 17509 7769 17543 7803
rect 18429 7769 18463 7803
rect 1869 7701 1903 7735
rect 2881 7701 2915 7735
rect 3249 7701 3283 7735
rect 3341 7701 3375 7735
rect 3801 7701 3835 7735
rect 4261 7701 4295 7735
rect 5825 7701 5859 7735
rect 7389 7701 7423 7735
rect 13645 7701 13679 7735
rect 14105 7701 14139 7735
rect 2973 7497 3007 7531
rect 3341 7497 3375 7531
rect 3893 7497 3927 7531
rect 4629 7497 4663 7531
rect 5089 7497 5123 7531
rect 6469 7497 6503 7531
rect 7941 7497 7975 7531
rect 12909 7497 12943 7531
rect 13369 7497 13403 7531
rect 13553 7497 13587 7531
rect 13737 7497 13771 7531
rect 15301 7497 15335 7531
rect 15485 7497 15519 7531
rect 15577 7497 15611 7531
rect 16221 7497 16255 7531
rect 16681 7497 16715 7531
rect 17141 7497 17175 7531
rect 17877 7497 17911 7531
rect 4537 7429 4571 7463
rect 4997 7429 5031 7463
rect 9404 7429 9438 7463
rect 11774 7429 11808 7463
rect 1685 7361 1719 7395
rect 2145 7361 2179 7395
rect 3801 7361 3835 7395
rect 5641 7361 5675 7395
rect 6828 7361 6862 7395
rect 11529 7361 11563 7395
rect 14850 7361 14884 7395
rect 15117 7361 15151 7395
rect 16129 7361 16163 7395
rect 17049 7361 17083 7395
rect 17969 7361 18003 7395
rect 1961 7293 1995 7327
rect 2053 7293 2087 7327
rect 2789 7293 2823 7327
rect 2881 7293 2915 7327
rect 3985 7293 4019 7327
rect 5273 7293 5307 7327
rect 6561 7293 6595 7327
rect 9137 7293 9171 7327
rect 11345 7293 11379 7327
rect 16313 7293 16347 7327
rect 17325 7293 17359 7327
rect 18061 7293 18095 7327
rect 18337 7293 18371 7327
rect 1501 7225 1535 7259
rect 8033 7225 8067 7259
rect 8217 7225 8251 7259
rect 10517 7225 10551 7259
rect 2513 7157 2547 7191
rect 3433 7157 3467 7191
rect 4353 7157 4387 7191
rect 5549 7157 5583 7191
rect 5917 7157 5951 7191
rect 10701 7157 10735 7191
rect 10977 7157 11011 7191
rect 11069 7157 11103 7191
rect 15761 7157 15795 7191
rect 17509 7157 17543 7191
rect 1685 6953 1719 6987
rect 2605 6953 2639 6987
rect 3893 6953 3927 6987
rect 7297 6953 7331 6987
rect 9965 6953 9999 6987
rect 11437 6953 11471 6987
rect 13829 6953 13863 6987
rect 18061 6953 18095 6987
rect 5825 6885 5859 6919
rect 7389 6885 7423 6919
rect 13737 6885 13771 6919
rect 2145 6817 2179 6851
rect 2973 6817 3007 6851
rect 3157 6817 3191 6851
rect 13093 6817 13127 6851
rect 14105 6817 14139 6851
rect 17601 6817 17635 6851
rect 1501 6749 1535 6783
rect 2053 6749 2087 6783
rect 3249 6749 3283 6783
rect 4077 6749 4111 6783
rect 4261 6749 4295 6783
rect 4445 6749 4479 6783
rect 5917 6749 5951 6783
rect 8769 6749 8803 6783
rect 11078 6749 11112 6783
rect 11345 6749 11379 6783
rect 12817 6749 12851 6783
rect 14361 6749 14395 6783
rect 16957 6749 16991 6783
rect 17509 6749 17543 6783
rect 17877 6749 17911 6783
rect 18245 6749 18279 6783
rect 2513 6681 2547 6715
rect 4712 6681 4746 6715
rect 6184 6681 6218 6715
rect 8524 6681 8558 6715
rect 12550 6681 12584 6715
rect 13369 6681 13403 6715
rect 13553 6681 13587 6715
rect 16712 6681 16746 6715
rect 1869 6613 1903 6647
rect 3617 6613 3651 6647
rect 9045 6613 9079 6647
rect 9137 6613 9171 6647
rect 13001 6613 13035 6647
rect 15485 6613 15519 6647
rect 15577 6613 15611 6647
rect 17049 6613 17083 6647
rect 17417 6613 17451 6647
rect 18429 6613 18463 6647
rect 2789 6409 2823 6443
rect 4353 6409 4387 6443
rect 4445 6409 4479 6443
rect 10609 6409 10643 6443
rect 10793 6409 10827 6443
rect 10977 6409 11011 6443
rect 11345 6409 11379 6443
rect 11621 6409 11655 6443
rect 11989 6409 12023 6443
rect 12173 6409 12207 6443
rect 13369 6409 13403 6443
rect 14933 6409 14967 6443
rect 16405 6409 16439 6443
rect 17233 6409 17267 6443
rect 17693 6409 17727 6443
rect 3801 6341 3835 6375
rect 9496 6341 9530 6375
rect 12633 6341 12667 6375
rect 14596 6341 14630 6375
rect 17785 6341 17819 6375
rect 1685 6273 1719 6307
rect 2053 6273 2087 6307
rect 2421 6273 2455 6307
rect 3157 6273 3191 6307
rect 3617 6273 3651 6307
rect 5080 6273 5114 6307
rect 7369 6273 7403 6307
rect 8677 6273 8711 6307
rect 9229 6273 9263 6307
rect 14841 6273 14875 6307
rect 16046 6273 16080 6307
rect 16313 6273 16347 6307
rect 18153 6273 18187 6307
rect 18337 6273 18371 6307
rect 3249 6205 3283 6239
rect 3433 6205 3467 6239
rect 4629 6205 4663 6239
rect 4813 6205 4847 6239
rect 7113 6205 7147 6239
rect 16773 6205 16807 6239
rect 17877 6205 17911 6239
rect 2237 6137 2271 6171
rect 6193 6137 6227 6171
rect 8493 6137 8527 6171
rect 13461 6137 13495 6171
rect 1501 6069 1535 6103
rect 1869 6069 1903 6103
rect 2697 6069 2731 6103
rect 3985 6069 4019 6103
rect 6377 6069 6411 6103
rect 6653 6069 6687 6103
rect 11713 6069 11747 6103
rect 12449 6069 12483 6103
rect 12817 6069 12851 6103
rect 13001 6069 13035 6103
rect 13185 6069 13219 6103
rect 16957 6069 16991 6103
rect 17325 6069 17359 6103
rect 1501 5865 1535 5899
rect 2329 5865 2363 5899
rect 3157 5865 3191 5899
rect 3617 5865 3651 5899
rect 11989 5865 12023 5899
rect 12081 5865 12115 5899
rect 13737 5865 13771 5899
rect 15577 5865 15611 5899
rect 15761 5865 15795 5899
rect 15945 5865 15979 5899
rect 6009 5797 6043 5831
rect 6101 5797 6135 5831
rect 2605 5729 2639 5763
rect 2697 5729 2731 5763
rect 3985 5729 4019 5763
rect 4629 5729 4663 5763
rect 16589 5729 16623 5763
rect 16773 5729 16807 5763
rect 17509 5729 17543 5763
rect 18337 5729 18371 5763
rect 2053 5661 2087 5695
rect 3341 5661 3375 5695
rect 4077 5661 4111 5695
rect 7481 5661 7515 5695
rect 7573 5661 7607 5695
rect 7757 5661 7791 5695
rect 8125 5661 8159 5695
rect 9137 5661 9171 5695
rect 10609 5661 10643 5695
rect 10876 5661 10910 5695
rect 13194 5661 13228 5695
rect 13461 5661 13495 5695
rect 13921 5661 13955 5695
rect 14105 5661 14139 5695
rect 16497 5661 16531 5695
rect 2789 5593 2823 5627
rect 4169 5593 4203 5627
rect 4896 5593 4930 5627
rect 7214 5593 7248 5627
rect 9382 5593 9416 5627
rect 14372 5593 14406 5627
rect 1593 5525 1627 5559
rect 1869 5525 1903 5559
rect 4537 5525 4571 5559
rect 10517 5525 10551 5559
rect 15485 5525 15519 5559
rect 16129 5525 16163 5559
rect 16957 5525 16991 5559
rect 17325 5525 17359 5559
rect 17417 5525 17451 5559
rect 17785 5525 17819 5559
rect 18153 5525 18187 5559
rect 18245 5525 18279 5559
rect 2605 5321 2639 5355
rect 3985 5321 4019 5355
rect 4077 5321 4111 5355
rect 4445 5321 4479 5355
rect 6101 5321 6135 5355
rect 6377 5321 6411 5355
rect 15945 5321 15979 5355
rect 16405 5321 16439 5355
rect 17417 5321 17451 5355
rect 18245 5321 18279 5355
rect 18337 5321 18371 5355
rect 9597 5253 9631 5287
rect 9781 5253 9815 5287
rect 11796 5253 11830 5287
rect 14114 5253 14148 5287
rect 17785 5253 17819 5287
rect 1685 5185 1719 5219
rect 2053 5185 2087 5219
rect 2421 5185 2455 5219
rect 3157 5185 3191 5219
rect 4813 5185 4847 5219
rect 5641 5185 5675 5219
rect 6653 5185 6687 5219
rect 6920 5185 6954 5219
rect 8125 5185 8159 5219
rect 8392 5185 8426 5219
rect 9965 5185 9999 5219
rect 10221 5185 10255 5219
rect 11529 5185 11563 5219
rect 14381 5185 14415 5219
rect 14473 5185 14507 5219
rect 14740 5185 14774 5219
rect 17049 5185 17083 5219
rect 17877 5185 17911 5219
rect 3249 5117 3283 5151
rect 3433 5117 3467 5151
rect 4261 5117 4295 5151
rect 4905 5117 4939 5151
rect 4997 5117 5031 5151
rect 5733 5117 5767 5151
rect 5825 5117 5859 5151
rect 16773 5117 16807 5151
rect 16957 5117 16991 5151
rect 17601 5117 17635 5151
rect 5273 5049 5307 5083
rect 8033 5049 8067 5083
rect 9505 5049 9539 5083
rect 12909 5049 12943 5083
rect 15853 5049 15887 5083
rect 1501 4981 1535 5015
rect 1869 4981 1903 5015
rect 2237 4981 2271 5015
rect 2789 4981 2823 5015
rect 3617 4981 3651 5015
rect 11345 4981 11379 5015
rect 13001 4981 13035 5015
rect 16313 4981 16347 5015
rect 1777 4777 1811 4811
rect 2881 4777 2915 4811
rect 4353 4777 4387 4811
rect 5825 4777 5859 4811
rect 9781 4777 9815 4811
rect 9965 4777 9999 4811
rect 13277 4777 13311 4811
rect 13461 4777 13495 4811
rect 13645 4777 13679 4811
rect 13829 4777 13863 4811
rect 14105 4777 14139 4811
rect 17969 4777 18003 4811
rect 18429 4777 18463 4811
rect 1593 4709 1627 4743
rect 5917 4709 5951 4743
rect 8769 4709 8803 4743
rect 10057 4709 10091 4743
rect 2145 4641 2179 4675
rect 2329 4641 2363 4675
rect 3341 4641 3375 4675
rect 3525 4641 3559 4675
rect 15485 4641 15519 4675
rect 16129 4641 16163 4675
rect 16957 4641 16991 4675
rect 17325 4641 17359 4675
rect 1961 4573 1995 4607
rect 4077 4573 4111 4607
rect 4445 4573 4479 4607
rect 7297 4573 7331 4607
rect 7389 4573 7423 4607
rect 7656 4573 7690 4607
rect 9413 4573 9447 4607
rect 9597 4573 9631 4607
rect 11437 4573 11471 4607
rect 11713 4573 11747 4607
rect 15945 4573 15979 4607
rect 17601 4573 17635 4607
rect 18061 4573 18095 4607
rect 2421 4505 2455 4539
rect 3249 4505 3283 4539
rect 4712 4505 4746 4539
rect 7030 4505 7064 4539
rect 9137 4505 9171 4539
rect 11170 4505 11204 4539
rect 11980 4505 12014 4539
rect 15218 4505 15252 4539
rect 16773 4505 16807 4539
rect 2789 4437 2823 4471
rect 3893 4437 3927 4471
rect 11621 4437 11655 4471
rect 13093 4437 13127 4471
rect 15577 4437 15611 4471
rect 16037 4437 16071 4471
rect 16405 4437 16439 4471
rect 16865 4437 16899 4471
rect 17509 4437 17543 4471
rect 18245 4437 18279 4471
rect 2697 4233 2731 4267
rect 2881 4233 2915 4267
rect 3065 4233 3099 4267
rect 4353 4233 4387 4267
rect 8401 4233 8435 4267
rect 11621 4233 11655 4267
rect 11805 4233 11839 4267
rect 11989 4233 12023 4267
rect 13645 4233 13679 4267
rect 16037 4233 16071 4267
rect 17141 4233 17175 4267
rect 17509 4233 17543 4267
rect 18153 4233 18187 4267
rect 1501 4165 1535 4199
rect 1685 4165 1719 4199
rect 3433 4165 3467 4199
rect 3525 4165 3559 4199
rect 9536 4165 9570 4199
rect 15945 4165 15979 4199
rect 2053 4097 2087 4131
rect 2421 4097 2455 4131
rect 4261 4097 4295 4131
rect 5080 4097 5114 4131
rect 6377 4097 6411 4131
rect 8042 4097 8076 4131
rect 9781 4097 9815 4131
rect 9873 4097 9907 4131
rect 10129 4097 10163 4131
rect 13286 4097 13320 4131
rect 13553 4097 13587 4131
rect 14105 4097 14139 4131
rect 14361 4097 14395 4131
rect 16405 4097 16439 4131
rect 16773 4097 16807 4131
rect 17969 4097 18003 4131
rect 18429 4097 18463 4131
rect 3341 4029 3375 4063
rect 4169 4029 4203 4063
rect 4813 4029 4847 4063
rect 6653 4029 6687 4063
rect 8309 4029 8343 4063
rect 13829 4029 13863 4063
rect 16129 4029 16163 4063
rect 17601 4029 17635 4063
rect 17693 4029 17727 4063
rect 6929 3961 6963 3995
rect 11253 3961 11287 3995
rect 16957 3961 16991 3995
rect 1869 3893 1903 3927
rect 2237 3893 2271 3927
rect 3893 3893 3927 3927
rect 4721 3893 4755 3927
rect 6193 3893 6227 3927
rect 12173 3893 12207 3927
rect 15485 3893 15519 3927
rect 15577 3893 15611 3927
rect 1501 3689 1535 3723
rect 1685 3689 1719 3723
rect 3893 3689 3927 3723
rect 4813 3689 4847 3723
rect 4997 3689 5031 3723
rect 11897 3689 11931 3723
rect 13461 3689 13495 3723
rect 13645 3689 13679 3723
rect 13829 3689 13863 3723
rect 14105 3689 14139 3723
rect 15577 3689 15611 3723
rect 17509 3689 17543 3723
rect 18337 3689 18371 3723
rect 1777 3621 1811 3655
rect 2053 3621 2087 3655
rect 2881 3621 2915 3655
rect 3985 3621 4019 3655
rect 5181 3621 5215 3655
rect 9045 3621 9079 3655
rect 2237 3553 2271 3587
rect 3341 3553 3375 3587
rect 3433 3553 3467 3587
rect 4629 3553 4663 3587
rect 13369 3553 13403 3587
rect 15485 3553 15519 3587
rect 18061 3553 18095 3587
rect 2789 3485 2823 3519
rect 3249 3485 3283 3519
rect 6561 3485 6595 3519
rect 8033 3485 8067 3519
rect 8125 3485 8159 3519
rect 8309 3485 8343 3519
rect 10425 3485 10459 3519
rect 10517 3485 10551 3519
rect 13113 3485 13147 3519
rect 16957 3485 16991 3519
rect 17141 3485 17175 3519
rect 2513 3417 2547 3451
rect 4445 3417 4479 3451
rect 6316 3417 6350 3451
rect 7788 3417 7822 3451
rect 8585 3417 8619 3451
rect 10158 3417 10192 3451
rect 10762 3417 10796 3451
rect 15240 3417 15274 3451
rect 16712 3417 16746 3451
rect 17877 3417 17911 3451
rect 4353 3349 4387 3383
rect 6653 3349 6687 3383
rect 11989 3349 12023 3383
rect 17325 3349 17359 3383
rect 17969 3349 18003 3383
rect 4261 3145 4295 3179
rect 4353 3145 4387 3179
rect 4721 3145 4755 3179
rect 9873 3145 9907 3179
rect 11529 3145 11563 3179
rect 14473 3145 14507 3179
rect 16957 3145 16991 3179
rect 17417 3145 17451 3179
rect 17785 3145 17819 3179
rect 18153 3145 18187 3179
rect 3065 3077 3099 3111
rect 8760 3077 8794 3111
rect 15586 3077 15620 3111
rect 1685 3009 1719 3043
rect 2237 3009 2271 3043
rect 2789 3009 2823 3043
rect 3341 3009 3375 3043
rect 3893 3009 3927 3043
rect 5926 3009 5960 3043
rect 7490 3009 7524 3043
rect 7757 3009 7791 3043
rect 8401 3009 8435 3043
rect 11078 3009 11112 3043
rect 11345 3009 11379 3043
rect 12642 3009 12676 3043
rect 12909 3009 12943 3043
rect 13001 3009 13035 3043
rect 13268 3009 13302 3043
rect 15853 3009 15887 3043
rect 15945 3009 15979 3043
rect 17325 3009 17359 3043
rect 2053 2941 2087 2975
rect 2605 2941 2639 2975
rect 3709 2941 3743 2975
rect 4169 2941 4203 2975
rect 6193 2941 6227 2975
rect 8217 2941 8251 2975
rect 8493 2941 8527 2975
rect 16129 2941 16163 2975
rect 17601 2941 17635 2975
rect 18245 2941 18279 2975
rect 18337 2941 18371 2975
rect 4813 2873 4847 2907
rect 14381 2873 14415 2907
rect 16865 2873 16899 2907
rect 1501 2805 1535 2839
rect 6377 2805 6411 2839
rect 9965 2805 9999 2839
rect 1501 2601 1535 2635
rect 2697 2601 2731 2635
rect 3065 2601 3099 2635
rect 6193 2601 6227 2635
rect 7021 2601 7055 2635
rect 8493 2601 8527 2635
rect 8677 2601 8711 2635
rect 8953 2601 8987 2635
rect 9321 2601 9355 2635
rect 11621 2601 11655 2635
rect 11713 2601 11747 2635
rect 14749 2601 14783 2635
rect 14841 2601 14875 2635
rect 15025 2601 15059 2635
rect 15853 2601 15887 2635
rect 16129 2601 16163 2635
rect 17049 2601 17083 2635
rect 18061 2601 18095 2635
rect 2329 2533 2363 2567
rect 2881 2533 2915 2567
rect 5089 2533 5123 2567
rect 16313 2533 16347 2567
rect 16773 2533 16807 2567
rect 1961 2465 1995 2499
rect 4077 2465 4111 2499
rect 4537 2465 4571 2499
rect 5365 2465 5399 2499
rect 5457 2465 5491 2499
rect 8401 2465 8435 2499
rect 9873 2465 9907 2499
rect 10241 2465 10275 2499
rect 11161 2465 11195 2499
rect 13921 2465 13955 2499
rect 2145 2397 2179 2431
rect 2513 2397 2547 2431
rect 3617 2397 3651 2431
rect 3801 2397 3835 2431
rect 4629 2397 4663 2431
rect 4721 2397 4755 2431
rect 5549 2397 5583 2431
rect 6469 2397 6503 2431
rect 9137 2397 9171 2431
rect 10333 2397 10367 2431
rect 12357 2397 12391 2431
rect 13654 2397 13688 2431
rect 14105 2397 14139 2431
rect 15485 2397 15519 2431
rect 15761 2397 15795 2431
rect 17141 2397 17175 2431
rect 17509 2397 17543 2431
rect 17877 2397 17911 2431
rect 18245 2397 18279 2431
rect 3341 2329 3375 2363
rect 6745 2329 6779 2363
rect 8156 2329 8190 2363
rect 9689 2329 9723 2363
rect 12081 2329 12115 2363
rect 14381 2329 14415 2363
rect 5917 2261 5951 2295
rect 9781 2261 9815 2295
rect 12541 2261 12575 2295
rect 16497 2261 16531 2295
rect 17325 2261 17359 2295
rect 17693 2261 17727 2295
rect 18429 2261 18463 2295
<< metal1 >>
rect 6270 15308 6276 15360
rect 6328 15348 6334 15360
rect 15194 15348 15200 15360
rect 6328 15320 15200 15348
rect 6328 15308 6334 15320
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 3418 15240 3424 15292
rect 3476 15280 3482 15292
rect 11238 15280 11244 15292
rect 3476 15252 11244 15280
rect 3476 15240 3482 15252
rect 11238 15240 11244 15252
rect 11296 15240 11302 15292
rect 3050 15172 3056 15224
rect 3108 15212 3114 15224
rect 3970 15212 3976 15224
rect 3108 15184 3976 15212
rect 3108 15172 3114 15184
rect 3970 15172 3976 15184
rect 4028 15212 4034 15224
rect 7006 15212 7012 15224
rect 4028 15184 7012 15212
rect 4028 15172 4034 15184
rect 7006 15172 7012 15184
rect 7064 15172 7070 15224
rect 13538 15172 13544 15224
rect 13596 15212 13602 15224
rect 15286 15212 15292 15224
rect 13596 15184 15292 15212
rect 13596 15172 13602 15184
rect 15286 15172 15292 15184
rect 15344 15172 15350 15224
rect 1104 14714 18860 14736
rect 1104 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 3302 14714
rect 3354 14662 3366 14714
rect 3418 14662 3430 14714
rect 3482 14662 7622 14714
rect 7674 14662 7686 14714
rect 7738 14662 7750 14714
rect 7802 14662 7814 14714
rect 7866 14662 7878 14714
rect 7930 14662 12070 14714
rect 12122 14662 12134 14714
rect 12186 14662 12198 14714
rect 12250 14662 12262 14714
rect 12314 14662 12326 14714
rect 12378 14662 16518 14714
rect 16570 14662 16582 14714
rect 16634 14662 16646 14714
rect 16698 14662 16710 14714
rect 16762 14662 16774 14714
rect 16826 14662 18860 14714
rect 1104 14640 18860 14662
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 5169 14603 5227 14609
rect 5169 14600 5181 14603
rect 4212 14572 5181 14600
rect 4212 14560 4218 14572
rect 5169 14569 5181 14572
rect 5215 14600 5227 14603
rect 5718 14600 5724 14612
rect 5215 14572 5724 14600
rect 5215 14569 5227 14572
rect 5169 14563 5227 14569
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 9766 14492 9772 14544
rect 9824 14532 9830 14544
rect 15286 14532 15292 14544
rect 9824 14504 15292 14532
rect 9824 14492 9830 14504
rect 15286 14492 15292 14504
rect 15344 14492 15350 14544
rect 1118 14424 1124 14476
rect 1176 14464 1182 14476
rect 10318 14464 10324 14476
rect 1176 14436 10324 14464
rect 1176 14424 1182 14436
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 14366 14424 14372 14476
rect 14424 14464 14430 14476
rect 15102 14464 15108 14476
rect 14424 14436 15108 14464
rect 14424 14424 14430 14436
rect 15102 14424 15108 14436
rect 15160 14424 15166 14476
rect 3418 14356 3424 14408
rect 3476 14396 3482 14408
rect 7374 14396 7380 14408
rect 3476 14368 7380 14396
rect 3476 14356 3482 14368
rect 7374 14356 7380 14368
rect 7432 14356 7438 14408
rect 10594 14356 10600 14408
rect 10652 14396 10658 14408
rect 15194 14396 15200 14408
rect 10652 14368 15200 14396
rect 10652 14356 10658 14368
rect 15194 14356 15200 14368
rect 15252 14356 15258 14408
rect 16666 14396 16672 14408
rect 16546 14368 16672 14396
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 16546 14328 16574 14368
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 3660 14300 16574 14328
rect 3660 14288 3666 14300
rect 4982 14260 4988 14272
rect 4943 14232 4988 14260
rect 4982 14220 4988 14232
rect 5040 14220 5046 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 14734 14260 14740 14272
rect 5592 14232 14740 14260
rect 5592 14220 5598 14232
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 1104 14170 18860 14192
rect 1104 14118 5398 14170
rect 5450 14118 5462 14170
rect 5514 14118 5526 14170
rect 5578 14118 5590 14170
rect 5642 14118 5654 14170
rect 5706 14118 9846 14170
rect 9898 14118 9910 14170
rect 9962 14118 9974 14170
rect 10026 14118 10038 14170
rect 10090 14118 10102 14170
rect 10154 14118 14294 14170
rect 14346 14118 14358 14170
rect 14410 14118 14422 14170
rect 14474 14118 14486 14170
rect 14538 14118 14550 14170
rect 14602 14118 18860 14170
rect 1104 14096 18860 14118
rect 3602 14016 3608 14068
rect 3660 14056 3666 14068
rect 4157 14059 4215 14065
rect 4157 14056 4169 14059
rect 3660 14028 4169 14056
rect 3660 14016 3666 14028
rect 4157 14025 4169 14028
rect 4203 14025 4215 14059
rect 4157 14019 4215 14025
rect 4525 14059 4583 14065
rect 4525 14025 4537 14059
rect 4571 14056 4583 14059
rect 4985 14059 5043 14065
rect 4985 14056 4997 14059
rect 4571 14028 4997 14056
rect 4571 14025 4583 14028
rect 4525 14019 4583 14025
rect 4985 14025 4997 14028
rect 5031 14025 5043 14059
rect 4985 14019 5043 14025
rect 5074 14016 5080 14068
rect 5132 14056 5138 14068
rect 5445 14059 5503 14065
rect 5445 14056 5457 14059
rect 5132 14028 5457 14056
rect 5132 14016 5138 14028
rect 5445 14025 5457 14028
rect 5491 14056 5503 14059
rect 5491 14028 6040 14056
rect 5491 14025 5503 14028
rect 5445 14019 5503 14025
rect 3510 13948 3516 14000
rect 3568 13988 3574 14000
rect 5902 13988 5908 14000
rect 3568 13960 5908 13988
rect 3568 13948 3574 13960
rect 5902 13948 5908 13960
rect 5960 13948 5966 14000
rect 4246 13880 4252 13932
rect 4304 13920 4310 13932
rect 5353 13923 5411 13929
rect 4304 13892 5120 13920
rect 4304 13880 4310 13892
rect 4614 13852 4620 13864
rect 4575 13824 4620 13852
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 4709 13855 4767 13861
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 4982 13852 4988 13864
rect 4755 13824 4988 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 4338 13744 4344 13796
rect 4396 13784 4402 13796
rect 4724 13784 4752 13815
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 5092 13852 5120 13892
rect 5353 13889 5365 13923
rect 5399 13920 5411 13923
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5399 13892 5825 13920
rect 5399 13889 5411 13892
rect 5353 13883 5411 13889
rect 5813 13889 5825 13892
rect 5859 13889 5871 13923
rect 6012 13920 6040 14028
rect 6454 14016 6460 14068
rect 6512 14056 6518 14068
rect 9766 14056 9772 14068
rect 6512 14028 9772 14056
rect 6512 14016 6518 14028
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10318 14056 10324 14068
rect 10279 14028 10324 14056
rect 10318 14016 10324 14028
rect 10376 14056 10382 14068
rect 14645 14059 14703 14065
rect 14645 14056 14657 14059
rect 10376 14028 10548 14056
rect 10376 14016 10382 14028
rect 6086 13948 6092 14000
rect 6144 13988 6150 14000
rect 9674 13988 9680 14000
rect 6144 13960 9680 13988
rect 6144 13948 6150 13960
rect 9674 13948 9680 13960
rect 9732 13948 9738 14000
rect 10410 13920 10416 13932
rect 6012 13892 6684 13920
rect 5813 13883 5871 13889
rect 6656 13861 6684 13892
rect 6886 13892 10416 13920
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5092 13824 5641 13852
rect 5629 13821 5641 13824
rect 5675 13852 5687 13855
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 5675 13824 6101 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 6089 13821 6101 13824
rect 6135 13821 6147 13855
rect 6089 13815 6147 13821
rect 6641 13855 6699 13861
rect 6641 13821 6653 13855
rect 6687 13852 6699 13855
rect 6886 13852 6914 13892
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 10520 13929 10548 14028
rect 14384 14028 14657 14056
rect 11974 13948 11980 14000
rect 12032 13988 12038 14000
rect 13081 13991 13139 13997
rect 13081 13988 13093 13991
rect 12032 13960 13093 13988
rect 12032 13948 12038 13960
rect 13081 13957 13093 13960
rect 13127 13957 13139 13991
rect 14274 13988 14280 14000
rect 14235 13960 14280 13988
rect 13081 13951 13139 13957
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 14384 13997 14412 14028
rect 14645 14025 14657 14028
rect 14691 14056 14703 14059
rect 16850 14056 16856 14068
rect 14691 14028 16856 14056
rect 14691 14025 14703 14028
rect 14645 14019 14703 14025
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 14369 13991 14427 13997
rect 14369 13957 14381 13991
rect 14415 13957 14427 13991
rect 15194 13988 15200 14000
rect 14369 13951 14427 13957
rect 15028 13960 15200 13988
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13889 10563 13923
rect 10870 13920 10876 13932
rect 10831 13892 10876 13920
rect 10505 13883 10563 13889
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 12802 13920 12808 13932
rect 12763 13892 12808 13920
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 15028 13929 15056 13960
rect 15194 13948 15200 13960
rect 15252 13948 15258 14000
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 16209 13991 16267 13997
rect 15344 13960 15389 13988
rect 15344 13948 15350 13960
rect 16209 13957 16221 13991
rect 16255 13988 16267 13991
rect 18782 13988 18788 14000
rect 16255 13960 18788 13988
rect 16255 13957 16267 13960
rect 16209 13951 16267 13957
rect 18782 13948 18788 13960
rect 18840 13948 18846 14000
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13889 15071 13923
rect 16666 13920 16672 13932
rect 16627 13892 16672 13920
rect 15013 13883 15071 13889
rect 16666 13880 16672 13892
rect 16724 13920 16730 13932
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 16724 13892 17049 13920
rect 16724 13880 16730 13892
rect 17037 13889 17049 13892
rect 17083 13889 17095 13923
rect 17037 13883 17095 13889
rect 6687 13824 6914 13852
rect 6687 13821 6699 13824
rect 6641 13815 6699 13821
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10888 13852 10916 13880
rect 10284 13824 10916 13852
rect 11241 13855 11299 13861
rect 10284 13812 10290 13824
rect 11241 13821 11253 13855
rect 11287 13852 11299 13855
rect 12434 13852 12440 13864
rect 11287 13824 12440 13852
rect 11287 13821 11299 13824
rect 11241 13815 11299 13821
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 13722 13852 13728 13864
rect 13683 13824 13728 13852
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 15197 13855 15255 13861
rect 14792 13824 14872 13852
rect 14792 13812 14798 13824
rect 4396 13756 4752 13784
rect 4396 13744 4402 13756
rect 5718 13744 5724 13796
rect 5776 13784 5782 13796
rect 6822 13784 6828 13796
rect 5776 13756 6828 13784
rect 5776 13744 5782 13756
rect 6822 13744 6828 13756
rect 6880 13744 6886 13796
rect 14844 13793 14872 13824
rect 15197 13821 15209 13855
rect 15243 13852 15255 13855
rect 16298 13852 16304 13864
rect 15243 13824 16304 13852
rect 15243 13821 15255 13824
rect 15197 13815 15255 13821
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 18874 13852 18880 13864
rect 16868 13824 18880 13852
rect 16868 13793 16896 13824
rect 18874 13812 18880 13824
rect 18932 13812 18938 13864
rect 14829 13787 14887 13793
rect 14829 13753 14841 13787
rect 14875 13753 14887 13787
rect 14829 13747 14887 13753
rect 16853 13787 16911 13793
rect 16853 13753 16865 13787
rect 16899 13753 16911 13787
rect 16853 13747 16911 13753
rect 2774 13676 2780 13728
rect 2832 13716 2838 13728
rect 5994 13716 6000 13728
rect 2832 13688 6000 13716
rect 2832 13676 2838 13688
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 6457 13719 6515 13725
rect 6457 13685 6469 13719
rect 6503 13716 6515 13719
rect 6730 13716 6736 13728
rect 6503 13688 6736 13716
rect 6503 13685 6515 13688
rect 6457 13679 6515 13685
rect 6730 13676 6736 13688
rect 6788 13676 6794 13728
rect 1104 13626 18860 13648
rect 1104 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 3302 13626
rect 3354 13574 3366 13626
rect 3418 13574 3430 13626
rect 3482 13574 7622 13626
rect 7674 13574 7686 13626
rect 7738 13574 7750 13626
rect 7802 13574 7814 13626
rect 7866 13574 7878 13626
rect 7930 13574 12070 13626
rect 12122 13574 12134 13626
rect 12186 13574 12198 13626
rect 12250 13574 12262 13626
rect 12314 13574 12326 13626
rect 12378 13574 16518 13626
rect 16570 13574 16582 13626
rect 16634 13574 16646 13626
rect 16698 13574 16710 13626
rect 16762 13574 16774 13626
rect 16826 13574 18860 13626
rect 1104 13552 18860 13574
rect 2774 13512 2780 13524
rect 2735 13484 2780 13512
rect 2774 13472 2780 13484
rect 2832 13472 2838 13524
rect 3605 13515 3663 13521
rect 3605 13481 3617 13515
rect 3651 13512 3663 13515
rect 4614 13512 4620 13524
rect 3651 13484 4620 13512
rect 3651 13481 3663 13484
rect 3605 13475 3663 13481
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 6270 13512 6276 13524
rect 5868 13484 6276 13512
rect 5868 13472 5874 13484
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 13403 13515 13461 13521
rect 13403 13481 13415 13515
rect 13449 13512 13461 13515
rect 14274 13512 14280 13524
rect 13449 13484 14280 13512
rect 13449 13481 13461 13484
rect 13403 13475 13461 13481
rect 14274 13472 14280 13484
rect 14332 13472 14338 13524
rect 10962 13444 10968 13456
rect 6472 13416 10968 13444
rect 2961 13379 3019 13385
rect 2961 13376 2973 13379
rect 2700 13348 2973 13376
rect 2406 13200 2412 13252
rect 2464 13240 2470 13252
rect 2700 13240 2728 13348
rect 2961 13345 2973 13348
rect 3007 13345 3019 13379
rect 5166 13376 5172 13388
rect 5127 13348 5172 13376
rect 2961 13339 3019 13345
rect 5166 13336 5172 13348
rect 5224 13376 5230 13388
rect 5905 13379 5963 13385
rect 5905 13376 5917 13379
rect 5224 13348 5917 13376
rect 5224 13336 5230 13348
rect 5905 13345 5917 13348
rect 5951 13345 5963 13379
rect 6472 13376 6500 13416
rect 10962 13404 10968 13416
rect 11020 13404 11026 13456
rect 5905 13339 5963 13345
rect 6104 13348 6500 13376
rect 6549 13379 6607 13385
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 2832 13280 3249 13308
rect 2832 13268 2838 13280
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 5718 13308 5724 13320
rect 3237 13271 3295 13277
rect 4356 13280 5028 13308
rect 5679 13280 5724 13308
rect 3881 13243 3939 13249
rect 3881 13240 3893 13243
rect 2464 13212 3893 13240
rect 2464 13200 2470 13212
rect 3881 13209 3893 13212
rect 3927 13240 3939 13243
rect 4246 13240 4252 13252
rect 3927 13212 4252 13240
rect 3927 13209 3939 13212
rect 3881 13203 3939 13209
rect 4246 13200 4252 13212
rect 4304 13200 4310 13252
rect 1302 13132 1308 13184
rect 1360 13172 1366 13184
rect 3145 13175 3203 13181
rect 3145 13172 3157 13175
rect 1360 13144 3157 13172
rect 1360 13132 1366 13144
rect 3145 13141 3157 13144
rect 3191 13172 3203 13175
rect 4065 13175 4123 13181
rect 4065 13172 4077 13175
rect 3191 13144 4077 13172
rect 3191 13141 3203 13144
rect 3145 13135 3203 13141
rect 4065 13141 4077 13144
rect 4111 13172 4123 13175
rect 4356 13172 4384 13280
rect 4433 13243 4491 13249
rect 4433 13209 4445 13243
rect 4479 13240 4491 13243
rect 4893 13243 4951 13249
rect 4893 13240 4905 13243
rect 4479 13212 4905 13240
rect 4479 13209 4491 13212
rect 4433 13203 4491 13209
rect 4893 13209 4905 13212
rect 4939 13209 4951 13243
rect 5000 13240 5028 13280
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 6104 13240 6132 13348
rect 6549 13345 6561 13379
rect 6595 13376 6607 13379
rect 7466 13376 7472 13388
rect 6595 13348 7472 13376
rect 6595 13345 6607 13348
rect 6549 13339 6607 13345
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 6638 13308 6644 13320
rect 5000 13212 6132 13240
rect 6196 13280 6644 13308
rect 4893 13203 4951 13209
rect 4111 13144 4384 13172
rect 4111 13141 4123 13144
rect 4065 13135 4123 13141
rect 4522 13132 4528 13184
rect 4580 13172 4586 13184
rect 4982 13172 4988 13184
rect 4580 13144 4625 13172
rect 4943 13144 4988 13172
rect 4580 13132 4586 13144
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5074 13132 5080 13184
rect 5132 13172 5138 13184
rect 5353 13175 5411 13181
rect 5353 13172 5365 13175
rect 5132 13144 5365 13172
rect 5132 13132 5138 13144
rect 5353 13141 5365 13144
rect 5399 13141 5411 13175
rect 5353 13135 5411 13141
rect 5813 13175 5871 13181
rect 5813 13141 5825 13175
rect 5859 13172 5871 13175
rect 6196 13172 6224 13280
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 6822 13268 6828 13320
rect 6880 13308 6886 13320
rect 6880 13268 6914 13308
rect 12434 13268 12440 13320
rect 12492 13308 12498 13320
rect 13332 13311 13390 13317
rect 13332 13308 13344 13311
rect 12492 13280 13344 13308
rect 12492 13268 12498 13280
rect 13332 13277 13344 13280
rect 13378 13308 13390 13311
rect 15102 13308 15108 13320
rect 13378 13280 15108 13308
rect 13378 13277 13390 13280
rect 13332 13271 13390 13277
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 6270 13200 6276 13252
rect 6328 13240 6334 13252
rect 6733 13243 6791 13249
rect 6733 13240 6745 13243
rect 6328 13212 6745 13240
rect 6328 13200 6334 13212
rect 6733 13209 6745 13212
rect 6779 13209 6791 13243
rect 6886 13240 6914 13268
rect 13906 13240 13912 13252
rect 6886 13212 13912 13240
rect 6733 13203 6791 13209
rect 13906 13200 13912 13212
rect 13964 13200 13970 13252
rect 6638 13172 6644 13184
rect 5859 13144 6224 13172
rect 6599 13144 6644 13172
rect 5859 13141 5871 13144
rect 5813 13135 5871 13141
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 7098 13172 7104 13184
rect 7059 13144 7104 13172
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 15194 13172 15200 13184
rect 15155 13144 15200 13172
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 1104 13082 18860 13104
rect 1104 13030 5398 13082
rect 5450 13030 5462 13082
rect 5514 13030 5526 13082
rect 5578 13030 5590 13082
rect 5642 13030 5654 13082
rect 5706 13030 9846 13082
rect 9898 13030 9910 13082
rect 9962 13030 9974 13082
rect 10026 13030 10038 13082
rect 10090 13030 10102 13082
rect 10154 13030 14294 13082
rect 14346 13030 14358 13082
rect 14410 13030 14422 13082
rect 14474 13030 14486 13082
rect 14538 13030 14550 13082
rect 14602 13030 18860 13082
rect 1104 13008 18860 13030
rect 4522 12968 4528 12980
rect 4483 12940 4528 12968
rect 4522 12928 4528 12940
rect 4580 12928 4586 12980
rect 4617 12971 4675 12977
rect 4617 12937 4629 12971
rect 4663 12968 4675 12971
rect 5074 12968 5080 12980
rect 4663 12940 5080 12968
rect 4663 12937 4675 12940
rect 4617 12931 4675 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5721 12971 5779 12977
rect 5721 12937 5733 12971
rect 5767 12968 5779 12971
rect 5810 12968 5816 12980
rect 5767 12940 5816 12968
rect 5767 12937 5779 12940
rect 5721 12931 5779 12937
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 6181 12971 6239 12977
rect 6181 12937 6193 12971
rect 6227 12968 6239 12971
rect 6270 12968 6276 12980
rect 6227 12940 6276 12968
rect 6227 12937 6239 12940
rect 6181 12931 6239 12937
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 6638 12928 6644 12980
rect 6696 12968 6702 12980
rect 7009 12971 7067 12977
rect 7009 12968 7021 12971
rect 6696 12940 7021 12968
rect 6696 12928 6702 12940
rect 7009 12937 7021 12940
rect 7055 12937 7067 12971
rect 7009 12931 7067 12937
rect 7190 12928 7196 12980
rect 7248 12968 7254 12980
rect 13449 12971 13507 12977
rect 13449 12968 13461 12971
rect 7248 12940 13461 12968
rect 7248 12928 7254 12940
rect 13449 12937 13461 12940
rect 13495 12968 13507 12971
rect 14185 12971 14243 12977
rect 14185 12968 14197 12971
rect 13495 12940 14197 12968
rect 13495 12937 13507 12940
rect 13449 12931 13507 12937
rect 14185 12937 14197 12940
rect 14231 12968 14243 12971
rect 15010 12968 15016 12980
rect 14231 12940 15016 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 15010 12928 15016 12940
rect 15068 12928 15074 12980
rect 17862 12968 17868 12980
rect 16546 12940 17868 12968
rect 2130 12900 2136 12912
rect 2043 12872 2136 12900
rect 2130 12860 2136 12872
rect 2188 12900 2194 12912
rect 4890 12900 4896 12912
rect 2188 12872 4896 12900
rect 2188 12860 2194 12872
rect 4890 12860 4896 12872
rect 4948 12900 4954 12912
rect 5353 12903 5411 12909
rect 5353 12900 5365 12903
rect 4948 12872 5365 12900
rect 4948 12860 4954 12872
rect 5353 12869 5365 12872
rect 5399 12900 5411 12903
rect 6730 12900 6736 12912
rect 5399 12872 6736 12900
rect 5399 12869 5411 12872
rect 5353 12863 5411 12869
rect 6730 12860 6736 12872
rect 6788 12900 6794 12912
rect 16546 12900 16574 12940
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 6788 12872 16574 12900
rect 6788 12860 6794 12872
rect 1670 12792 1676 12844
rect 1728 12832 1734 12844
rect 4982 12832 4988 12844
rect 1728 12804 4988 12832
rect 1728 12792 1734 12804
rect 4982 12792 4988 12804
rect 5040 12832 5046 12844
rect 5169 12835 5227 12841
rect 5169 12832 5181 12835
rect 5040 12804 5181 12832
rect 5040 12792 5046 12804
rect 5169 12801 5181 12804
rect 5215 12832 5227 12835
rect 5813 12835 5871 12841
rect 5215 12804 5764 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 4706 12764 4712 12776
rect 4667 12736 4712 12764
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 5629 12767 5687 12773
rect 5629 12733 5641 12767
rect 5675 12733 5687 12767
rect 5736 12764 5764 12804
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 5859 12804 6561 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 7006 12792 7012 12844
rect 7064 12832 7070 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 7064 12804 7389 12832
rect 7064 12792 7070 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12832 7527 12835
rect 7558 12832 7564 12844
rect 7515 12804 7564 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 7558 12792 7564 12804
rect 7616 12832 7622 12844
rect 8110 12832 8116 12844
rect 7616 12804 8116 12832
rect 7616 12792 7622 12804
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 13354 12832 13360 12844
rect 13315 12804 13360 12832
rect 13354 12792 13360 12804
rect 13412 12792 13418 12844
rect 13906 12832 13912 12844
rect 13867 12804 13912 12832
rect 13906 12792 13912 12804
rect 13964 12832 13970 12844
rect 14458 12832 14464 12844
rect 13964 12804 14464 12832
rect 13964 12792 13970 12804
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 7190 12764 7196 12776
rect 5736 12736 7196 12764
rect 5629 12727 5687 12733
rect 2038 12656 2044 12708
rect 2096 12696 2102 12708
rect 2593 12699 2651 12705
rect 2593 12696 2605 12699
rect 2096 12668 2605 12696
rect 2096 12656 2102 12668
rect 2593 12665 2605 12668
rect 2639 12665 2651 12699
rect 5644 12696 5672 12727
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12764 7711 12767
rect 8202 12764 8208 12776
rect 7699 12736 8208 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 7668 12696 7696 12727
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 14826 12764 14832 12776
rect 13679 12736 14832 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 5644 12668 7696 12696
rect 2593 12659 2651 12665
rect 2501 12631 2559 12637
rect 2501 12597 2513 12631
rect 2547 12628 2559 12631
rect 2958 12628 2964 12640
rect 2547 12600 2964 12628
rect 2547 12597 2559 12600
rect 2501 12591 2559 12597
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 3510 12588 3516 12640
rect 3568 12628 3574 12640
rect 4157 12631 4215 12637
rect 4157 12628 4169 12631
rect 3568 12600 4169 12628
rect 3568 12588 3574 12600
rect 4157 12597 4169 12600
rect 4203 12597 4215 12631
rect 4157 12591 4215 12597
rect 5902 12588 5908 12640
rect 5960 12628 5966 12640
rect 6365 12631 6423 12637
rect 6365 12628 6377 12631
rect 5960 12600 6377 12628
rect 5960 12588 5966 12600
rect 6365 12597 6377 12600
rect 6411 12628 6423 12631
rect 6822 12628 6828 12640
rect 6411 12600 6828 12628
rect 6411 12597 6423 12600
rect 6365 12591 6423 12597
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 6917 12631 6975 12637
rect 6917 12597 6929 12631
rect 6963 12628 6975 12631
rect 7006 12628 7012 12640
rect 6963 12600 7012 12628
rect 6963 12597 6975 12600
rect 6917 12591 6975 12597
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 7374 12588 7380 12640
rect 7432 12628 7438 12640
rect 7929 12631 7987 12637
rect 7929 12628 7941 12631
rect 7432 12600 7941 12628
rect 7432 12588 7438 12600
rect 7929 12597 7941 12600
rect 7975 12628 7987 12631
rect 8110 12628 8116 12640
rect 7975 12600 8116 12628
rect 7975 12597 7987 12600
rect 7929 12591 7987 12597
rect 8110 12588 8116 12600
rect 8168 12588 8174 12640
rect 9677 12631 9735 12637
rect 9677 12597 9689 12631
rect 9723 12628 9735 12631
rect 10502 12628 10508 12640
rect 9723 12600 10508 12628
rect 9723 12597 9735 12600
rect 9677 12591 9735 12597
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 12986 12628 12992 12640
rect 12947 12600 12992 12628
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 1104 12538 18860 12560
rect 1104 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 3302 12538
rect 3354 12486 3366 12538
rect 3418 12486 3430 12538
rect 3482 12486 7622 12538
rect 7674 12486 7686 12538
rect 7738 12486 7750 12538
rect 7802 12486 7814 12538
rect 7866 12486 7878 12538
rect 7930 12486 12070 12538
rect 12122 12486 12134 12538
rect 12186 12486 12198 12538
rect 12250 12486 12262 12538
rect 12314 12486 12326 12538
rect 12378 12486 16518 12538
rect 16570 12486 16582 12538
rect 16634 12486 16646 12538
rect 16698 12486 16710 12538
rect 16762 12486 16774 12538
rect 16826 12486 18860 12538
rect 1104 12464 18860 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 11790 12424 11796 12436
rect 2832 12396 11796 12424
rect 2832 12384 2838 12396
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 6822 12316 6828 12368
rect 6880 12316 6886 12368
rect 6914 12316 6920 12368
rect 6972 12356 6978 12368
rect 9398 12356 9404 12368
rect 6972 12328 9404 12356
rect 6972 12316 6978 12328
rect 9398 12316 9404 12328
rect 9456 12316 9462 12368
rect 14918 12356 14924 12368
rect 9508 12328 10456 12356
rect 2225 12291 2283 12297
rect 2225 12257 2237 12291
rect 2271 12288 2283 12291
rect 2682 12288 2688 12300
rect 2271 12260 2688 12288
rect 2271 12257 2283 12260
rect 2225 12251 2283 12257
rect 2682 12248 2688 12260
rect 2740 12288 2746 12300
rect 3326 12288 3332 12300
rect 2740 12260 3332 12288
rect 2740 12248 2746 12260
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 3421 12291 3479 12297
rect 3421 12257 3433 12291
rect 3467 12288 3479 12291
rect 4433 12291 4491 12297
rect 3467 12260 3740 12288
rect 3467 12257 3479 12260
rect 3421 12251 3479 12257
rect 3712 12232 3740 12260
rect 4433 12257 4445 12291
rect 4479 12288 4491 12291
rect 4706 12288 4712 12300
rect 4479 12260 4712 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 4801 12291 4859 12297
rect 4801 12257 4813 12291
rect 4847 12288 4859 12291
rect 5997 12291 6055 12297
rect 5997 12288 6009 12291
rect 4847 12260 6009 12288
rect 4847 12257 4859 12260
rect 4801 12251 4859 12257
rect 5997 12257 6009 12260
rect 6043 12288 6055 12291
rect 6840 12288 6868 12316
rect 7009 12291 7067 12297
rect 7009 12288 7021 12291
rect 6043 12260 6776 12288
rect 6840 12260 7021 12288
rect 6043 12257 6055 12260
rect 5997 12251 6055 12257
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12220 2007 12223
rect 2130 12220 2136 12232
rect 1995 12192 2136 12220
rect 1995 12189 2007 12192
rect 1949 12183 2007 12189
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12220 3295 12223
rect 3510 12220 3516 12232
rect 3283 12192 3516 12220
rect 3283 12189 3295 12192
rect 3237 12183 3295 12189
rect 3510 12180 3516 12192
rect 3568 12180 3574 12232
rect 3694 12180 3700 12232
rect 3752 12180 3758 12232
rect 4890 12220 4896 12232
rect 4851 12192 4896 12220
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 5902 12220 5908 12232
rect 5863 12192 5908 12220
rect 5902 12180 5908 12192
rect 5960 12180 5966 12232
rect 2317 12155 2375 12161
rect 2317 12121 2329 12155
rect 2363 12152 2375 12155
rect 2590 12152 2596 12164
rect 2363 12124 2596 12152
rect 2363 12121 2375 12124
rect 2317 12115 2375 12121
rect 2590 12112 2596 12124
rect 2648 12112 2654 12164
rect 4522 12152 4528 12164
rect 2792 12124 4528 12152
rect 934 12044 940 12096
rect 992 12084 998 12096
rect 1765 12087 1823 12093
rect 1765 12084 1777 12087
rect 992 12056 1777 12084
rect 992 12044 998 12056
rect 1765 12053 1777 12056
rect 1811 12053 1823 12087
rect 1765 12047 1823 12053
rect 2409 12087 2467 12093
rect 2409 12053 2421 12087
rect 2455 12084 2467 12087
rect 2498 12084 2504 12096
rect 2455 12056 2504 12084
rect 2455 12053 2467 12056
rect 2409 12047 2467 12053
rect 2498 12044 2504 12056
rect 2556 12044 2562 12096
rect 2792 12093 2820 12124
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 4798 12112 4804 12164
rect 4856 12152 4862 12164
rect 6270 12152 6276 12164
rect 4856 12124 6276 12152
rect 4856 12112 4862 12124
rect 6270 12112 6276 12124
rect 6328 12112 6334 12164
rect 6748 12152 6776 12260
rect 7009 12257 7021 12260
rect 7055 12257 7067 12291
rect 7834 12288 7840 12300
rect 7795 12260 7840 12288
rect 7009 12251 7067 12257
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 9508 12297 9536 12328
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12257 9551 12291
rect 10226 12288 10232 12300
rect 10187 12260 10232 12288
rect 9493 12251 9551 12257
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 10428 12297 10456 12328
rect 12820 12328 14412 12356
rect 10413 12291 10471 12297
rect 10413 12257 10425 12291
rect 10459 12288 10471 12291
rect 10778 12288 10784 12300
rect 10459 12260 10784 12288
rect 10459 12257 10471 12260
rect 10413 12251 10471 12257
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 12066 12248 12072 12300
rect 12124 12288 12130 12300
rect 12529 12291 12587 12297
rect 12529 12288 12541 12291
rect 12124 12260 12541 12288
rect 12124 12248 12130 12260
rect 12529 12257 12541 12260
rect 12575 12257 12587 12291
rect 12529 12251 12587 12257
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 7098 12220 7104 12232
rect 6871 12192 7104 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 8018 12180 8024 12232
rect 8076 12220 8082 12232
rect 8202 12220 8208 12232
rect 8076 12192 8208 12220
rect 8076 12180 8082 12192
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 10244 12220 10272 12248
rect 10597 12223 10655 12229
rect 10597 12220 10609 12223
rect 10244 12192 10609 12220
rect 10597 12189 10609 12192
rect 10643 12189 10655 12223
rect 10597 12183 10655 12189
rect 11790 12180 11796 12232
rect 11848 12220 11854 12232
rect 12437 12223 12495 12229
rect 12437 12220 12449 12223
rect 11848 12192 12449 12220
rect 11848 12180 11854 12192
rect 12437 12189 12449 12192
rect 12483 12220 12495 12223
rect 12820 12220 12848 12328
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12288 12955 12291
rect 13078 12288 13084 12300
rect 12943 12260 13084 12288
rect 12943 12257 12955 12260
rect 12897 12251 12955 12257
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 13354 12248 13360 12300
rect 13412 12288 13418 12300
rect 13633 12291 13691 12297
rect 13633 12288 13645 12291
rect 13412 12260 13645 12288
rect 13412 12248 13418 12260
rect 13633 12257 13645 12260
rect 13679 12257 13691 12291
rect 13633 12251 13691 12257
rect 12483 12192 12848 12220
rect 12483 12189 12495 12192
rect 12437 12183 12495 12189
rect 12986 12180 12992 12232
rect 13044 12220 13050 12232
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 13044 12192 13185 12220
rect 13044 12180 13050 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 14384 12220 14412 12328
rect 14568 12328 14924 12356
rect 14568 12297 14596 12328
rect 14918 12316 14924 12328
rect 14976 12316 14982 12368
rect 15010 12316 15016 12368
rect 15068 12356 15074 12368
rect 18138 12356 18144 12368
rect 15068 12328 18144 12356
rect 15068 12316 15074 12328
rect 18138 12316 18144 12328
rect 18196 12316 18202 12368
rect 14553 12291 14611 12297
rect 14553 12257 14565 12291
rect 14599 12257 14611 12291
rect 14553 12251 14611 12257
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12288 14795 12291
rect 14826 12288 14832 12300
rect 14783 12260 14832 12288
rect 14783 12257 14795 12260
rect 14737 12251 14795 12257
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 17586 12248 17592 12300
rect 17644 12288 17650 12300
rect 17773 12291 17831 12297
rect 17773 12288 17785 12291
rect 17644 12260 17785 12288
rect 17644 12248 17650 12260
rect 17773 12257 17785 12260
rect 17819 12257 17831 12291
rect 17773 12251 17831 12257
rect 17494 12220 17500 12232
rect 14384 12192 17500 12220
rect 13173 12183 13231 12189
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12220 17739 12223
rect 17862 12220 17868 12232
rect 17727 12192 17868 12220
rect 17727 12189 17739 12192
rect 17681 12183 17739 12189
rect 17862 12180 17868 12192
rect 17920 12220 17926 12232
rect 18049 12223 18107 12229
rect 18049 12220 18061 12223
rect 17920 12192 18061 12220
rect 17920 12180 17926 12192
rect 18049 12189 18061 12192
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 8297 12155 8355 12161
rect 8297 12152 8309 12155
rect 6748 12124 7144 12152
rect 7116 12096 7144 12124
rect 7760 12124 8309 12152
rect 7760 12096 7788 12124
rect 8297 12121 8309 12124
rect 8343 12152 8355 12155
rect 13081 12155 13139 12161
rect 8343 12124 12388 12152
rect 8343 12121 8355 12124
rect 8297 12115 8355 12121
rect 12360 12096 12388 12124
rect 13081 12121 13093 12155
rect 13127 12152 13139 12155
rect 13127 12124 14136 12152
rect 13127 12121 13139 12124
rect 13081 12115 13139 12121
rect 2777 12087 2835 12093
rect 2777 12053 2789 12087
rect 2823 12053 2835 12087
rect 2777 12047 2835 12053
rect 2866 12044 2872 12096
rect 2924 12084 2930 12096
rect 3329 12087 3387 12093
rect 2924 12056 2969 12084
rect 2924 12044 2930 12056
rect 3329 12053 3341 12087
rect 3375 12084 3387 12087
rect 3789 12087 3847 12093
rect 3789 12084 3801 12087
rect 3375 12056 3801 12084
rect 3375 12053 3387 12056
rect 3329 12047 3387 12053
rect 3789 12053 3801 12056
rect 3835 12053 3847 12087
rect 3789 12047 3847 12053
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 4157 12087 4215 12093
rect 4157 12084 4169 12087
rect 4120 12056 4169 12084
rect 4120 12044 4126 12056
rect 4157 12053 4169 12056
rect 4203 12053 4215 12087
rect 4157 12047 4215 12053
rect 4246 12044 4252 12096
rect 4304 12084 4310 12096
rect 4304 12056 4349 12084
rect 4304 12044 4310 12056
rect 4430 12044 4436 12096
rect 4488 12084 4494 12096
rect 4982 12084 4988 12096
rect 4488 12056 4988 12084
rect 4488 12044 4494 12056
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 5258 12044 5264 12096
rect 5316 12084 5322 12096
rect 5353 12087 5411 12093
rect 5353 12084 5365 12087
rect 5316 12056 5365 12084
rect 5316 12044 5322 12056
rect 5353 12053 5365 12056
rect 5399 12053 5411 12087
rect 5353 12047 5411 12053
rect 5445 12087 5503 12093
rect 5445 12053 5457 12087
rect 5491 12084 5503 12087
rect 5718 12084 5724 12096
rect 5491 12056 5724 12084
rect 5491 12053 5503 12056
rect 5445 12047 5503 12053
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 5810 12044 5816 12096
rect 5868 12084 5874 12096
rect 6454 12084 6460 12096
rect 5868 12056 5913 12084
rect 6415 12056 6460 12084
rect 5868 12044 5874 12056
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 6972 12056 7017 12084
rect 6972 12044 6978 12056
rect 7098 12044 7104 12096
rect 7156 12044 7162 12096
rect 7282 12084 7288 12096
rect 7243 12056 7288 12084
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 7650 12084 7656 12096
rect 7611 12056 7656 12084
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 7800 12056 7845 12084
rect 7800 12044 7806 12056
rect 7926 12044 7932 12096
rect 7984 12084 7990 12096
rect 8113 12087 8171 12093
rect 8113 12084 8125 12087
rect 7984 12056 8125 12084
rect 7984 12044 7990 12056
rect 8113 12053 8125 12056
rect 8159 12053 8171 12087
rect 8938 12084 8944 12096
rect 8899 12056 8944 12084
rect 8113 12047 8171 12053
rect 8938 12044 8944 12056
rect 8996 12044 9002 12096
rect 9306 12084 9312 12096
rect 9267 12056 9312 12084
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 9490 12084 9496 12096
rect 9447 12056 9496 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 9766 12084 9772 12096
rect 9727 12056 9772 12084
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 10137 12087 10195 12093
rect 10137 12053 10149 12087
rect 10183 12084 10195 12087
rect 10502 12084 10508 12096
rect 10183 12056 10508 12084
rect 10183 12053 10195 12056
rect 10137 12047 10195 12053
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 11974 12084 11980 12096
rect 11935 12056 11980 12084
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12342 12084 12348 12096
rect 12303 12056 12348 12084
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 13538 12084 13544 12096
rect 13499 12056 13544 12084
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 14108 12093 14136 12124
rect 14093 12087 14151 12093
rect 14093 12053 14105 12087
rect 14139 12053 14151 12087
rect 14458 12084 14464 12096
rect 14371 12056 14464 12084
rect 14093 12047 14151 12053
rect 14458 12044 14464 12056
rect 14516 12084 14522 12096
rect 15010 12084 15016 12096
rect 14516 12056 15016 12084
rect 14516 12044 14522 12056
rect 15010 12044 15016 12056
rect 15068 12044 15074 12096
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17037 12087 17095 12093
rect 17037 12084 17049 12087
rect 17000 12056 17049 12084
rect 17000 12044 17006 12056
rect 17037 12053 17049 12056
rect 17083 12053 17095 12087
rect 17037 12047 17095 12053
rect 17126 12044 17132 12096
rect 17184 12084 17190 12096
rect 17221 12087 17279 12093
rect 17221 12084 17233 12087
rect 17184 12056 17233 12084
rect 17184 12044 17190 12056
rect 17221 12053 17233 12056
rect 17267 12053 17279 12087
rect 17221 12047 17279 12053
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 17589 12087 17647 12093
rect 17589 12084 17601 12087
rect 17368 12056 17601 12084
rect 17368 12044 17374 12056
rect 17589 12053 17601 12056
rect 17635 12053 17647 12087
rect 17589 12047 17647 12053
rect 17678 12044 17684 12096
rect 17736 12084 17742 12096
rect 18233 12087 18291 12093
rect 18233 12084 18245 12087
rect 17736 12056 18245 12084
rect 17736 12044 17742 12056
rect 18233 12053 18245 12056
rect 18279 12053 18291 12087
rect 18233 12047 18291 12053
rect 1104 11994 18860 12016
rect 1104 11942 5398 11994
rect 5450 11942 5462 11994
rect 5514 11942 5526 11994
rect 5578 11942 5590 11994
rect 5642 11942 5654 11994
rect 5706 11942 9846 11994
rect 9898 11942 9910 11994
rect 9962 11942 9974 11994
rect 10026 11942 10038 11994
rect 10090 11942 10102 11994
rect 10154 11942 14294 11994
rect 14346 11942 14358 11994
rect 14410 11942 14422 11994
rect 14474 11942 14486 11994
rect 14538 11942 14550 11994
rect 14602 11942 18860 11994
rect 1104 11920 18860 11942
rect 2498 11880 2504 11892
rect 2459 11852 2504 11880
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 2590 11840 2596 11892
rect 2648 11880 2654 11892
rect 2958 11880 2964 11892
rect 2648 11852 2693 11880
rect 2746 11852 2964 11880
rect 2648 11840 2654 11852
rect 1118 11772 1124 11824
rect 1176 11812 1182 11824
rect 2041 11815 2099 11821
rect 2041 11812 2053 11815
rect 1176 11784 2053 11812
rect 1176 11772 1182 11784
rect 2041 11781 2053 11784
rect 2087 11781 2099 11815
rect 2746 11812 2774 11852
rect 2958 11840 2964 11852
rect 3016 11880 3022 11892
rect 3053 11883 3111 11889
rect 3053 11880 3065 11883
rect 3016 11852 3065 11880
rect 3016 11840 3022 11852
rect 3053 11849 3065 11852
rect 3099 11849 3111 11883
rect 4062 11880 4068 11892
rect 4023 11852 4068 11880
rect 3053 11843 3111 11849
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 4522 11840 4528 11892
rect 4580 11880 4586 11892
rect 4798 11880 4804 11892
rect 4580 11852 4804 11880
rect 4580 11840 4586 11852
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 4982 11880 4988 11892
rect 4943 11852 4988 11880
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 5316 11852 5457 11880
rect 5316 11840 5322 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 5445 11843 5503 11849
rect 5537 11883 5595 11889
rect 5537 11849 5549 11883
rect 5583 11880 5595 11883
rect 5718 11880 5724 11892
rect 5583 11852 5724 11880
rect 5583 11849 5595 11852
rect 5537 11843 5595 11849
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 5810 11840 5816 11892
rect 5868 11880 5874 11892
rect 5997 11883 6055 11889
rect 5997 11880 6009 11883
rect 5868 11852 6009 11880
rect 5868 11840 5874 11852
rect 5997 11849 6009 11852
rect 6043 11849 6055 11883
rect 6914 11880 6920 11892
rect 6875 11852 6920 11880
rect 5997 11843 6055 11849
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 7285 11883 7343 11889
rect 7285 11849 7297 11883
rect 7331 11880 7343 11883
rect 7745 11883 7803 11889
rect 7745 11880 7757 11883
rect 7331 11852 7757 11880
rect 7331 11849 7343 11852
rect 7285 11843 7343 11849
rect 7745 11849 7757 11852
rect 7791 11849 7803 11883
rect 7745 11843 7803 11849
rect 8113 11883 8171 11889
rect 8113 11849 8125 11883
rect 8159 11880 8171 11883
rect 8202 11880 8208 11892
rect 8159 11852 8208 11880
rect 8159 11849 8171 11852
rect 8113 11843 8171 11849
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8938 11880 8944 11892
rect 8899 11852 8944 11880
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 9306 11840 9312 11892
rect 9364 11880 9370 11892
rect 9401 11883 9459 11889
rect 9401 11880 9413 11883
rect 9364 11852 9413 11880
rect 9364 11840 9370 11852
rect 9401 11849 9413 11852
rect 9447 11849 9459 11883
rect 9401 11843 9459 11849
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 10781 11883 10839 11889
rect 9548 11852 9904 11880
rect 9548 11840 9554 11852
rect 2041 11775 2099 11781
rect 2516 11784 2774 11812
rect 2516 11756 2544 11784
rect 3326 11772 3332 11824
rect 3384 11812 3390 11824
rect 6086 11812 6092 11824
rect 3384 11784 6092 11812
rect 3384 11772 3390 11784
rect 6086 11772 6092 11784
rect 6144 11812 6150 11824
rect 6144 11784 6316 11812
rect 6144 11772 6150 11784
rect 1670 11744 1676 11756
rect 1631 11716 1676 11744
rect 1670 11704 1676 11716
rect 1728 11704 1734 11756
rect 2130 11744 2136 11756
rect 2091 11716 2136 11744
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 2498 11704 2504 11756
rect 2556 11704 2562 11756
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11744 3019 11747
rect 3421 11747 3479 11753
rect 3421 11744 3433 11747
rect 3007 11716 3433 11744
rect 3007 11713 3019 11716
rect 2961 11707 3019 11713
rect 3421 11713 3433 11716
rect 3467 11744 3479 11747
rect 3973 11747 4031 11753
rect 3467 11716 3924 11744
rect 3467 11713 3479 11716
rect 3421 11707 3479 11713
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11645 2007 11679
rect 3237 11679 3295 11685
rect 3237 11676 3249 11679
rect 1949 11639 2007 11645
rect 2700 11648 3249 11676
rect 1964 11608 1992 11639
rect 2700 11608 2728 11648
rect 3237 11645 3249 11648
rect 3283 11676 3295 11679
rect 3510 11676 3516 11688
rect 3283 11648 3516 11676
rect 3283 11645 3295 11648
rect 3237 11639 3295 11645
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 1964 11580 2728 11608
rect 3896 11608 3924 11716
rect 3973 11713 3985 11747
rect 4019 11744 4031 11747
rect 4154 11744 4160 11756
rect 4019 11716 4160 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 4154 11704 4160 11716
rect 4212 11744 4218 11756
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 4212 11716 4445 11744
rect 4212 11704 4218 11716
rect 4433 11713 4445 11716
rect 4479 11744 4491 11747
rect 5718 11744 5724 11756
rect 4479 11716 5724 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 5718 11704 5724 11716
rect 5776 11704 5782 11756
rect 6288 11744 6316 11784
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 6457 11815 6515 11821
rect 6457 11812 6469 11815
rect 6420 11784 6469 11812
rect 6420 11772 6426 11784
rect 6457 11781 6469 11784
rect 6503 11812 6515 11815
rect 6638 11812 6644 11824
rect 6503 11784 6644 11812
rect 6503 11781 6515 11784
rect 6457 11775 6515 11781
rect 6638 11772 6644 11784
rect 6696 11772 6702 11824
rect 9033 11815 9091 11821
rect 9033 11781 9045 11815
rect 9079 11812 9091 11815
rect 9766 11812 9772 11824
rect 9079 11784 9772 11812
rect 9079 11781 9091 11784
rect 9033 11775 9091 11781
rect 9766 11772 9772 11784
rect 9824 11772 9830 11824
rect 9876 11821 9904 11852
rect 10781 11849 10793 11883
rect 10827 11880 10839 11883
rect 11974 11880 11980 11892
rect 10827 11852 11980 11880
rect 10827 11849 10839 11852
rect 10781 11843 10839 11849
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 12897 11883 12955 11889
rect 12897 11880 12909 11883
rect 12400 11852 12909 11880
rect 12400 11840 12406 11852
rect 12897 11849 12909 11852
rect 12943 11880 12955 11883
rect 15102 11880 15108 11892
rect 12943 11852 15108 11880
rect 12943 11849 12955 11852
rect 12897 11843 12955 11849
rect 15102 11840 15108 11852
rect 15160 11840 15166 11892
rect 17126 11880 17132 11892
rect 17087 11852 17132 11880
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 17681 11883 17739 11889
rect 17681 11880 17693 11883
rect 17552 11852 17693 11880
rect 17552 11840 17558 11852
rect 17681 11849 17693 11852
rect 17727 11880 17739 11883
rect 17770 11880 17776 11892
rect 17727 11852 17776 11880
rect 17727 11849 17739 11852
rect 17681 11843 17739 11849
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 17954 11880 17960 11892
rect 17915 11852 17960 11880
rect 17954 11840 17960 11852
rect 18012 11840 18018 11892
rect 9861 11815 9919 11821
rect 9861 11781 9873 11815
rect 9907 11812 9919 11815
rect 15010 11812 15016 11824
rect 9907 11784 15016 11812
rect 9907 11781 9919 11784
rect 9861 11775 9919 11781
rect 15010 11772 15016 11784
rect 15068 11772 15074 11824
rect 18049 11815 18107 11821
rect 18049 11812 18061 11815
rect 15304 11784 18061 11812
rect 6914 11744 6920 11756
rect 6288 11716 6920 11744
rect 6914 11704 6920 11716
rect 6972 11744 6978 11756
rect 7834 11744 7840 11756
rect 6972 11716 7840 11744
rect 6972 11704 6978 11716
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11744 8263 11747
rect 8938 11744 8944 11756
rect 8251 11716 8944 11744
rect 8251 11713 8263 11716
rect 8205 11707 8263 11713
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 9732 11716 10241 11744
rect 9732 11704 9738 11716
rect 10229 11713 10241 11716
rect 10275 11744 10287 11747
rect 10686 11744 10692 11756
rect 10275 11716 10692 11744
rect 10275 11713 10287 11716
rect 10229 11707 10287 11713
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11885 11747 11943 11753
rect 11885 11744 11897 11747
rect 11664 11716 11897 11744
rect 11664 11704 11670 11716
rect 11885 11713 11897 11716
rect 11931 11744 11943 11747
rect 13449 11747 13507 11753
rect 11931 11716 12480 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 4522 11676 4528 11688
rect 4483 11648 4528 11676
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11676 4767 11679
rect 4798 11676 4804 11688
rect 4755 11648 4804 11676
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 4798 11636 4804 11648
rect 4856 11676 4862 11688
rect 5166 11676 5172 11688
rect 4856 11648 5172 11676
rect 4856 11636 4862 11648
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 5353 11679 5411 11685
rect 5353 11645 5365 11679
rect 5399 11676 5411 11679
rect 6362 11676 6368 11688
rect 5399 11648 6368 11676
rect 5399 11645 5411 11648
rect 5353 11639 5411 11645
rect 6362 11636 6368 11648
rect 6420 11636 6426 11688
rect 6730 11636 6736 11688
rect 6788 11676 6794 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6788 11648 6837 11676
rect 6788 11636 6794 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 7374 11676 7380 11688
rect 7335 11648 7380 11676
rect 6825 11639 6883 11645
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 7524 11648 7569 11676
rect 7524 11636 7530 11648
rect 8110 11636 8116 11688
rect 8168 11676 8174 11688
rect 8297 11679 8355 11685
rect 8297 11676 8309 11679
rect 8168 11648 8309 11676
rect 8168 11636 8174 11648
rect 8297 11645 8309 11648
rect 8343 11645 8355 11679
rect 9122 11676 9128 11688
rect 9083 11648 9128 11676
rect 8297 11639 8355 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 10778 11636 10784 11688
rect 10836 11676 10842 11688
rect 10873 11679 10931 11685
rect 10873 11676 10885 11679
rect 10836 11648 10885 11676
rect 10836 11636 10842 11648
rect 10873 11645 10885 11648
rect 10919 11645 10931 11679
rect 10873 11639 10931 11645
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 11977 11679 12035 11685
rect 11977 11676 11989 11679
rect 11848 11648 11989 11676
rect 11848 11636 11854 11648
rect 11977 11645 11989 11648
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 12124 11648 12217 11676
rect 12124 11636 12130 11648
rect 4338 11608 4344 11620
rect 3896 11580 4344 11608
rect 4338 11568 4344 11580
rect 4396 11608 4402 11620
rect 5074 11608 5080 11620
rect 4396 11580 5080 11608
rect 4396 11568 4402 11580
rect 5074 11568 5080 11580
rect 5132 11568 5138 11620
rect 5810 11608 5816 11620
rect 5736 11580 5816 11608
rect 1486 11540 1492 11552
rect 1447 11512 1492 11540
rect 1486 11500 1492 11512
rect 1544 11500 1550 11552
rect 3694 11500 3700 11552
rect 3752 11540 3758 11552
rect 3789 11543 3847 11549
rect 3789 11540 3801 11543
rect 3752 11512 3801 11540
rect 3752 11500 3758 11512
rect 3789 11509 3801 11512
rect 3835 11540 3847 11543
rect 3878 11540 3884 11552
rect 3835 11512 3884 11540
rect 3835 11509 3847 11512
rect 3789 11503 3847 11509
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 5736 11540 5764 11580
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 9674 11608 9680 11620
rect 7984 11580 9680 11608
rect 7984 11568 7990 11580
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 11422 11568 11428 11620
rect 11480 11608 11486 11620
rect 12084 11608 12112 11636
rect 12452 11617 12480 11716
rect 13449 11713 13461 11747
rect 13495 11744 13507 11747
rect 13722 11744 13728 11756
rect 13495 11716 13728 11744
rect 13495 11713 13507 11716
rect 13449 11707 13507 11713
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 15304 11753 15332 11784
rect 18049 11781 18061 11784
rect 18095 11812 18107 11815
rect 18230 11812 18236 11824
rect 18095 11784 18236 11812
rect 18095 11781 18107 11784
rect 18049 11775 18107 11781
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 15289 11747 15347 11753
rect 15289 11744 15301 11747
rect 14792 11716 15301 11744
rect 14792 11704 14798 11716
rect 15289 11713 15301 11716
rect 15335 11713 15347 11747
rect 17034 11744 17040 11756
rect 16995 11716 17040 11744
rect 15289 11707 15347 11713
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 13541 11679 13599 11685
rect 13541 11676 13553 11679
rect 13320 11648 13553 11676
rect 13320 11636 13326 11648
rect 13541 11645 13553 11648
rect 13587 11645 13599 11679
rect 13541 11639 13599 11645
rect 13630 11636 13636 11688
rect 13688 11676 13694 11688
rect 15102 11685 15108 11688
rect 15059 11679 15108 11685
rect 13688 11648 13733 11676
rect 13688 11636 13694 11648
rect 15059 11645 15071 11679
rect 15105 11645 15108 11679
rect 15059 11639 15108 11645
rect 15102 11636 15108 11639
rect 15160 11636 15166 11688
rect 15197 11679 15255 11685
rect 15197 11645 15209 11679
rect 15243 11645 15255 11679
rect 15197 11639 15255 11645
rect 11480 11580 12112 11608
rect 12437 11611 12495 11617
rect 11480 11568 11486 11580
rect 12437 11577 12449 11611
rect 12483 11608 12495 11611
rect 15212 11608 15240 11639
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 17221 11679 17279 11685
rect 15712 11648 16712 11676
rect 15712 11636 15718 11648
rect 15841 11611 15899 11617
rect 15841 11608 15853 11611
rect 12483 11580 15853 11608
rect 12483 11577 12495 11580
rect 12437 11571 12495 11577
rect 15841 11577 15853 11580
rect 15887 11608 15899 11611
rect 16390 11608 16396 11620
rect 15887 11580 16396 11608
rect 15887 11577 15899 11580
rect 15841 11571 15899 11577
rect 16390 11568 16396 11580
rect 16448 11568 16454 11620
rect 16684 11617 16712 11648
rect 17221 11645 17233 11679
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 16669 11611 16727 11617
rect 16669 11577 16681 11611
rect 16715 11577 16727 11611
rect 16669 11571 16727 11577
rect 5902 11540 5908 11552
rect 4028 11512 5764 11540
rect 5863 11512 5908 11540
rect 4028 11500 4034 11512
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 8352 11512 8585 11540
rect 8352 11500 8358 11512
rect 8573 11509 8585 11512
rect 8619 11509 8631 11543
rect 10318 11540 10324 11552
rect 10279 11512 10324 11540
rect 8573 11503 8631 11509
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 11146 11540 11152 11552
rect 10468 11512 11152 11540
rect 10468 11500 10474 11512
rect 11146 11500 11152 11512
rect 11204 11540 11210 11552
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 11204 11512 11253 11540
rect 11204 11500 11210 11512
rect 11241 11509 11253 11512
rect 11287 11509 11299 11543
rect 11241 11503 11299 11509
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 11517 11543 11575 11549
rect 11517 11540 11529 11543
rect 11388 11512 11529 11540
rect 11388 11500 11394 11512
rect 11517 11509 11529 11512
rect 11563 11509 11575 11543
rect 13078 11540 13084 11552
rect 13039 11512 13084 11540
rect 11517 11503 11575 11509
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 13446 11540 13452 11552
rect 13320 11512 13452 11540
rect 13320 11500 13326 11512
rect 13446 11500 13452 11512
rect 13504 11540 13510 11552
rect 13909 11543 13967 11549
rect 13909 11540 13921 11543
rect 13504 11512 13921 11540
rect 13504 11500 13510 11512
rect 13909 11509 13921 11512
rect 13955 11509 13967 11543
rect 14734 11540 14740 11552
rect 14695 11512 14740 11540
rect 13909 11503 13967 11509
rect 14734 11500 14740 11512
rect 14792 11500 14798 11552
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 15657 11543 15715 11549
rect 15657 11540 15669 11543
rect 15528 11512 15669 11540
rect 15528 11500 15534 11512
rect 15657 11509 15669 11512
rect 15703 11509 15715 11543
rect 15657 11503 15715 11509
rect 15930 11500 15936 11552
rect 15988 11540 15994 11552
rect 17236 11540 17264 11639
rect 15988 11512 17264 11540
rect 15988 11500 15994 11512
rect 17862 11500 17868 11552
rect 17920 11540 17926 11552
rect 18325 11543 18383 11549
rect 18325 11540 18337 11543
rect 17920 11512 18337 11540
rect 17920 11500 17926 11512
rect 18325 11509 18337 11512
rect 18371 11509 18383 11543
rect 18325 11503 18383 11509
rect 1104 11450 18860 11472
rect 1104 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 3302 11450
rect 3354 11398 3366 11450
rect 3418 11398 3430 11450
rect 3482 11398 7622 11450
rect 7674 11398 7686 11450
rect 7738 11398 7750 11450
rect 7802 11398 7814 11450
rect 7866 11398 7878 11450
rect 7930 11398 12070 11450
rect 12122 11398 12134 11450
rect 12186 11398 12198 11450
rect 12250 11398 12262 11450
rect 12314 11398 12326 11450
rect 12378 11398 16518 11450
rect 16570 11398 16582 11450
rect 16634 11398 16646 11450
rect 16698 11398 16710 11450
rect 16762 11398 16774 11450
rect 16826 11398 18860 11450
rect 1104 11376 18860 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2593 11339 2651 11345
rect 2593 11305 2605 11339
rect 2639 11336 2651 11339
rect 2774 11336 2780 11348
rect 2639 11308 2780 11336
rect 2639 11305 2651 11308
rect 2593 11299 2651 11305
rect 2774 11296 2780 11308
rect 2832 11336 2838 11348
rect 2832 11308 3096 11336
rect 2832 11296 2838 11308
rect 1394 11228 1400 11280
rect 1452 11268 1458 11280
rect 2133 11271 2191 11277
rect 2133 11268 2145 11271
rect 1452 11240 2145 11268
rect 1452 11228 1458 11240
rect 2133 11237 2145 11240
rect 2179 11237 2191 11271
rect 2133 11231 2191 11237
rect 2682 11160 2688 11212
rect 2740 11200 2746 11212
rect 2777 11203 2835 11209
rect 2777 11200 2789 11203
rect 2740 11172 2789 11200
rect 2740 11160 2746 11172
rect 2777 11169 2789 11172
rect 2823 11169 2835 11203
rect 2777 11163 2835 11169
rect 1949 11135 2007 11141
rect 1949 11101 1961 11135
rect 1995 11132 2007 11135
rect 2314 11132 2320 11144
rect 1995 11104 2320 11132
rect 1995 11101 2007 11104
rect 1949 11095 2007 11101
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 3068 11141 3096 11308
rect 4246 11296 4252 11348
rect 4304 11336 4310 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4304 11308 4537 11336
rect 4304 11296 4310 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 6178 11336 6184 11348
rect 4525 11299 4583 11305
rect 4724 11308 6184 11336
rect 3421 11271 3479 11277
rect 3421 11237 3433 11271
rect 3467 11268 3479 11271
rect 3467 11240 4292 11268
rect 3467 11237 3479 11240
rect 3421 11231 3479 11237
rect 3973 11203 4031 11209
rect 3973 11169 3985 11203
rect 4019 11169 4031 11203
rect 3973 11163 4031 11169
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 2682 11024 2688 11076
rect 2740 11064 2746 11076
rect 2961 11067 3019 11073
rect 2961 11064 2973 11067
rect 2740 11036 2973 11064
rect 2740 11024 2746 11036
rect 2961 11033 2973 11036
rect 3007 11033 3019 11067
rect 3988 11064 4016 11163
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11132 4123 11135
rect 4154 11132 4160 11144
rect 4111 11104 4160 11132
rect 4111 11101 4123 11104
rect 4065 11095 4123 11101
rect 4154 11092 4160 11104
rect 4212 11092 4218 11144
rect 4264 11132 4292 11240
rect 4724 11209 4752 11308
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7834 11336 7840 11348
rect 7248 11308 7840 11336
rect 7248 11296 7254 11308
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 8478 11336 8484 11348
rect 7944 11308 8484 11336
rect 5166 11228 5172 11280
rect 5224 11268 5230 11280
rect 5537 11271 5595 11277
rect 5537 11268 5549 11271
rect 5224 11240 5549 11268
rect 5224 11228 5230 11240
rect 5537 11237 5549 11240
rect 5583 11237 5595 11271
rect 6365 11271 6423 11277
rect 6365 11268 6377 11271
rect 5537 11231 5595 11237
rect 5920 11240 6377 11268
rect 4709 11203 4767 11209
rect 4709 11169 4721 11203
rect 4755 11169 4767 11203
rect 4890 11200 4896 11212
rect 4851 11172 4896 11200
rect 4709 11163 4767 11169
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 5920 11141 5948 11240
rect 6365 11237 6377 11240
rect 6411 11237 6423 11271
rect 6365 11231 6423 11237
rect 6546 11228 6552 11280
rect 6604 11268 6610 11280
rect 7944 11268 7972 11308
rect 8478 11296 8484 11308
rect 8536 11336 8542 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8536 11308 8953 11336
rect 8536 11296 8542 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 14734 11336 14740 11348
rect 9180 11308 10272 11336
rect 9180 11296 9186 11308
rect 6604 11240 7972 11268
rect 8021 11271 8079 11277
rect 6604 11228 6610 11240
rect 8021 11237 8033 11271
rect 8067 11237 8079 11271
rect 9309 11271 9367 11277
rect 9309 11268 9321 11271
rect 8021 11231 8079 11237
rect 8496 11240 9321 11268
rect 6178 11200 6184 11212
rect 6139 11172 6184 11200
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6638 11160 6644 11212
rect 6696 11200 6702 11212
rect 6825 11203 6883 11209
rect 6825 11200 6837 11203
rect 6696 11172 6837 11200
rect 6696 11160 6702 11172
rect 6825 11169 6837 11172
rect 6871 11169 6883 11203
rect 6825 11163 6883 11169
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 6972 11172 7017 11200
rect 6972 11160 6978 11172
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 7742 11200 7748 11212
rect 7156 11172 7748 11200
rect 7156 11160 7162 11172
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 8036 11144 8064 11231
rect 8496 11209 8524 11240
rect 9309 11237 9321 11240
rect 9355 11237 9367 11271
rect 10137 11271 10195 11277
rect 10137 11268 10149 11271
rect 9309 11231 9367 11237
rect 9784 11240 10149 11268
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11169 8539 11203
rect 8481 11163 8539 11169
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 9784 11209 9812 11240
rect 10137 11237 10149 11240
rect 10183 11237 10195 11271
rect 10137 11231 10195 11237
rect 9769 11203 9827 11209
rect 8628 11172 8673 11200
rect 8628 11160 8634 11172
rect 9769 11169 9781 11203
rect 9815 11169 9827 11203
rect 9769 11163 9827 11169
rect 9953 11203 10011 11209
rect 9953 11169 9965 11203
rect 9999 11200 10011 11203
rect 10244 11200 10272 11308
rect 9999 11172 10272 11200
rect 10428 11308 14740 11336
rect 9999 11169 10011 11172
rect 9953 11163 10011 11169
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4264 11104 4997 11132
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11101 5963 11135
rect 6730 11132 6736 11144
rect 6691 11104 6736 11132
rect 5905 11095 5963 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 8018 11092 8024 11144
rect 8076 11092 8082 11144
rect 9677 11135 9735 11141
rect 8588 11104 9536 11132
rect 4798 11064 4804 11076
rect 3988 11036 4804 11064
rect 2961 11027 3019 11033
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 5997 11067 6055 11073
rect 5997 11033 6009 11067
rect 6043 11064 6055 11067
rect 7282 11064 7288 11076
rect 6043 11036 7288 11064
rect 6043 11033 6055 11036
rect 5997 11027 6055 11033
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 7650 11064 7656 11076
rect 7611 11036 7656 11064
rect 7650 11024 7656 11036
rect 7708 11064 7714 11076
rect 7926 11064 7932 11076
rect 7708 11036 7932 11064
rect 7708 11024 7714 11036
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 8588 11064 8616 11104
rect 8036 11036 8616 11064
rect 1118 10956 1124 11008
rect 1176 10996 1182 11008
rect 1489 10999 1547 11005
rect 1489 10996 1501 10999
rect 1176 10968 1501 10996
rect 1176 10956 1182 10968
rect 1489 10965 1501 10968
rect 1535 10965 1547 10999
rect 1489 10959 1547 10965
rect 2590 10956 2596 11008
rect 2648 10996 2654 11008
rect 2866 10996 2872 11008
rect 2648 10968 2872 10996
rect 2648 10956 2654 10968
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 4157 10999 4215 11005
rect 4157 10965 4169 10999
rect 4203 10996 4215 10999
rect 4246 10996 4252 11008
rect 4203 10968 4252 10996
rect 4203 10965 4215 10968
rect 4157 10959 4215 10965
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 4430 10956 4436 11008
rect 4488 10996 4494 11008
rect 4982 10996 4988 11008
rect 4488 10968 4988 10996
rect 4488 10956 4494 10968
rect 4982 10956 4988 10968
rect 5040 10956 5046 11008
rect 5258 10956 5264 11008
rect 5316 10996 5322 11008
rect 5353 10999 5411 11005
rect 5353 10996 5365 10999
rect 5316 10968 5365 10996
rect 5316 10956 5322 10968
rect 5353 10965 5365 10968
rect 5399 10965 5411 10999
rect 5353 10959 5411 10965
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 7193 10999 7251 11005
rect 7193 10996 7205 10999
rect 6512 10968 7205 10996
rect 6512 10956 6518 10968
rect 7193 10965 7205 10968
rect 7239 10965 7251 10999
rect 7558 10996 7564 11008
rect 7519 10968 7564 10996
rect 7193 10959 7251 10965
rect 7558 10956 7564 10968
rect 7616 10996 7622 11008
rect 8036 10996 8064 11036
rect 8662 11024 8668 11076
rect 8720 11064 8726 11076
rect 9125 11067 9183 11073
rect 9125 11064 9137 11067
rect 8720 11036 9137 11064
rect 8720 11024 8726 11036
rect 9125 11033 9137 11036
rect 9171 11064 9183 11067
rect 9398 11064 9404 11076
rect 9171 11036 9404 11064
rect 9171 11033 9183 11036
rect 9125 11027 9183 11033
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 9508 11064 9536 11104
rect 9677 11101 9689 11135
rect 9723 11132 9735 11135
rect 10318 11132 10324 11144
rect 9723 11104 10324 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 10428 11064 10456 11308
rect 14734 11296 14740 11308
rect 14792 11296 14798 11348
rect 14826 11296 14832 11348
rect 14884 11336 14890 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 14884 11308 14933 11336
rect 14884 11296 14890 11308
rect 14921 11305 14933 11308
rect 14967 11336 14979 11339
rect 15010 11336 15016 11348
rect 14967 11308 15016 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 15102 11296 15108 11348
rect 15160 11336 15166 11348
rect 17034 11336 17040 11348
rect 15160 11308 16896 11336
rect 16995 11308 17040 11336
rect 15160 11296 15166 11308
rect 10965 11271 11023 11277
rect 10965 11268 10977 11271
rect 10612 11240 10977 11268
rect 10612 11209 10640 11240
rect 10965 11237 10977 11240
rect 11011 11237 11023 11271
rect 14093 11271 14151 11277
rect 14093 11268 14105 11271
rect 10965 11231 11023 11237
rect 13004 11240 14105 11268
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11169 10655 11203
rect 10778 11200 10784 11212
rect 10739 11172 10784 11200
rect 10597 11163 10655 11169
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 11422 11160 11428 11212
rect 11480 11200 11486 11212
rect 13004 11209 13032 11240
rect 14093 11237 14105 11240
rect 14139 11237 14151 11271
rect 14093 11231 14151 11237
rect 14182 11228 14188 11280
rect 14240 11268 14246 11280
rect 16485 11271 16543 11277
rect 16485 11268 16497 11271
rect 14240 11240 16497 11268
rect 14240 11228 14246 11240
rect 16485 11237 16497 11240
rect 16531 11268 16543 11271
rect 16758 11268 16764 11280
rect 16531 11240 16764 11268
rect 16531 11237 16543 11240
rect 16485 11231 16543 11237
rect 16758 11228 16764 11240
rect 16816 11228 16822 11280
rect 16868 11268 16896 11308
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 18049 11339 18107 11345
rect 18049 11305 18061 11339
rect 18095 11336 18107 11339
rect 18874 11336 18880 11348
rect 18095 11308 18880 11336
rect 18095 11305 18107 11308
rect 18049 11299 18107 11305
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 17954 11268 17960 11280
rect 16868 11240 17960 11268
rect 11517 11203 11575 11209
rect 11517 11200 11529 11203
rect 11480 11172 11529 11200
rect 11480 11160 11486 11172
rect 11517 11169 11529 11172
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 12897 11203 12955 11209
rect 12897 11169 12909 11203
rect 12943 11169 12955 11203
rect 12897 11163 12955 11169
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11169 13047 11203
rect 12989 11163 13047 11169
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11132 10563 11135
rect 11330 11132 11336 11144
rect 10551 11104 11336 11132
rect 10551 11101 10563 11104
rect 10505 11095 10563 11101
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 9508 11036 10456 11064
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 11425 11067 11483 11073
rect 11425 11064 11437 11067
rect 11112 11036 11437 11064
rect 11112 11024 11118 11036
rect 11425 11033 11437 11036
rect 11471 11064 11483 11067
rect 11974 11064 11980 11076
rect 11471 11036 11980 11064
rect 11471 11033 11483 11036
rect 11425 11027 11483 11033
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 12710 11064 12716 11076
rect 12084 11036 12716 11064
rect 7616 10968 8064 10996
rect 7616 10956 7622 10968
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 8389 10999 8447 11005
rect 8389 10996 8401 10999
rect 8352 10968 8401 10996
rect 8352 10956 8358 10968
rect 8389 10965 8401 10968
rect 8435 10965 8447 10999
rect 8389 10959 8447 10965
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 11333 10999 11391 11005
rect 11333 10996 11345 10999
rect 8536 10968 11345 10996
rect 8536 10956 8542 10968
rect 11333 10965 11345 10968
rect 11379 10996 11391 10999
rect 11793 10999 11851 11005
rect 11793 10996 11805 10999
rect 11379 10968 11805 10996
rect 11379 10965 11391 10968
rect 11333 10959 11391 10965
rect 11793 10965 11805 10968
rect 11839 10996 11851 10999
rect 12084 10996 12112 11036
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 12912 11064 12940 11163
rect 13630 11160 13636 11212
rect 13688 11200 13694 11212
rect 14645 11203 14703 11209
rect 14645 11200 14657 11203
rect 13688 11172 14657 11200
rect 13688 11160 13694 11172
rect 14645 11169 14657 11172
rect 14691 11200 14703 11203
rect 15562 11200 15568 11212
rect 14691 11172 15568 11200
rect 14691 11169 14703 11172
rect 14645 11163 14703 11169
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11200 15807 11203
rect 15838 11200 15844 11212
rect 15795 11172 15844 11200
rect 15795 11169 15807 11172
rect 15749 11163 15807 11169
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 17512 11209 17540 11240
rect 17954 11228 17960 11240
rect 18012 11228 18018 11280
rect 18417 11271 18475 11277
rect 18417 11237 18429 11271
rect 18463 11268 18475 11271
rect 18690 11268 18696 11280
rect 18463 11240 18696 11268
rect 18463 11237 18475 11240
rect 18417 11231 18475 11237
rect 18690 11228 18696 11240
rect 18748 11228 18754 11280
rect 17497 11203 17555 11209
rect 17497 11169 17509 11203
rect 17543 11169 17555 11203
rect 17497 11163 17555 11169
rect 17586 11160 17592 11212
rect 17644 11200 17650 11212
rect 17644 11172 17689 11200
rect 17644 11160 17650 11172
rect 13078 11132 13084 11144
rect 13039 11104 13084 11132
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 13228 11104 13768 11132
rect 13228 11092 13234 11104
rect 13630 11064 13636 11076
rect 12912 11036 13636 11064
rect 13630 11024 13636 11036
rect 13688 11024 13694 11076
rect 13740 11064 13768 11104
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 13909 11135 13967 11141
rect 13909 11132 13921 11135
rect 13872 11104 13921 11132
rect 13872 11092 13878 11104
rect 13909 11101 13921 11104
rect 13955 11132 13967 11135
rect 14458 11132 14464 11144
rect 13955 11104 14464 11132
rect 13955 11101 13967 11104
rect 13909 11095 13967 11101
rect 14458 11092 14464 11104
rect 14516 11092 14522 11144
rect 16022 11132 16028 11144
rect 15488 11104 16028 11132
rect 14553 11067 14611 11073
rect 13740 11036 13952 11064
rect 13924 11008 13952 11036
rect 14553 11033 14565 11067
rect 14599 11064 14611 11067
rect 15488 11064 15516 11104
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 16114 11092 16120 11144
rect 16172 11132 16178 11144
rect 16669 11135 16727 11141
rect 16669 11132 16681 11135
rect 16172 11104 16681 11132
rect 16172 11092 16178 11104
rect 16669 11101 16681 11104
rect 16715 11132 16727 11135
rect 16850 11132 16856 11144
rect 16715 11104 16856 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 16850 11092 16856 11104
rect 16908 11092 16914 11144
rect 17770 11092 17776 11144
rect 17828 11132 17834 11144
rect 17865 11135 17923 11141
rect 17865 11132 17877 11135
rect 17828 11104 17877 11132
rect 17828 11092 17834 11104
rect 17865 11101 17877 11104
rect 17911 11101 17923 11135
rect 18230 11132 18236 11144
rect 18191 11104 18236 11132
rect 17865 11095 17923 11101
rect 18230 11092 18236 11104
rect 18288 11092 18294 11144
rect 14599 11036 15516 11064
rect 15565 11067 15623 11073
rect 14599 11033 14611 11036
rect 14553 11027 14611 11033
rect 15565 11033 15577 11067
rect 15611 11064 15623 11067
rect 16574 11064 16580 11076
rect 15611 11036 16580 11064
rect 15611 11033 15623 11036
rect 15565 11027 15623 11033
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 13446 10996 13452 11008
rect 11839 10968 12112 10996
rect 13407 10968 13452 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 13446 10956 13452 10968
rect 13504 10956 13510 11008
rect 13906 10956 13912 11008
rect 13964 10956 13970 11008
rect 15102 10996 15108 11008
rect 15063 10968 15108 10996
rect 15102 10956 15108 10968
rect 15160 10956 15166 11008
rect 15470 10996 15476 11008
rect 15431 10968 15476 10996
rect 15470 10956 15476 10968
rect 15528 10956 15534 11008
rect 16206 10996 16212 11008
rect 16167 10968 16212 10996
rect 16206 10956 16212 10968
rect 16264 10956 16270 11008
rect 16850 10956 16856 11008
rect 16908 10996 16914 11008
rect 17126 10996 17132 11008
rect 16908 10968 17132 10996
rect 16908 10956 16914 10968
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 17402 10996 17408 11008
rect 17363 10968 17408 10996
rect 17402 10956 17408 10968
rect 17460 10956 17466 11008
rect 1104 10906 18860 10928
rect 1104 10854 5398 10906
rect 5450 10854 5462 10906
rect 5514 10854 5526 10906
rect 5578 10854 5590 10906
rect 5642 10854 5654 10906
rect 5706 10854 9846 10906
rect 9898 10854 9910 10906
rect 9962 10854 9974 10906
rect 10026 10854 10038 10906
rect 10090 10854 10102 10906
rect 10154 10854 14294 10906
rect 14346 10854 14358 10906
rect 14410 10854 14422 10906
rect 14474 10854 14486 10906
rect 14538 10854 14550 10906
rect 14602 10854 18860 10906
rect 1104 10832 18860 10854
rect 2406 10752 2412 10804
rect 2464 10792 2470 10804
rect 2501 10795 2559 10801
rect 2501 10792 2513 10795
rect 2464 10764 2513 10792
rect 2464 10752 2470 10764
rect 2501 10761 2513 10764
rect 2547 10761 2559 10795
rect 2682 10792 2688 10804
rect 2643 10764 2688 10792
rect 2501 10755 2559 10761
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 3050 10752 3056 10804
rect 3108 10752 3114 10804
rect 3145 10795 3203 10801
rect 3145 10761 3157 10795
rect 3191 10792 3203 10795
rect 3418 10792 3424 10804
rect 3191 10764 3424 10792
rect 3191 10761 3203 10764
rect 3145 10755 3203 10761
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 4249 10795 4307 10801
rect 4249 10761 4261 10795
rect 4295 10792 4307 10795
rect 4522 10792 4528 10804
rect 4295 10764 4528 10792
rect 4295 10761 4307 10764
rect 4249 10755 4307 10761
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 4890 10792 4896 10804
rect 4764 10764 4896 10792
rect 4764 10752 4770 10764
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5074 10752 5080 10804
rect 5132 10792 5138 10804
rect 5261 10795 5319 10801
rect 5261 10792 5273 10795
rect 5132 10764 5273 10792
rect 5132 10752 5138 10764
rect 5261 10761 5273 10764
rect 5307 10792 5319 10795
rect 5626 10792 5632 10804
rect 5307 10764 5632 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 6089 10795 6147 10801
rect 6089 10792 6101 10795
rect 5776 10764 6101 10792
rect 5776 10752 5782 10764
rect 6089 10761 6101 10764
rect 6135 10792 6147 10795
rect 7558 10792 7564 10804
rect 6135 10764 7564 10792
rect 6135 10761 6147 10764
rect 6089 10755 6147 10761
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 7650 10752 7656 10804
rect 7708 10752 7714 10804
rect 7745 10795 7803 10801
rect 7745 10761 7757 10795
rect 7791 10792 7803 10795
rect 8113 10795 8171 10801
rect 8113 10792 8125 10795
rect 7791 10764 8125 10792
rect 7791 10761 7803 10764
rect 7745 10755 7803 10761
rect 8113 10761 8125 10764
rect 8159 10761 8171 10795
rect 8478 10792 8484 10804
rect 8439 10764 8484 10792
rect 8113 10755 8171 10761
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 8938 10792 8944 10804
rect 8899 10764 8944 10792
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9398 10792 9404 10804
rect 9359 10764 9404 10792
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 10229 10795 10287 10801
rect 10229 10761 10241 10795
rect 10275 10792 10287 10795
rect 10594 10792 10600 10804
rect 10275 10764 10600 10792
rect 10275 10761 10287 10764
rect 10229 10755 10287 10761
rect 10594 10752 10600 10764
rect 10652 10752 10658 10804
rect 10873 10795 10931 10801
rect 10873 10761 10885 10795
rect 10919 10792 10931 10795
rect 11054 10792 11060 10804
rect 10919 10764 11060 10792
rect 10919 10761 10931 10764
rect 10873 10755 10931 10761
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11238 10792 11244 10804
rect 11199 10764 11244 10792
rect 11238 10752 11244 10764
rect 11296 10792 11302 10804
rect 11885 10795 11943 10801
rect 11885 10792 11897 10795
rect 11296 10764 11897 10792
rect 11296 10752 11302 10764
rect 11885 10761 11897 10764
rect 11931 10792 11943 10795
rect 11931 10764 12756 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 1581 10727 1639 10733
rect 1581 10693 1593 10727
rect 1627 10724 1639 10727
rect 2041 10727 2099 10733
rect 2041 10724 2053 10727
rect 1627 10696 2053 10724
rect 1627 10693 1639 10696
rect 1581 10687 1639 10693
rect 2041 10693 2053 10696
rect 2087 10724 2099 10727
rect 3068 10724 3096 10752
rect 3605 10727 3663 10733
rect 3605 10724 3617 10727
rect 2087 10696 3096 10724
rect 3160 10696 3617 10724
rect 2087 10693 2099 10696
rect 2041 10687 2099 10693
rect 2406 10656 2412 10668
rect 1780 10628 2412 10656
rect 1780 10597 1808 10628
rect 2406 10616 2412 10628
rect 2464 10656 2470 10668
rect 2682 10656 2688 10668
rect 2464 10628 2688 10656
rect 2464 10616 2470 10628
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3160 10656 3188 10696
rect 3605 10693 3617 10696
rect 3651 10724 3663 10727
rect 4062 10724 4068 10736
rect 3651 10696 4068 10724
rect 3651 10693 3663 10696
rect 3605 10687 3663 10693
rect 4062 10684 4068 10696
rect 4120 10724 4126 10736
rect 4617 10727 4675 10733
rect 4617 10724 4629 10727
rect 4120 10696 4629 10724
rect 4120 10684 4126 10696
rect 4617 10693 4629 10696
rect 4663 10724 4675 10727
rect 5644 10724 5672 10752
rect 6546 10724 6552 10736
rect 4663 10696 5212 10724
rect 5644 10696 6552 10724
rect 4663 10693 4675 10696
rect 4617 10687 4675 10693
rect 3099 10628 3188 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3418 10616 3424 10668
rect 3476 10656 3482 10668
rect 4706 10656 4712 10668
rect 3476 10628 4712 10656
rect 3476 10616 3482 10628
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10557 1823 10591
rect 1946 10588 1952 10600
rect 1907 10560 1952 10588
rect 1765 10551 1823 10557
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 3510 10588 3516 10600
rect 3375 10560 3516 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 3510 10548 3516 10560
rect 3568 10548 3574 10600
rect 4172 10597 4200 10628
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 4157 10591 4215 10597
rect 4157 10557 4169 10591
rect 4203 10557 4215 10591
rect 4157 10551 4215 10557
rect 4430 10548 4436 10600
rect 4488 10588 4494 10600
rect 5184 10597 5212 10696
rect 6546 10684 6552 10696
rect 6604 10684 6610 10736
rect 7282 10684 7288 10736
rect 7340 10724 7346 10736
rect 7668 10724 7696 10752
rect 7340 10696 7696 10724
rect 7340 10684 7346 10696
rect 8202 10684 8208 10736
rect 8260 10724 8266 10736
rect 12618 10724 12624 10736
rect 8260 10696 12624 10724
rect 8260 10684 8266 10696
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 12728 10724 12756 10764
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12860 10764 12909 10792
rect 12860 10752 12866 10764
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 12897 10755 12955 10761
rect 13265 10795 13323 10801
rect 13265 10761 13277 10795
rect 13311 10792 13323 10795
rect 13446 10792 13452 10804
rect 13311 10764 13452 10792
rect 13311 10761 13323 10764
rect 13265 10755 13323 10761
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 13722 10792 13728 10804
rect 13683 10764 13728 10792
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 14461 10795 14519 10801
rect 14461 10761 14473 10795
rect 14507 10792 14519 10795
rect 15102 10792 15108 10804
rect 14507 10764 15108 10792
rect 14507 10761 14519 10764
rect 14461 10755 14519 10761
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 15289 10795 15347 10801
rect 15289 10761 15301 10795
rect 15335 10792 15347 10795
rect 15749 10795 15807 10801
rect 15749 10792 15761 10795
rect 15335 10764 15761 10792
rect 15335 10761 15347 10764
rect 15289 10755 15347 10761
rect 15749 10761 15761 10764
rect 15795 10761 15807 10795
rect 15749 10755 15807 10761
rect 16574 10752 16580 10804
rect 16632 10792 16638 10804
rect 16669 10795 16727 10801
rect 16669 10792 16681 10795
rect 16632 10764 16681 10792
rect 16632 10752 16638 10764
rect 16669 10761 16681 10764
rect 16715 10761 16727 10795
rect 16669 10755 16727 10761
rect 16758 10752 16764 10804
rect 16816 10792 16822 10804
rect 17037 10795 17095 10801
rect 17037 10792 17049 10795
rect 16816 10764 17049 10792
rect 16816 10752 16822 10764
rect 17037 10761 17049 10764
rect 17083 10761 17095 10795
rect 17037 10755 17095 10761
rect 17402 10752 17408 10804
rect 17460 10792 17466 10804
rect 17497 10795 17555 10801
rect 17497 10792 17509 10795
rect 17460 10764 17509 10792
rect 17460 10752 17466 10764
rect 17497 10761 17509 10764
rect 17543 10761 17555 10795
rect 17497 10755 17555 10761
rect 13814 10724 13820 10736
rect 12728 10696 13820 10724
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 14369 10727 14427 10733
rect 14369 10693 14381 10727
rect 14415 10724 14427 10727
rect 14415 10696 14964 10724
rect 14415 10693 14427 10696
rect 14369 10687 14427 10693
rect 5994 10656 6000 10668
rect 5907 10628 6000 10656
rect 5994 10616 6000 10628
rect 6052 10656 6058 10668
rect 6730 10656 6736 10668
rect 6052 10628 6736 10656
rect 6052 10616 6058 10628
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 7558 10656 7564 10668
rect 6840 10628 7564 10656
rect 4801 10591 4859 10597
rect 4801 10588 4813 10591
rect 4488 10560 4813 10588
rect 4488 10548 4494 10560
rect 4801 10557 4813 10560
rect 4847 10557 4859 10591
rect 4801 10551 4859 10557
rect 5169 10591 5227 10597
rect 5169 10557 5181 10591
rect 5215 10588 5227 10591
rect 5350 10588 5356 10600
rect 5215 10560 5356 10588
rect 5215 10557 5227 10560
rect 5169 10551 5227 10557
rect 5350 10548 5356 10560
rect 5408 10548 5414 10600
rect 6840 10597 6868 10628
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 7653 10659 7711 10665
rect 7653 10625 7665 10659
rect 7699 10656 7711 10659
rect 8294 10656 8300 10668
rect 7699 10628 8300 10656
rect 7699 10625 7711 10628
rect 7653 10619 7711 10625
rect 8294 10616 8300 10628
rect 8352 10616 8358 10668
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 9858 10656 9864 10668
rect 9355 10628 9864 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10137 10659 10195 10665
rect 10137 10656 10149 10659
rect 10008 10628 10149 10656
rect 10008 10616 10014 10628
rect 10137 10625 10149 10628
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 13357 10659 13415 10665
rect 13357 10625 13369 10659
rect 13403 10656 13415 10659
rect 14826 10656 14832 10668
rect 13403 10628 14832 10656
rect 13403 10625 13415 10628
rect 13357 10619 13415 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 14936 10656 14964 10696
rect 15010 10684 15016 10736
rect 15068 10724 15074 10736
rect 15197 10727 15255 10733
rect 15197 10724 15209 10727
rect 15068 10696 15209 10724
rect 15068 10684 15074 10696
rect 15197 10693 15209 10696
rect 15243 10724 15255 10727
rect 18138 10724 18144 10736
rect 15243 10696 18144 10724
rect 15243 10693 15255 10696
rect 15197 10687 15255 10693
rect 18138 10684 18144 10696
rect 18196 10724 18202 10736
rect 18417 10727 18475 10733
rect 18417 10724 18429 10727
rect 18196 10696 18429 10724
rect 18196 10684 18202 10696
rect 18417 10693 18429 10696
rect 18463 10693 18475 10727
rect 18417 10687 18475 10693
rect 15654 10656 15660 10668
rect 14936 10628 15660 10656
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 16114 10656 16120 10668
rect 16075 10628 16120 10656
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 17862 10656 17868 10668
rect 17823 10628 17868 10656
rect 17862 10616 17868 10628
rect 17920 10656 17926 10668
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 17920 10628 18245 10656
rect 17920 10616 17926 10628
rect 18233 10625 18245 10628
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10588 6975 10591
rect 7190 10588 7196 10600
rect 6963 10560 7196 10588
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 7837 10591 7895 10597
rect 7837 10588 7849 10591
rect 7800 10560 7849 10588
rect 7800 10548 7806 10560
rect 7837 10557 7849 10560
rect 7883 10557 7895 10591
rect 7837 10551 7895 10557
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8444 10560 8585 10588
rect 8444 10548 8450 10560
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10557 8723 10591
rect 9490 10588 9496 10600
rect 9451 10560 9496 10588
rect 8665 10551 8723 10557
rect 3878 10480 3884 10532
rect 3936 10520 3942 10532
rect 6365 10523 6423 10529
rect 6365 10520 6377 10523
rect 3936 10492 6377 10520
rect 3936 10480 3942 10492
rect 6365 10489 6377 10492
rect 6411 10489 6423 10523
rect 6365 10483 6423 10489
rect 7006 10480 7012 10532
rect 7064 10520 7070 10532
rect 8680 10520 8708 10551
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 10318 10588 10324 10600
rect 10279 10560 10324 10588
rect 10318 10548 10324 10560
rect 10376 10548 10382 10600
rect 11977 10591 12035 10597
rect 11977 10557 11989 10591
rect 12023 10557 12035 10591
rect 11977 10551 12035 10557
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 12986 10588 12992 10600
rect 12207 10560 12992 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 7064 10492 8708 10520
rect 7064 10480 7070 10492
rect 9398 10480 9404 10532
rect 9456 10520 9462 10532
rect 11054 10520 11060 10532
rect 9456 10492 11060 10520
rect 9456 10480 9462 10492
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 11992 10520 12020 10551
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10588 13599 10591
rect 13722 10588 13728 10600
rect 13587 10560 13728 10588
rect 13587 10557 13599 10560
rect 13541 10551 13599 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 13872 10560 14565 10588
rect 13872 10548 13878 10560
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 15381 10591 15439 10597
rect 15381 10588 15393 10591
rect 14976 10560 15393 10588
rect 14976 10548 14982 10560
rect 15381 10557 15393 10560
rect 15427 10557 15439 10591
rect 16206 10588 16212 10600
rect 16167 10560 16212 10588
rect 15381 10551 15439 10557
rect 16206 10548 16212 10560
rect 16264 10548 16270 10600
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 17126 10588 17132 10600
rect 16356 10560 16401 10588
rect 17087 10560 17132 10588
rect 16356 10548 16362 10560
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 17221 10591 17279 10597
rect 17221 10557 17233 10591
rect 17267 10588 17279 10591
rect 17586 10588 17592 10600
rect 17267 10560 17592 10588
rect 17267 10557 17279 10560
rect 17221 10551 17279 10557
rect 12437 10523 12495 10529
rect 12437 10520 12449 10523
rect 11992 10492 12449 10520
rect 12437 10489 12449 10492
rect 12483 10520 12495 10523
rect 15286 10520 15292 10532
rect 12483 10492 15292 10520
rect 12483 10489 12495 10492
rect 12437 10483 12495 10489
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 2406 10452 2412 10464
rect 2367 10424 2412 10452
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 5534 10452 5540 10464
rect 5495 10424 5540 10452
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 6972 10424 7297 10452
rect 6972 10412 6978 10424
rect 7285 10421 7297 10424
rect 7331 10421 7343 10455
rect 7285 10415 7343 10421
rect 7558 10412 7564 10464
rect 7616 10452 7622 10464
rect 8202 10452 8208 10464
rect 7616 10424 8208 10452
rect 7616 10412 7622 10424
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8478 10412 8484 10464
rect 8536 10452 8542 10464
rect 9769 10455 9827 10461
rect 9769 10452 9781 10455
rect 8536 10424 9781 10452
rect 8536 10412 8542 10424
rect 9769 10421 9781 10424
rect 9815 10421 9827 10455
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 9769 10415 9827 10421
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 12618 10452 12624 10464
rect 12579 10424 12624 10452
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 13998 10452 14004 10464
rect 13959 10424 14004 10452
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 14829 10455 14887 10461
rect 14829 10452 14841 10455
rect 14516 10424 14841 10452
rect 14516 10412 14522 10424
rect 14829 10421 14841 10424
rect 14875 10421 14887 10455
rect 14829 10415 14887 10421
rect 15102 10412 15108 10464
rect 15160 10452 15166 10464
rect 17236 10452 17264 10551
rect 17586 10548 17592 10560
rect 17644 10548 17650 10600
rect 18049 10523 18107 10529
rect 18049 10489 18061 10523
rect 18095 10520 18107 10523
rect 18782 10520 18788 10532
rect 18095 10492 18788 10520
rect 18095 10489 18107 10492
rect 18049 10483 18107 10489
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 18966 10480 18972 10532
rect 19024 10520 19030 10532
rect 19242 10520 19248 10532
rect 19024 10492 19248 10520
rect 19024 10480 19030 10492
rect 19242 10480 19248 10492
rect 19300 10480 19306 10532
rect 15160 10424 17264 10452
rect 15160 10412 15166 10424
rect 1104 10362 18860 10384
rect 1104 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 3430 10362
rect 3482 10310 7622 10362
rect 7674 10310 7686 10362
rect 7738 10310 7750 10362
rect 7802 10310 7814 10362
rect 7866 10310 7878 10362
rect 7930 10310 12070 10362
rect 12122 10310 12134 10362
rect 12186 10310 12198 10362
rect 12250 10310 12262 10362
rect 12314 10310 12326 10362
rect 12378 10310 16518 10362
rect 16570 10310 16582 10362
rect 16634 10310 16646 10362
rect 16698 10310 16710 10362
rect 16762 10310 16774 10362
rect 16826 10310 18860 10362
rect 1104 10288 18860 10310
rect 2222 10248 2228 10260
rect 2183 10220 2228 10248
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 2593 10251 2651 10257
rect 2593 10217 2605 10251
rect 2639 10248 2651 10251
rect 2774 10248 2780 10260
rect 2639 10220 2780 10248
rect 2639 10217 2651 10220
rect 2593 10211 2651 10217
rect 2774 10208 2780 10220
rect 2832 10208 2838 10260
rect 3973 10251 4031 10257
rect 3973 10217 3985 10251
rect 4019 10248 4031 10251
rect 4246 10248 4252 10260
rect 4019 10220 4252 10248
rect 4019 10217 4031 10220
rect 3973 10211 4031 10217
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 5868 10220 7328 10248
rect 5868 10208 5874 10220
rect 3694 10140 3700 10192
rect 3752 10180 3758 10192
rect 4801 10183 4859 10189
rect 4801 10180 4813 10183
rect 3752 10152 4813 10180
rect 3752 10140 3758 10152
rect 4801 10149 4813 10152
rect 4847 10149 4859 10183
rect 4801 10143 4859 10149
rect 6362 10140 6368 10192
rect 6420 10180 6426 10192
rect 7300 10180 7328 10220
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 7432 10220 7665 10248
rect 7432 10208 7438 10220
rect 7653 10217 7665 10220
rect 7699 10217 7711 10251
rect 7653 10211 7711 10217
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 8202 10248 8208 10260
rect 7800 10220 8208 10248
rect 7800 10208 7806 10220
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 9858 10208 9864 10260
rect 9916 10248 9922 10260
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 9916 10220 10149 10248
rect 9916 10208 9922 10220
rect 10137 10217 10149 10220
rect 10183 10248 10195 10251
rect 10962 10248 10968 10260
rect 10183 10220 10968 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 17313 10251 17371 10257
rect 17313 10248 17325 10251
rect 11112 10220 17325 10248
rect 11112 10208 11118 10220
rect 17313 10217 17325 10220
rect 17359 10217 17371 10251
rect 17313 10211 17371 10217
rect 7469 10183 7527 10189
rect 7469 10180 7481 10183
rect 6420 10152 7052 10180
rect 7300 10152 7481 10180
rect 6420 10140 6426 10152
rect 3050 10072 3056 10124
rect 3108 10112 3114 10124
rect 3789 10115 3847 10121
rect 3789 10112 3801 10115
rect 3108 10084 3801 10112
rect 3108 10072 3114 10084
rect 3789 10081 3801 10084
rect 3835 10081 3847 10115
rect 3789 10075 3847 10081
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10044 2099 10047
rect 2222 10044 2228 10056
rect 2087 10016 2228 10044
rect 2087 10013 2099 10016
rect 2041 10007 2099 10013
rect 2222 10004 2228 10016
rect 2280 10004 2286 10056
rect 3804 9976 3832 10075
rect 4430 10072 4436 10124
rect 4488 10112 4494 10124
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 4488 10084 4537 10112
rect 4488 10072 4494 10084
rect 4525 10081 4537 10084
rect 4571 10081 4583 10115
rect 5258 10112 5264 10124
rect 5219 10084 5264 10112
rect 4525 10075 4583 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 5442 10112 5448 10124
rect 5403 10084 5448 10112
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 6270 10112 6276 10124
rect 6231 10084 6276 10112
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 7024 10112 7052 10152
rect 7469 10149 7481 10152
rect 7515 10180 7527 10183
rect 8294 10180 8300 10192
rect 7515 10152 8300 10180
rect 7515 10149 7527 10152
rect 7469 10143 7527 10149
rect 8294 10140 8300 10152
rect 8352 10180 8358 10192
rect 10410 10180 10416 10192
rect 8352 10152 10416 10180
rect 8352 10140 8358 10152
rect 10410 10140 10416 10152
rect 10468 10140 10474 10192
rect 10520 10152 11744 10180
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 6512 10084 6592 10112
rect 7024 10084 7113 10112
rect 6512 10072 6518 10084
rect 4341 10047 4399 10053
rect 4341 10013 4353 10047
rect 4387 10044 4399 10047
rect 4890 10044 4896 10056
rect 4387 10016 4896 10044
rect 4387 10013 4399 10016
rect 4341 10007 4399 10013
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 5626 10004 5632 10056
rect 5684 10044 5690 10056
rect 5994 10044 6000 10056
rect 5684 10016 6000 10044
rect 5684 10004 5690 10016
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6564 10044 6592 10084
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 7374 10072 7380 10124
rect 7432 10112 7438 10124
rect 8110 10112 8116 10124
rect 7432 10084 8116 10112
rect 7432 10072 7438 10084
rect 8110 10072 8116 10084
rect 8168 10112 8174 10124
rect 8205 10115 8263 10121
rect 8205 10112 8217 10115
rect 8168 10084 8217 10112
rect 8168 10072 8174 10084
rect 8205 10081 8217 10084
rect 8251 10081 8263 10115
rect 8205 10075 8263 10081
rect 8386 10072 8392 10124
rect 8444 10072 8450 10124
rect 9306 10072 9312 10124
rect 9364 10112 9370 10124
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 9364 10084 9505 10112
rect 9364 10072 9370 10084
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9950 10112 9956 10124
rect 9911 10084 9956 10112
rect 9493 10075 9551 10081
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 10520 10121 10548 10152
rect 11716 10124 11744 10152
rect 11790 10140 11796 10192
rect 11848 10180 11854 10192
rect 11848 10152 13492 10180
rect 11848 10140 11854 10152
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10081 10563 10115
rect 10505 10075 10563 10081
rect 10597 10115 10655 10121
rect 10597 10081 10609 10115
rect 10643 10112 10655 10115
rect 11514 10112 11520 10124
rect 10643 10084 11520 10112
rect 10643 10081 10655 10084
rect 10597 10075 10655 10081
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 11698 10072 11704 10124
rect 11756 10112 11762 10124
rect 12713 10115 12771 10121
rect 11756 10084 11849 10112
rect 11756 10072 11762 10084
rect 12713 10081 12725 10115
rect 12759 10112 12771 10115
rect 12986 10112 12992 10124
rect 12759 10084 12992 10112
rect 12759 10081 12771 10084
rect 12713 10075 12771 10081
rect 12986 10072 12992 10084
rect 13044 10072 13050 10124
rect 13464 10121 13492 10152
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10081 13507 10115
rect 13449 10075 13507 10081
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 14645 10115 14703 10121
rect 14645 10112 14657 10115
rect 13964 10084 14657 10112
rect 13964 10072 13970 10084
rect 14645 10081 14657 10084
rect 14691 10081 14703 10115
rect 14645 10075 14703 10081
rect 14918 10072 14924 10124
rect 14976 10112 14982 10124
rect 15473 10115 15531 10121
rect 15473 10112 15485 10115
rect 14976 10084 15485 10112
rect 14976 10072 14982 10084
rect 15473 10081 15485 10084
rect 15519 10081 15531 10115
rect 15473 10075 15531 10081
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 16301 10115 16359 10121
rect 16301 10112 16313 10115
rect 15620 10084 16313 10112
rect 15620 10072 15626 10084
rect 16301 10081 16313 10084
rect 16347 10081 16359 10115
rect 16574 10112 16580 10124
rect 16535 10084 16580 10112
rect 16301 10075 16359 10081
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 16758 10072 16764 10124
rect 16816 10112 16822 10124
rect 17037 10115 17095 10121
rect 17037 10112 17049 10115
rect 16816 10084 17049 10112
rect 16816 10072 16822 10084
rect 17037 10081 17049 10084
rect 17083 10081 17095 10115
rect 17037 10075 17095 10081
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6564 10016 6837 10044
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 8404 10044 8432 10072
rect 8481 10047 8539 10053
rect 8481 10044 8493 10047
rect 6825 10007 6883 10013
rect 7668 10016 8493 10044
rect 4433 9979 4491 9985
rect 4433 9976 4445 9979
rect 3804 9948 4445 9976
rect 4433 9945 4445 9948
rect 4479 9945 4491 9979
rect 4433 9939 4491 9945
rect 1762 9868 1768 9920
rect 1820 9908 1826 9920
rect 1857 9911 1915 9917
rect 1857 9908 1869 9911
rect 1820 9880 1869 9908
rect 1820 9868 1826 9880
rect 1857 9877 1869 9880
rect 1903 9877 1915 9911
rect 4448 9908 4476 9939
rect 4522 9936 4528 9988
rect 4580 9976 4586 9988
rect 5534 9976 5540 9988
rect 4580 9948 5540 9976
rect 4580 9936 4586 9948
rect 5534 9936 5540 9948
rect 5592 9976 5598 9988
rect 6089 9979 6147 9985
rect 6089 9976 6101 9979
rect 5592 9948 6101 9976
rect 5592 9936 5598 9948
rect 6089 9945 6101 9948
rect 6135 9945 6147 9979
rect 6089 9939 6147 9945
rect 7190 9936 7196 9988
rect 7248 9976 7254 9988
rect 7668 9976 7696 10016
rect 8481 10013 8493 10016
rect 8527 10013 8539 10047
rect 8481 10007 8539 10013
rect 7248 9948 7696 9976
rect 8021 9979 8079 9985
rect 7248 9936 7254 9948
rect 8021 9945 8033 9979
rect 8067 9976 8079 9979
rect 8386 9976 8392 9988
rect 8067 9948 8392 9976
rect 8067 9945 8079 9948
rect 8021 9939 8079 9945
rect 8386 9936 8392 9948
rect 8444 9936 8450 9988
rect 8496 9976 8524 10007
rect 8662 10004 8668 10056
rect 8720 10044 8726 10056
rect 9214 10044 9220 10056
rect 8720 10016 9220 10044
rect 8720 10004 8726 10016
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 9674 10044 9680 10056
rect 9447 10016 9680 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10044 10747 10047
rect 12342 10044 12348 10056
rect 10735 10016 12348 10044
rect 10735 10013 10747 10016
rect 10689 10007 10747 10013
rect 12342 10004 12348 10016
rect 12400 10004 12406 10056
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10044 13323 10047
rect 13538 10044 13544 10056
rect 13311 10016 13544 10044
rect 13311 10013 13323 10016
rect 13265 10007 13323 10013
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 14458 10044 14464 10056
rect 14419 10016 14464 10044
rect 14458 10004 14464 10016
rect 14516 10004 14522 10056
rect 17328 10044 17356 10211
rect 17681 10183 17739 10189
rect 17681 10149 17693 10183
rect 17727 10180 17739 10183
rect 18966 10180 18972 10192
rect 17727 10152 18972 10180
rect 17727 10149 17739 10152
rect 17681 10143 17739 10149
rect 18966 10140 18972 10152
rect 19024 10140 19030 10192
rect 17497 10047 17555 10053
rect 17497 10044 17509 10047
rect 14752 10016 16804 10044
rect 17328 10016 17509 10044
rect 11238 9976 11244 9988
rect 8496 9948 11244 9976
rect 11238 9936 11244 9948
rect 11296 9936 11302 9988
rect 11517 9979 11575 9985
rect 11517 9945 11529 9979
rect 11563 9976 11575 9979
rect 12437 9979 12495 9985
rect 11563 9948 12112 9976
rect 11563 9945 11575 9948
rect 11517 9939 11575 9945
rect 5074 9908 5080 9920
rect 4448 9880 5080 9908
rect 1857 9871 1915 9877
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5629 9911 5687 9917
rect 5629 9877 5641 9911
rect 5675 9908 5687 9911
rect 5718 9908 5724 9920
rect 5675 9880 5724 9908
rect 5675 9877 5687 9880
rect 5629 9871 5687 9877
rect 5718 9868 5724 9880
rect 5776 9868 5782 9920
rect 6454 9908 6460 9920
rect 6415 9880 6460 9908
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7377 9911 7435 9917
rect 6972 9880 7017 9908
rect 6972 9868 6978 9880
rect 7377 9877 7389 9911
rect 7423 9908 7435 9911
rect 7558 9908 7564 9920
rect 7423 9880 7564 9908
rect 7423 9877 7435 9880
rect 7377 9871 7435 9877
rect 7558 9868 7564 9880
rect 7616 9908 7622 9920
rect 7742 9908 7748 9920
rect 7616 9880 7748 9908
rect 7616 9868 7622 9880
rect 7742 9868 7748 9880
rect 7800 9868 7806 9920
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 8113 9911 8171 9917
rect 8113 9908 8125 9911
rect 7892 9880 8125 9908
rect 7892 9868 7898 9880
rect 8113 9877 8125 9880
rect 8159 9877 8171 9911
rect 8113 9871 8171 9877
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 8662 9908 8668 9920
rect 8352 9880 8668 9908
rect 8352 9868 8358 9880
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 8938 9908 8944 9920
rect 8899 9880 8944 9908
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 9214 9868 9220 9920
rect 9272 9908 9278 9920
rect 9309 9911 9367 9917
rect 9309 9908 9321 9911
rect 9272 9880 9321 9908
rect 9272 9868 9278 9880
rect 9309 9877 9321 9880
rect 9355 9908 9367 9911
rect 9582 9908 9588 9920
rect 9355 9880 9588 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 11054 9908 11060 9920
rect 11015 9880 11060 9908
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 11606 9908 11612 9920
rect 11204 9880 11249 9908
rect 11567 9880 11612 9908
rect 11204 9868 11210 9880
rect 11606 9868 11612 9880
rect 11664 9868 11670 9920
rect 12084 9917 12112 9948
rect 12437 9945 12449 9979
rect 12483 9976 12495 9979
rect 12618 9976 12624 9988
rect 12483 9948 12624 9976
rect 12483 9945 12495 9948
rect 12437 9939 12495 9945
rect 12618 9936 12624 9948
rect 12676 9976 12682 9988
rect 14752 9976 14780 10016
rect 12676 9948 14780 9976
rect 16209 9979 16267 9985
rect 12676 9936 12682 9948
rect 16209 9945 16221 9979
rect 16255 9976 16267 9979
rect 16666 9976 16672 9988
rect 16255 9948 16672 9976
rect 16255 9945 16267 9948
rect 16209 9939 16267 9945
rect 16666 9936 16672 9948
rect 16724 9936 16730 9988
rect 16776 9976 16804 10016
rect 17497 10013 17509 10016
rect 17543 10013 17555 10047
rect 17497 10007 17555 10013
rect 17865 10047 17923 10053
rect 17865 10013 17877 10047
rect 17911 10044 17923 10047
rect 18046 10044 18052 10056
rect 17911 10016 18052 10044
rect 17911 10013 17923 10016
rect 17865 10007 17923 10013
rect 17880 9976 17908 10007
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 18138 10004 18144 10056
rect 18196 10044 18202 10056
rect 18233 10047 18291 10053
rect 18233 10044 18245 10047
rect 18196 10016 18245 10044
rect 18196 10004 18202 10016
rect 18233 10013 18245 10016
rect 18279 10013 18291 10047
rect 18233 10007 18291 10013
rect 16776 9948 17908 9976
rect 12069 9911 12127 9917
rect 12069 9877 12081 9911
rect 12115 9877 12127 9911
rect 12069 9871 12127 9877
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 12894 9908 12900 9920
rect 12584 9880 12629 9908
rect 12855 9880 12900 9908
rect 12584 9868 12590 9880
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 13357 9911 13415 9917
rect 13357 9877 13369 9911
rect 13403 9908 13415 9911
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 13403 9880 14105 9908
rect 13403 9877 13415 9880
rect 13357 9871 13415 9877
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 14093 9871 14151 9877
rect 14553 9911 14611 9917
rect 14553 9877 14565 9911
rect 14599 9908 14611 9911
rect 14921 9911 14979 9917
rect 14921 9908 14933 9911
rect 14599 9880 14933 9908
rect 14599 9877 14611 9880
rect 14553 9871 14611 9877
rect 14921 9877 14933 9880
rect 14967 9877 14979 9911
rect 14921 9871 14979 9877
rect 15010 9868 15016 9920
rect 15068 9908 15074 9920
rect 15289 9911 15347 9917
rect 15289 9908 15301 9911
rect 15068 9880 15301 9908
rect 15068 9868 15074 9880
rect 15289 9877 15301 9880
rect 15335 9877 15347 9911
rect 15289 9871 15347 9877
rect 15378 9868 15384 9920
rect 15436 9908 15442 9920
rect 15746 9908 15752 9920
rect 15436 9880 15481 9908
rect 15707 9880 15752 9908
rect 15436 9868 15442 9880
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 16117 9911 16175 9917
rect 16117 9877 16129 9911
rect 16163 9908 16175 9911
rect 16853 9911 16911 9917
rect 16853 9908 16865 9911
rect 16163 9880 16865 9908
rect 16163 9877 16175 9880
rect 16117 9871 16175 9877
rect 16853 9877 16865 9880
rect 16899 9908 16911 9911
rect 17402 9908 17408 9920
rect 16899 9880 17408 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 17402 9868 17408 9880
rect 17460 9868 17466 9920
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 18049 9911 18107 9917
rect 18049 9908 18061 9911
rect 18012 9880 18061 9908
rect 18012 9868 18018 9880
rect 18049 9877 18061 9880
rect 18095 9877 18107 9911
rect 18049 9871 18107 9877
rect 18417 9911 18475 9917
rect 18417 9877 18429 9911
rect 18463 9908 18475 9911
rect 18598 9908 18604 9920
rect 18463 9880 18604 9908
rect 18463 9877 18475 9880
rect 18417 9871 18475 9877
rect 18598 9868 18604 9880
rect 18656 9868 18662 9920
rect 1104 9818 18860 9840
rect 1104 9766 5398 9818
rect 5450 9766 5462 9818
rect 5514 9766 5526 9818
rect 5578 9766 5590 9818
rect 5642 9766 5654 9818
rect 5706 9766 9846 9818
rect 9898 9766 9910 9818
rect 9962 9766 9974 9818
rect 10026 9766 10038 9818
rect 10090 9766 10102 9818
rect 10154 9766 14294 9818
rect 14346 9766 14358 9818
rect 14410 9766 14422 9818
rect 14474 9766 14486 9818
rect 14538 9766 14550 9818
rect 14602 9766 18860 9818
rect 1104 9744 18860 9766
rect 2225 9707 2283 9713
rect 2225 9673 2237 9707
rect 2271 9704 2283 9707
rect 2406 9704 2412 9716
rect 2271 9676 2412 9704
rect 2271 9673 2283 9676
rect 2225 9667 2283 9673
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 4338 9704 4344 9716
rect 4299 9676 4344 9704
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 5629 9707 5687 9713
rect 5629 9673 5641 9707
rect 5675 9704 5687 9707
rect 5718 9704 5724 9716
rect 5675 9676 5724 9704
rect 5675 9673 5687 9676
rect 5629 9667 5687 9673
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6089 9707 6147 9713
rect 6089 9704 6101 9707
rect 6052 9676 6101 9704
rect 6052 9664 6058 9676
rect 6089 9673 6101 9676
rect 6135 9673 6147 9707
rect 6089 9667 6147 9673
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6512 9676 6837 9704
rect 6512 9664 6518 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 6825 9667 6883 9673
rect 7834 9664 7840 9716
rect 7892 9704 7898 9716
rect 7929 9707 7987 9713
rect 7929 9704 7941 9707
rect 7892 9676 7941 9704
rect 7892 9664 7898 9676
rect 7929 9673 7941 9676
rect 7975 9673 7987 9707
rect 8297 9707 8355 9713
rect 8297 9704 8309 9707
rect 7929 9667 7987 9673
rect 8128 9676 8309 9704
rect 3142 9636 3148 9648
rect 2792 9608 3148 9636
rect 2792 9577 2820 9608
rect 3142 9596 3148 9608
rect 3200 9596 3206 9648
rect 3513 9639 3571 9645
rect 3513 9605 3525 9639
rect 3559 9636 3571 9639
rect 3602 9636 3608 9648
rect 3559 9608 3608 9636
rect 3559 9605 3571 9608
rect 3513 9599 3571 9605
rect 3602 9596 3608 9608
rect 3660 9596 3666 9648
rect 4522 9596 4528 9648
rect 4580 9596 4586 9648
rect 5810 9596 5816 9648
rect 5868 9596 5874 9648
rect 5902 9596 5908 9648
rect 5960 9636 5966 9648
rect 6733 9639 6791 9645
rect 6733 9636 6745 9639
rect 5960 9608 6745 9636
rect 5960 9596 5966 9608
rect 6733 9605 6745 9608
rect 6779 9605 6791 9639
rect 6733 9599 6791 9605
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 7558 9636 7564 9648
rect 6972 9608 7564 9636
rect 6972 9596 6978 9608
rect 7558 9596 7564 9608
rect 7616 9596 7622 9648
rect 8128 9636 8156 9676
rect 8297 9673 8309 9676
rect 8343 9704 8355 9707
rect 9030 9704 9036 9716
rect 8343 9676 9036 9704
rect 8343 9673 8355 9676
rect 8297 9667 8355 9673
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 9858 9704 9864 9716
rect 9819 9676 9864 9704
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 11149 9707 11207 9713
rect 11149 9673 11161 9707
rect 11195 9704 11207 9707
rect 11606 9704 11612 9716
rect 11195 9676 11612 9704
rect 11195 9673 11207 9676
rect 11149 9667 11207 9673
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 11885 9707 11943 9713
rect 11885 9673 11897 9707
rect 11931 9704 11943 9707
rect 12158 9704 12164 9716
rect 11931 9676 12164 9704
rect 11931 9673 11943 9676
rect 11885 9667 11943 9673
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12342 9704 12348 9716
rect 12303 9676 12348 9704
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 13173 9707 13231 9713
rect 13173 9704 13185 9707
rect 12584 9676 13185 9704
rect 12584 9664 12590 9676
rect 13173 9673 13185 9676
rect 13219 9673 13231 9707
rect 13538 9704 13544 9716
rect 13451 9676 13544 9704
rect 13173 9667 13231 9673
rect 13538 9664 13544 9676
rect 13596 9704 13602 9716
rect 14642 9704 14648 9716
rect 13596 9676 14648 9704
rect 13596 9664 13602 9676
rect 14642 9664 14648 9676
rect 14700 9664 14706 9716
rect 14826 9704 14832 9716
rect 14787 9676 14832 9704
rect 14826 9664 14832 9676
rect 14884 9664 14890 9716
rect 15197 9707 15255 9713
rect 15197 9673 15209 9707
rect 15243 9704 15255 9707
rect 15746 9704 15752 9716
rect 15243 9676 15752 9704
rect 15243 9673 15255 9676
rect 15197 9667 15255 9673
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 16666 9704 16672 9716
rect 16627 9676 16672 9704
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 17862 9704 17868 9716
rect 17823 9676 17868 9704
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 18046 9664 18052 9716
rect 18104 9704 18110 9716
rect 18325 9707 18383 9713
rect 18325 9704 18337 9707
rect 18104 9676 18337 9704
rect 18104 9664 18110 9676
rect 18325 9673 18337 9676
rect 18371 9673 18383 9707
rect 18325 9667 18383 9673
rect 7852 9608 8156 9636
rect 9125 9639 9183 9645
rect 2777 9571 2835 9577
rect 2777 9568 2789 9571
rect 1964 9540 2789 9568
rect 1964 9509 1992 9540
rect 2777 9537 2789 9540
rect 2823 9537 2835 9571
rect 2777 9531 2835 9537
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 4433 9571 4491 9577
rect 4433 9568 4445 9571
rect 2924 9540 4445 9568
rect 2924 9528 2930 9540
rect 4433 9537 4445 9540
rect 4479 9568 4491 9571
rect 4540 9568 4568 9596
rect 5074 9568 5080 9580
rect 4479 9540 4568 9568
rect 4987 9540 5080 9568
rect 4479 9537 4491 9540
rect 4433 9531 4491 9537
rect 5074 9528 5080 9540
rect 5132 9568 5138 9580
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5132 9540 5549 9568
rect 5132 9528 5138 9540
rect 5537 9537 5549 9540
rect 5583 9568 5595 9571
rect 5828 9568 5856 9596
rect 7650 9568 7656 9580
rect 5583 9540 5856 9568
rect 7611 9540 7656 9568
rect 5583 9537 5595 9540
rect 5537 9531 5595 9537
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7852 9577 7880 9608
rect 9125 9605 9137 9639
rect 9171 9636 9183 9639
rect 9214 9636 9220 9648
rect 9171 9608 9220 9636
rect 9171 9605 9183 9608
rect 9125 9599 9183 9605
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 10318 9636 10324 9648
rect 9600 9608 10324 9636
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9537 7895 9571
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 7837 9531 7895 9537
rect 8036 9540 8401 9568
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9469 2007 9503
rect 1949 9463 2007 9469
rect 2038 9460 2044 9512
rect 2096 9500 2102 9512
rect 2133 9503 2191 9509
rect 2133 9500 2145 9503
rect 2096 9472 2145 9500
rect 2096 9460 2102 9472
rect 2133 9469 2145 9472
rect 2179 9469 2191 9503
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 2133 9463 2191 9469
rect 2746 9472 3617 9500
rect 2593 9435 2651 9441
rect 2593 9401 2605 9435
rect 2639 9432 2651 9435
rect 2746 9432 2774 9472
rect 3605 9469 3617 9472
rect 3651 9469 3663 9503
rect 3605 9463 3663 9469
rect 3789 9503 3847 9509
rect 3789 9469 3801 9503
rect 3835 9500 3847 9503
rect 4062 9500 4068 9512
rect 3835 9472 4068 9500
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 4338 9460 4344 9512
rect 4396 9500 4402 9512
rect 4525 9503 4583 9509
rect 4525 9500 4537 9503
rect 4396 9472 4537 9500
rect 4396 9460 4402 9472
rect 4525 9469 4537 9472
rect 4571 9469 4583 9503
rect 4525 9463 4583 9469
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9500 5871 9503
rect 6454 9500 6460 9512
rect 5859 9472 6460 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 6454 9460 6460 9472
rect 6512 9460 6518 9512
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6696 9472 6929 9500
rect 6696 9460 6702 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 2639 9404 2774 9432
rect 2639 9401 2651 9404
rect 2593 9395 2651 9401
rect 2866 9392 2872 9444
rect 2924 9432 2930 9444
rect 2961 9435 3019 9441
rect 2961 9432 2973 9435
rect 2924 9404 2973 9432
rect 2924 9392 2930 9404
rect 2961 9401 2973 9404
rect 3007 9401 3019 9435
rect 3973 9435 4031 9441
rect 2961 9395 3019 9401
rect 3068 9404 3832 9432
rect 2222 9324 2228 9376
rect 2280 9364 2286 9376
rect 3068 9364 3096 9404
rect 2280 9336 3096 9364
rect 3145 9367 3203 9373
rect 2280 9324 2286 9336
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 3694 9364 3700 9376
rect 3191 9336 3700 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 3804 9364 3832 9404
rect 3973 9401 3985 9435
rect 4019 9432 4031 9435
rect 4154 9432 4160 9444
rect 4019 9404 4160 9432
rect 4019 9401 4031 9404
rect 3973 9395 4031 9401
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 4801 9435 4859 9441
rect 4801 9401 4813 9435
rect 4847 9432 4859 9435
rect 4890 9432 4896 9444
rect 4847 9404 4896 9432
rect 4847 9401 4859 9404
rect 4801 9395 4859 9401
rect 4816 9364 4844 9395
rect 4890 9392 4896 9404
rect 4948 9432 4954 9444
rect 5442 9432 5448 9444
rect 4948 9404 5448 9432
rect 4948 9392 4954 9404
rect 5442 9392 5448 9404
rect 5500 9392 5506 9444
rect 5626 9392 5632 9444
rect 5684 9432 5690 9444
rect 7377 9435 7435 9441
rect 7377 9432 7389 9435
rect 5684 9404 7389 9432
rect 5684 9392 5690 9404
rect 7377 9401 7389 9404
rect 7423 9432 7435 9435
rect 8036 9432 8064 9540
rect 8389 9537 8401 9540
rect 8435 9568 8447 9571
rect 9600 9568 9628 9608
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 11333 9639 11391 9645
rect 11333 9636 11345 9639
rect 10428 9608 11345 9636
rect 9950 9568 9956 9580
rect 8435 9540 9352 9568
rect 8435 9537 8447 9540
rect 8389 9531 8447 9537
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 8662 9500 8668 9512
rect 8619 9472 8668 9500
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 8662 9460 8668 9472
rect 8720 9500 8726 9512
rect 9214 9500 9220 9512
rect 8720 9472 8984 9500
rect 9175 9472 9220 9500
rect 8720 9460 8726 9472
rect 7423 9404 8064 9432
rect 7423 9401 7435 9404
rect 7377 9395 7435 9401
rect 5166 9364 5172 9376
rect 3804 9336 4844 9364
rect 5127 9336 5172 9364
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 6328 9336 6377 9364
rect 6328 9324 6334 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 6604 9336 7205 9364
rect 6604 9324 6610 9336
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 7193 9327 7251 9333
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 8294 9364 8300 9376
rect 7616 9336 8300 9364
rect 7616 9324 7622 9336
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 8754 9324 8760 9376
rect 8812 9364 8818 9376
rect 8956 9364 8984 9472
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 9324 9432 9352 9540
rect 9508 9540 9628 9568
rect 9911 9540 9956 9568
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 9508 9500 9536 9540
rect 9950 9528 9956 9540
rect 10008 9528 10014 9580
rect 9447 9472 9536 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 10428 9500 10456 9608
rect 11333 9605 11345 9608
rect 11379 9636 11391 9639
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 11379 9608 11989 9636
rect 11379 9605 11391 9608
rect 11333 9599 11391 9605
rect 11977 9605 11989 9608
rect 12023 9605 12035 9639
rect 14366 9636 14372 9648
rect 11977 9599 12035 9605
rect 12084 9608 13759 9636
rect 14279 9608 14372 9636
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 9824 9472 9869 9500
rect 10244 9472 10456 9500
rect 10520 9540 10793 9568
rect 9824 9460 9830 9472
rect 10244 9432 10272 9472
rect 9324 9404 10272 9432
rect 10321 9435 10379 9441
rect 10321 9401 10333 9435
rect 10367 9432 10379 9435
rect 10520 9432 10548 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10597 9503 10655 9509
rect 10597 9469 10609 9503
rect 10643 9469 10655 9503
rect 10597 9463 10655 9469
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9500 10747 9503
rect 10735 9472 11560 9500
rect 10735 9469 10747 9472
rect 10689 9463 10747 9469
rect 10367 9404 10548 9432
rect 10367 9401 10379 9404
rect 10321 9395 10379 9401
rect 9490 9364 9496 9376
rect 8812 9336 8857 9364
rect 8956 9336 9496 9364
rect 8812 9324 8818 9336
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 10612 9364 10640 9463
rect 11532 9441 11560 9472
rect 11517 9435 11575 9441
rect 11517 9401 11529 9435
rect 11563 9401 11575 9435
rect 11992 9432 12020 9599
rect 12084 9512 12112 9608
rect 12710 9568 12716 9580
rect 12671 9540 12716 9568
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 12805 9571 12863 9577
rect 12805 9537 12817 9571
rect 12851 9568 12863 9571
rect 13262 9568 13268 9580
rect 12851 9540 13268 9568
rect 12851 9537 12863 9540
rect 12805 9531 12863 9537
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 12066 9460 12072 9512
rect 12124 9500 12130 9512
rect 12894 9500 12900 9512
rect 12124 9472 12169 9500
rect 12855 9472 12900 9500
rect 12124 9460 12130 9472
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 12986 9460 12992 9512
rect 13044 9500 13050 9512
rect 13731 9509 13759 9608
rect 14366 9596 14372 9608
rect 14424 9636 14430 9648
rect 15286 9636 15292 9648
rect 14424 9608 15292 9636
rect 14424 9596 14430 9608
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 15470 9596 15476 9648
rect 15528 9636 15534 9648
rect 15930 9636 15936 9648
rect 15528 9608 15936 9636
rect 15528 9596 15534 9608
rect 15930 9596 15936 9608
rect 15988 9596 15994 9648
rect 16025 9639 16083 9645
rect 16025 9605 16037 9639
rect 16071 9636 16083 9639
rect 16574 9636 16580 9648
rect 16071 9608 16580 9636
rect 16071 9605 16083 9608
rect 16025 9599 16083 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 17034 9636 17040 9648
rect 16995 9608 17040 9636
rect 17034 9596 17040 9608
rect 17092 9636 17098 9648
rect 17586 9636 17592 9648
rect 17092 9608 17592 9636
rect 17092 9596 17098 9608
rect 17586 9596 17592 9608
rect 17644 9596 17650 9648
rect 17770 9568 17776 9580
rect 14660 9540 17776 9568
rect 13633 9503 13691 9509
rect 13633 9500 13645 9503
rect 13044 9472 13645 9500
rect 13044 9460 13050 9472
rect 13633 9469 13645 9472
rect 13679 9469 13691 9503
rect 13633 9463 13691 9469
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9469 13783 9503
rect 14090 9500 14096 9512
rect 14051 9472 14096 9500
rect 13725 9463 13783 9469
rect 14090 9460 14096 9472
rect 14148 9460 14154 9512
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 14277 9503 14335 9509
rect 14277 9500 14289 9503
rect 14240 9472 14289 9500
rect 14240 9460 14246 9472
rect 14277 9469 14289 9472
rect 14323 9469 14335 9503
rect 14277 9463 14335 9469
rect 12618 9432 12624 9444
rect 11992 9404 12624 9432
rect 11517 9395 11575 9401
rect 12618 9392 12624 9404
rect 12676 9432 12682 9444
rect 14660 9432 14688 9540
rect 17770 9528 17776 9540
rect 17828 9568 17834 9580
rect 17828 9540 17908 9568
rect 17828 9528 17834 9540
rect 14826 9460 14832 9512
rect 14884 9500 14890 9512
rect 15289 9503 15347 9509
rect 15289 9500 15301 9503
rect 14884 9472 15301 9500
rect 14884 9460 14890 9472
rect 15289 9469 15301 9472
rect 15335 9469 15347 9503
rect 15289 9463 15347 9469
rect 15381 9503 15439 9509
rect 15381 9469 15393 9503
rect 15427 9469 15439 9503
rect 15381 9463 15439 9469
rect 12676 9404 14688 9432
rect 14737 9435 14795 9441
rect 12676 9392 12682 9404
rect 14737 9401 14749 9435
rect 14783 9432 14795 9435
rect 15010 9432 15016 9444
rect 14783 9404 15016 9432
rect 14783 9401 14795 9404
rect 14737 9395 14795 9401
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 11882 9364 11888 9376
rect 10612 9336 11888 9364
rect 11882 9324 11888 9336
rect 11940 9364 11946 9376
rect 12894 9364 12900 9376
rect 11940 9336 12900 9364
rect 11940 9324 11946 9336
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13630 9324 13636 9376
rect 13688 9364 13694 9376
rect 14642 9364 14648 9376
rect 13688 9336 14648 9364
rect 13688 9324 13694 9336
rect 14642 9324 14648 9336
rect 14700 9364 14706 9376
rect 15396 9364 15424 9463
rect 15654 9460 15660 9512
rect 15712 9500 15718 9512
rect 15749 9503 15807 9509
rect 15749 9500 15761 9503
rect 15712 9472 15761 9500
rect 15712 9460 15718 9472
rect 15749 9469 15761 9472
rect 15795 9469 15807 9503
rect 15749 9463 15807 9469
rect 16758 9460 16764 9512
rect 16816 9500 16822 9512
rect 17034 9500 17040 9512
rect 16816 9472 17040 9500
rect 16816 9460 16822 9472
rect 17034 9460 17040 9472
rect 17092 9500 17098 9512
rect 17129 9503 17187 9509
rect 17129 9500 17141 9503
rect 17092 9472 17141 9500
rect 17092 9460 17098 9472
rect 17129 9469 17141 9472
rect 17175 9469 17187 9503
rect 17310 9500 17316 9512
rect 17271 9472 17316 9500
rect 17129 9463 17187 9469
rect 17310 9460 17316 9472
rect 17368 9460 17374 9512
rect 17880 9500 17908 9540
rect 17957 9503 18015 9509
rect 17957 9500 17969 9503
rect 17880 9472 17969 9500
rect 17957 9469 17969 9472
rect 18003 9469 18015 9503
rect 17957 9463 18015 9469
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 15470 9392 15476 9444
rect 15528 9432 15534 9444
rect 16022 9432 16028 9444
rect 15528 9404 16028 9432
rect 15528 9392 15534 9404
rect 16022 9392 16028 9404
rect 16080 9392 16086 9444
rect 17328 9432 17356 9460
rect 18064 9432 18092 9463
rect 17328 9404 18092 9432
rect 16390 9364 16396 9376
rect 14700 9336 15424 9364
rect 16351 9336 16396 9364
rect 14700 9324 14706 9336
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 1104 9274 18860 9296
rect 1104 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 3430 9274
rect 3482 9222 7622 9274
rect 7674 9222 7686 9274
rect 7738 9222 7750 9274
rect 7802 9222 7814 9274
rect 7866 9222 7878 9274
rect 7930 9222 12070 9274
rect 12122 9222 12134 9274
rect 12186 9222 12198 9274
rect 12250 9222 12262 9274
rect 12314 9222 12326 9274
rect 12378 9222 16518 9274
rect 16570 9222 16582 9274
rect 16634 9222 16646 9274
rect 16698 9222 16710 9274
rect 16762 9222 16774 9274
rect 16826 9222 18860 9274
rect 1104 9200 18860 9222
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 3145 9163 3203 9169
rect 3145 9160 3157 9163
rect 3016 9132 3157 9160
rect 3016 9120 3022 9132
rect 3145 9129 3157 9132
rect 3191 9160 3203 9163
rect 4982 9160 4988 9172
rect 3191 9132 4988 9160
rect 3191 9129 3203 9132
rect 3145 9123 3203 9129
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 8444 9132 8953 9160
rect 8444 9120 8450 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 8941 9123 8999 9129
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 9732 9132 9904 9160
rect 9732 9120 9738 9132
rect 3970 9092 3976 9104
rect 1872 9064 3976 9092
rect 1872 8965 1900 9064
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 4706 9092 4712 9104
rect 4448 9064 4712 9092
rect 2314 8984 2320 9036
rect 2372 9024 2378 9036
rect 2409 9027 2467 9033
rect 2409 9024 2421 9027
rect 2372 8996 2421 9024
rect 2372 8984 2378 8996
rect 2409 8993 2421 8996
rect 2455 8993 2467 9027
rect 2590 9024 2596 9036
rect 2551 8996 2596 9024
rect 2409 8987 2467 8993
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 4448 9033 4476 9064
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 5902 9052 5908 9104
rect 5960 9092 5966 9104
rect 6178 9092 6184 9104
rect 5960 9064 6184 9092
rect 5960 9052 5966 9064
rect 6178 9052 6184 9064
rect 6236 9052 6242 9104
rect 7929 9095 7987 9101
rect 7929 9061 7941 9095
rect 7975 9092 7987 9095
rect 8662 9092 8668 9104
rect 7975 9064 8668 9092
rect 7975 9061 7987 9064
rect 7929 9055 7987 9061
rect 8662 9052 8668 9064
rect 8720 9052 8726 9104
rect 9876 9101 9904 9132
rect 9950 9120 9956 9172
rect 10008 9160 10014 9172
rect 10505 9163 10563 9169
rect 10505 9160 10517 9163
rect 10008 9132 10517 9160
rect 10008 9120 10014 9132
rect 10505 9129 10517 9132
rect 10551 9160 10563 9163
rect 11609 9163 11667 9169
rect 11609 9160 11621 9163
rect 10551 9132 11621 9160
rect 10551 9129 10563 9132
rect 10505 9123 10563 9129
rect 11609 9129 11621 9132
rect 11655 9160 11667 9163
rect 13446 9160 13452 9172
rect 11655 9132 13452 9160
rect 11655 9129 11667 9132
rect 11609 9123 11667 9129
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 14185 9163 14243 9169
rect 14185 9129 14197 9163
rect 14231 9160 14243 9163
rect 14734 9160 14740 9172
rect 14231 9132 14740 9160
rect 14231 9129 14243 9132
rect 14185 9123 14243 9129
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 14826 9120 14832 9172
rect 14884 9160 14890 9172
rect 15381 9163 15439 9169
rect 15381 9160 15393 9163
rect 14884 9132 15393 9160
rect 14884 9120 14890 9132
rect 15381 9129 15393 9132
rect 15427 9129 15439 9163
rect 17034 9160 17040 9172
rect 15381 9123 15439 9129
rect 15764 9132 17040 9160
rect 9861 9095 9919 9101
rect 9861 9061 9873 9095
rect 9907 9092 9919 9095
rect 11514 9092 11520 9104
rect 9907 9064 11520 9092
rect 9907 9061 9919 9064
rect 9861 9055 9919 9061
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 12434 9092 12440 9104
rect 12347 9064 12440 9092
rect 12434 9052 12440 9064
rect 12492 9092 12498 9104
rect 13354 9092 13360 9104
rect 12492 9064 13360 9092
rect 12492 9052 12498 9064
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 14366 9092 14372 9104
rect 14327 9064 14372 9092
rect 14366 9052 14372 9064
rect 14424 9052 14430 9104
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 8993 4491 9027
rect 4433 8987 4491 8993
rect 4522 8984 4528 9036
rect 4580 9024 4586 9036
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 4580 8996 5181 9024
rect 4580 8984 4586 8996
rect 5169 8993 5181 8996
rect 5215 8993 5227 9027
rect 5534 9024 5540 9036
rect 5495 8996 5540 9024
rect 5169 8987 5227 8993
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 8113 9027 8171 9033
rect 8113 8993 8125 9027
rect 8159 8993 8171 9027
rect 8113 8987 8171 8993
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 9024 8355 9027
rect 8754 9024 8760 9036
rect 8343 8996 8760 9024
rect 8343 8993 8355 8996
rect 8297 8987 8355 8993
rect 1489 8959 1547 8965
rect 1489 8925 1501 8959
rect 1535 8956 1547 8959
rect 1857 8959 1915 8965
rect 1857 8956 1869 8959
rect 1535 8928 1869 8956
rect 1535 8925 1547 8928
rect 1489 8919 1547 8925
rect 1857 8925 1869 8928
rect 1903 8925 1915 8959
rect 1857 8919 1915 8925
rect 3142 8916 3148 8968
rect 3200 8956 3206 8968
rect 3605 8959 3663 8965
rect 3605 8956 3617 8959
rect 3200 8928 3617 8956
rect 3200 8916 3206 8928
rect 3605 8925 3617 8928
rect 3651 8956 3663 8959
rect 4249 8959 4307 8965
rect 4249 8956 4261 8959
rect 3651 8928 4261 8956
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 4249 8925 4261 8928
rect 4295 8956 4307 8959
rect 4614 8956 4620 8968
rect 4295 8928 4620 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 6546 8956 6552 8968
rect 5500 8928 6316 8956
rect 6507 8928 6552 8956
rect 5500 8916 5506 8928
rect 3421 8891 3479 8897
rect 3421 8857 3433 8891
rect 3467 8888 3479 8891
rect 4157 8891 4215 8897
rect 4157 8888 4169 8891
rect 3467 8860 4169 8888
rect 3467 8857 3479 8860
rect 3421 8851 3479 8857
rect 4157 8857 4169 8860
rect 4203 8857 4215 8891
rect 5626 8888 5632 8900
rect 4157 8851 4215 8857
rect 4264 8860 5632 8888
rect 1670 8820 1676 8832
rect 1631 8792 1676 8820
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 2317 8823 2375 8829
rect 2317 8789 2329 8823
rect 2363 8820 2375 8823
rect 2869 8823 2927 8829
rect 2869 8820 2881 8823
rect 2363 8792 2881 8820
rect 2363 8789 2375 8792
rect 2317 8783 2375 8789
rect 2869 8789 2881 8792
rect 2915 8820 2927 8823
rect 2958 8820 2964 8832
rect 2915 8792 2964 8820
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3786 8820 3792 8832
rect 3747 8792 3792 8820
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 4264 8820 4292 8860
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 5810 8888 5816 8900
rect 5771 8860 5816 8888
rect 5810 8848 5816 8860
rect 5868 8848 5874 8900
rect 4028 8792 4292 8820
rect 4028 8780 4034 8792
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 4617 8823 4675 8829
rect 4617 8820 4629 8823
rect 4488 8792 4629 8820
rect 4488 8780 4494 8792
rect 4617 8789 4629 8792
rect 4663 8789 4675 8823
rect 4982 8820 4988 8832
rect 4943 8792 4988 8820
rect 4617 8783 4675 8789
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 5718 8820 5724 8832
rect 5132 8792 5177 8820
rect 5679 8792 5724 8820
rect 5132 8780 5138 8792
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 6178 8820 6184 8832
rect 6139 8792 6184 8820
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 6288 8820 6316 8928
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 6638 8916 6644 8968
rect 6696 8916 6702 8968
rect 6805 8959 6863 8965
rect 6805 8925 6817 8959
rect 6851 8925 6863 8959
rect 8128 8956 8156 8987
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 11146 9024 11152 9036
rect 9548 8996 9593 9024
rect 11107 8996 11152 9024
rect 9548 8984 9554 8996
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 11333 9027 11391 9033
rect 11333 8993 11345 9027
rect 11379 9024 11391 9027
rect 11422 9024 11428 9036
rect 11379 8996 11428 9024
rect 11379 8993 11391 8996
rect 11333 8987 11391 8993
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 9024 12035 9027
rect 12710 9024 12716 9036
rect 12023 8996 12716 9024
rect 12023 8993 12035 8996
rect 11977 8987 12035 8993
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 14090 8984 14096 9036
rect 14148 9024 14154 9036
rect 14645 9027 14703 9033
rect 14645 9024 14657 9027
rect 14148 8996 14657 9024
rect 14148 8984 14154 8996
rect 14645 8993 14657 8996
rect 14691 8993 14703 9027
rect 15764 9024 15792 9132
rect 17034 9120 17040 9132
rect 17092 9120 17098 9172
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 17405 9163 17463 9169
rect 17405 9160 17417 9163
rect 17184 9132 17417 9160
rect 17184 9120 17190 9132
rect 17405 9129 17417 9132
rect 17451 9129 17463 9163
rect 17405 9123 17463 9129
rect 17494 9092 17500 9104
rect 15856 9064 17500 9092
rect 15856 9033 15884 9064
rect 17494 9052 17500 9064
rect 17552 9052 17558 9104
rect 14645 8987 14703 8993
rect 14936 8996 15792 9024
rect 15841 9027 15899 9033
rect 8389 8959 8447 8965
rect 8128 8928 8340 8956
rect 6805 8919 6863 8925
rect 6656 8888 6684 8916
rect 6820 8888 6848 8919
rect 6656 8860 6848 8888
rect 6457 8823 6515 8829
rect 6457 8820 6469 8823
rect 6288 8792 6469 8820
rect 6457 8789 6469 8792
rect 6503 8820 6515 8823
rect 6730 8820 6736 8832
rect 6503 8792 6736 8820
rect 6503 8789 6515 8792
rect 6457 8783 6515 8789
rect 6730 8780 6736 8792
rect 6788 8820 6794 8832
rect 7282 8820 7288 8832
rect 6788 8792 7288 8820
rect 6788 8780 6794 8792
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 8312 8820 8340 8928
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 8478 8956 8484 8968
rect 8435 8928 8484 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 9858 8956 9864 8968
rect 9692 8928 9864 8956
rect 8938 8848 8944 8900
rect 8996 8888 9002 8900
rect 9401 8891 9459 8897
rect 9401 8888 9413 8891
rect 8996 8860 9413 8888
rect 8996 8848 9002 8860
rect 9401 8857 9413 8860
rect 9447 8888 9459 8891
rect 9692 8888 9720 8928
rect 9858 8916 9864 8928
rect 9916 8956 9922 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9916 8928 10149 8956
rect 9916 8916 9922 8928
rect 10137 8925 10149 8928
rect 10183 8956 10195 8959
rect 11054 8956 11060 8968
rect 10183 8928 10824 8956
rect 11015 8928 11060 8956
rect 10183 8925 10195 8928
rect 10137 8919 10195 8925
rect 9447 8860 9720 8888
rect 9447 8857 9459 8860
rect 9401 8851 9459 8857
rect 8478 8820 8484 8832
rect 8312 8792 8484 8820
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 8754 8820 8760 8832
rect 8715 8792 8760 8820
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 9309 8823 9367 8829
rect 9309 8820 9321 8823
rect 8904 8792 9321 8820
rect 8904 8780 8910 8792
rect 9309 8789 9321 8792
rect 9355 8789 9367 8823
rect 9309 8783 9367 8789
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 9950 8820 9956 8832
rect 9640 8792 9956 8820
rect 9640 8780 9646 8792
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 10045 8823 10103 8829
rect 10045 8789 10057 8823
rect 10091 8820 10103 8823
rect 10410 8820 10416 8832
rect 10091 8792 10416 8820
rect 10091 8789 10103 8792
rect 10045 8783 10103 8789
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 10686 8820 10692 8832
rect 10647 8792 10692 8820
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 10796 8820 10824 8928
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 12066 8916 12072 8968
rect 12124 8956 12130 8968
rect 12124 8928 12756 8956
rect 12124 8916 12130 8928
rect 12728 8888 12756 8928
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 14936 8965 14964 8996
rect 15841 8993 15853 9027
rect 15887 8993 15899 9027
rect 15841 8987 15899 8993
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 8993 15991 9027
rect 15933 8987 15991 8993
rect 16761 9027 16819 9033
rect 16761 8993 16773 9027
rect 16807 8993 16819 9027
rect 17957 9027 18015 9033
rect 17957 9024 17969 9027
rect 16761 8987 16819 8993
rect 16960 8996 17969 9024
rect 14921 8959 14979 8965
rect 14921 8956 14933 8959
rect 12860 8928 14933 8956
rect 12860 8916 12866 8928
rect 14921 8925 14933 8928
rect 14967 8925 14979 8959
rect 14921 8919 14979 8925
rect 15562 8916 15568 8968
rect 15620 8956 15626 8968
rect 15948 8956 15976 8987
rect 15620 8928 15976 8956
rect 15620 8916 15626 8928
rect 16390 8916 16396 8968
rect 16448 8956 16454 8968
rect 16577 8959 16635 8965
rect 16577 8956 16589 8959
rect 16448 8928 16589 8956
rect 16448 8916 16454 8928
rect 16577 8925 16589 8928
rect 16623 8925 16635 8959
rect 16776 8956 16804 8987
rect 16850 8956 16856 8968
rect 16776 8928 16856 8956
rect 16577 8919 16635 8925
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 13725 8891 13783 8897
rect 13725 8888 13737 8891
rect 12728 8860 13737 8888
rect 13725 8857 13737 8860
rect 13771 8888 13783 8891
rect 13771 8860 14872 8888
rect 13771 8857 13783 8860
rect 13725 8851 13783 8857
rect 14844 8832 14872 8860
rect 16022 8848 16028 8900
rect 16080 8888 16086 8900
rect 16080 8860 16804 8888
rect 16080 8848 16086 8860
rect 11974 8820 11980 8832
rect 10796 8792 11980 8820
rect 11974 8780 11980 8792
rect 12032 8780 12038 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 12986 8820 12992 8832
rect 12492 8792 12992 8820
rect 12492 8780 12498 8792
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 13262 8820 13268 8832
rect 13223 8792 13268 8820
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 13909 8823 13967 8829
rect 13909 8789 13921 8823
rect 13955 8820 13967 8823
rect 14182 8820 14188 8832
rect 13955 8792 14188 8820
rect 13955 8789 13967 8792
rect 13909 8783 13967 8789
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 14826 8820 14832 8832
rect 14787 8792 14832 8820
rect 14826 8780 14832 8792
rect 14884 8780 14890 8832
rect 15289 8823 15347 8829
rect 15289 8789 15301 8823
rect 15335 8820 15347 8823
rect 15378 8820 15384 8832
rect 15335 8792 15384 8820
rect 15335 8789 15347 8792
rect 15289 8783 15347 8789
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15746 8820 15752 8832
rect 15707 8792 15752 8820
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 16206 8820 16212 8832
rect 16167 8792 16212 8820
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 16632 8792 16681 8820
rect 16632 8780 16638 8792
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 16776 8820 16804 8860
rect 16960 8820 16988 8996
rect 17957 8993 17969 8996
rect 18003 8993 18015 9027
rect 17957 8987 18015 8993
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17678 8956 17684 8968
rect 17092 8928 17684 8956
rect 17092 8916 17098 8928
rect 17678 8916 17684 8928
rect 17736 8956 17742 8968
rect 17773 8959 17831 8965
rect 17773 8956 17785 8959
rect 17736 8928 17785 8956
rect 17736 8916 17742 8928
rect 17773 8925 17785 8928
rect 17819 8925 17831 8959
rect 18230 8956 18236 8968
rect 18191 8928 18236 8956
rect 17773 8919 17831 8925
rect 18230 8916 18236 8928
rect 18288 8916 18294 8968
rect 17126 8848 17132 8900
rect 17184 8888 17190 8900
rect 17221 8891 17279 8897
rect 17221 8888 17233 8891
rect 17184 8860 17233 8888
rect 17184 8848 17190 8860
rect 17221 8857 17233 8860
rect 17267 8857 17279 8891
rect 17221 8851 17279 8857
rect 16776 8792 16988 8820
rect 16669 8783 16727 8789
rect 17034 8780 17040 8832
rect 17092 8820 17098 8832
rect 17494 8820 17500 8832
rect 17092 8792 17500 8820
rect 17092 8780 17098 8792
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 17678 8780 17684 8832
rect 17736 8820 17742 8832
rect 17865 8823 17923 8829
rect 17865 8820 17877 8823
rect 17736 8792 17877 8820
rect 17736 8780 17742 8792
rect 17865 8789 17877 8792
rect 17911 8789 17923 8823
rect 18414 8820 18420 8832
rect 18375 8792 18420 8820
rect 17865 8783 17923 8789
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 1104 8730 18860 8752
rect 1104 8678 5398 8730
rect 5450 8678 5462 8730
rect 5514 8678 5526 8730
rect 5578 8678 5590 8730
rect 5642 8678 5654 8730
rect 5706 8678 9846 8730
rect 9898 8678 9910 8730
rect 9962 8678 9974 8730
rect 10026 8678 10038 8730
rect 10090 8678 10102 8730
rect 10154 8678 14294 8730
rect 14346 8678 14358 8730
rect 14410 8678 14422 8730
rect 14474 8678 14486 8730
rect 14538 8678 14550 8730
rect 14602 8678 18860 8730
rect 1104 8656 18860 8678
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 3142 8616 3148 8628
rect 2188 8588 3148 8616
rect 2188 8576 2194 8588
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 3237 8619 3295 8625
rect 3237 8585 3249 8619
rect 3283 8616 3295 8619
rect 3786 8616 3792 8628
rect 3283 8588 3792 8616
rect 3283 8585 3295 8588
rect 3237 8579 3295 8585
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 3878 8576 3884 8628
rect 3936 8576 3942 8628
rect 4430 8616 4436 8628
rect 4391 8588 4436 8616
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 6365 8619 6423 8625
rect 6365 8616 6377 8619
rect 5316 8588 6377 8616
rect 5316 8576 5322 8588
rect 6365 8585 6377 8588
rect 6411 8585 6423 8619
rect 6365 8579 6423 8585
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 6788 8588 6837 8616
rect 6788 8576 6794 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 6825 8579 6883 8585
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 10502 8616 10508 8628
rect 8619 8588 10364 8616
rect 10463 8588 10508 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 1673 8551 1731 8557
rect 1673 8517 1685 8551
rect 1719 8548 1731 8551
rect 1946 8548 1952 8560
rect 1719 8520 1952 8548
rect 1719 8517 1731 8520
rect 1673 8511 1731 8517
rect 1946 8508 1952 8520
rect 2004 8508 2010 8560
rect 2501 8551 2559 8557
rect 2501 8517 2513 8551
rect 2547 8548 2559 8551
rect 3329 8551 3387 8557
rect 2547 8520 2636 8548
rect 2547 8517 2559 8520
rect 2501 8511 2559 8517
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2314 8480 2320 8492
rect 1903 8452 2320 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2608 8480 2636 8520
rect 3329 8517 3341 8551
rect 3375 8548 3387 8551
rect 3896 8548 3924 8576
rect 3375 8520 3924 8548
rect 3375 8517 3387 8520
rect 3329 8511 3387 8517
rect 4246 8508 4252 8560
rect 4304 8548 4310 8560
rect 4614 8548 4620 8560
rect 4304 8520 4620 8548
rect 4304 8508 4310 8520
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 5902 8548 5908 8560
rect 4816 8520 5908 8548
rect 2958 8480 2964 8492
rect 2608 8452 2964 8480
rect 2409 8443 2467 8449
rect 1118 8372 1124 8424
rect 1176 8412 1182 8424
rect 2424 8412 2452 8443
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 4816 8489 4844 8520
rect 5902 8508 5908 8520
rect 5960 8548 5966 8560
rect 6546 8548 6552 8560
rect 5960 8520 6552 8548
rect 5960 8508 5966 8520
rect 6546 8508 6552 8520
rect 6604 8548 6610 8560
rect 6604 8520 7236 8548
rect 6604 8508 6610 8520
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 2682 8412 2688 8424
rect 1176 8384 2452 8412
rect 2643 8384 2688 8412
rect 1176 8372 1182 8384
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 3418 8372 3424 8424
rect 3476 8412 3482 8424
rect 3881 8415 3939 8421
rect 3476 8384 3521 8412
rect 3476 8372 3482 8384
rect 3881 8381 3893 8415
rect 3927 8412 3939 8415
rect 4246 8412 4252 8424
rect 3927 8384 4252 8412
rect 3927 8381 3939 8384
rect 3881 8375 3939 8381
rect 4246 8372 4252 8384
rect 4304 8372 4310 8424
rect 4356 8356 4384 8443
rect 4890 8440 4896 8492
rect 4948 8440 4954 8492
rect 5068 8483 5126 8489
rect 5068 8449 5080 8483
rect 5114 8480 5126 8483
rect 5810 8480 5816 8492
rect 5114 8452 5816 8480
rect 5114 8449 5126 8452
rect 5068 8443 5126 8449
rect 5810 8440 5816 8452
rect 5868 8480 5874 8492
rect 6362 8480 6368 8492
rect 5868 8452 6368 8480
rect 5868 8440 5874 8452
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 7208 8489 7236 8520
rect 7282 8508 7288 8560
rect 7340 8548 7346 8560
rect 7438 8551 7496 8557
rect 7438 8548 7450 8551
rect 7340 8520 7450 8548
rect 7340 8508 7346 8520
rect 7438 8517 7450 8520
rect 7484 8517 7496 8551
rect 7438 8511 7496 8517
rect 8386 8508 8392 8560
rect 8444 8548 8450 8560
rect 8849 8551 8907 8557
rect 8849 8548 8861 8551
rect 8444 8520 8861 8548
rect 8444 8508 8450 8520
rect 8849 8517 8861 8520
rect 8895 8548 8907 8551
rect 8938 8548 8944 8560
rect 8895 8520 8944 8548
rect 8895 8517 8907 8520
rect 8849 8511 8907 8517
rect 8938 8508 8944 8520
rect 8996 8508 9002 8560
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 9370 8551 9428 8557
rect 9370 8548 9382 8551
rect 9272 8520 9382 8548
rect 9272 8508 9278 8520
rect 9370 8517 9382 8520
rect 9416 8517 9428 8551
rect 9370 8511 9428 8517
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 7193 8483 7251 8489
rect 6779 8452 7144 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 4617 8415 4675 8421
rect 4617 8381 4629 8415
rect 4663 8412 4675 8415
rect 4908 8412 4936 8440
rect 4663 8384 4936 8412
rect 4663 8381 4675 8384
rect 4617 8375 4675 8381
rect 6454 8372 6460 8424
rect 6512 8412 6518 8424
rect 6917 8415 6975 8421
rect 6512 8384 6776 8412
rect 6512 8372 6518 8384
rect 6748 8356 6776 8384
rect 6917 8381 6929 8415
rect 6963 8381 6975 8415
rect 6917 8375 6975 8381
rect 7116 8412 7144 8452
rect 7193 8449 7205 8483
rect 7239 8449 7251 8483
rect 8202 8480 8208 8492
rect 7193 8443 7251 8449
rect 7300 8452 8208 8480
rect 7300 8412 7328 8452
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 10336 8480 10364 8588
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 11609 8619 11667 8625
rect 11609 8585 11621 8619
rect 11655 8616 11667 8619
rect 11790 8616 11796 8628
rect 11655 8588 11796 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 14829 8619 14887 8625
rect 14829 8616 14841 8619
rect 14700 8588 14841 8616
rect 14700 8576 14706 8588
rect 14829 8585 14841 8588
rect 14875 8585 14887 8619
rect 14829 8579 14887 8585
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 16669 8619 16727 8625
rect 16669 8616 16681 8619
rect 16632 8588 16681 8616
rect 16632 8576 16638 8588
rect 16669 8585 16681 8588
rect 16715 8585 16727 8619
rect 16669 8579 16727 8585
rect 16942 8576 16948 8628
rect 17000 8616 17006 8628
rect 17000 8588 17908 8616
rect 17000 8576 17006 8588
rect 12744 8551 12802 8557
rect 12744 8517 12756 8551
rect 12790 8548 12802 8551
rect 13906 8548 13912 8560
rect 12790 8520 13912 8548
rect 12790 8517 12802 8520
rect 12744 8511 12802 8517
rect 13906 8508 13912 8520
rect 13964 8508 13970 8560
rect 15562 8548 15568 8560
rect 14016 8520 15568 8548
rect 11054 8480 11060 8492
rect 10336 8452 11060 8480
rect 11054 8440 11060 8452
rect 11112 8480 11118 8492
rect 11330 8480 11336 8492
rect 11112 8452 11336 8480
rect 11112 8440 11118 8452
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 13716 8483 13774 8489
rect 13716 8449 13728 8483
rect 13762 8480 13774 8483
rect 14016 8480 14044 8520
rect 15562 8508 15568 8520
rect 15620 8508 15626 8560
rect 15654 8508 15660 8560
rect 15712 8548 15718 8560
rect 15712 8520 17172 8548
rect 15712 8508 15718 8520
rect 13762 8452 14044 8480
rect 13762 8449 13774 8452
rect 13716 8443 13774 8449
rect 14090 8440 14096 8492
rect 14148 8480 14154 8492
rect 16034 8483 16092 8489
rect 16034 8480 16046 8483
rect 14148 8452 16046 8480
rect 14148 8440 14154 8452
rect 16034 8449 16046 8452
rect 16080 8480 16092 8483
rect 16206 8480 16212 8492
rect 16080 8452 16212 8480
rect 16080 8449 16092 8452
rect 16034 8443 16092 8449
rect 16206 8440 16212 8452
rect 16264 8440 16270 8492
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 17034 8480 17040 8492
rect 16816 8452 17040 8480
rect 16816 8440 16822 8452
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 17144 8480 17172 8520
rect 17586 8508 17592 8560
rect 17644 8548 17650 8560
rect 17681 8551 17739 8557
rect 17681 8548 17693 8551
rect 17644 8520 17693 8548
rect 17644 8508 17650 8520
rect 17681 8517 17693 8520
rect 17727 8548 17739 8551
rect 17770 8548 17776 8560
rect 17727 8520 17776 8548
rect 17727 8517 17739 8520
rect 17681 8511 17739 8517
rect 17770 8508 17776 8520
rect 17828 8508 17834 8560
rect 17880 8489 17908 8588
rect 17865 8483 17923 8489
rect 17144 8452 17264 8480
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 7116 8384 7328 8412
rect 8956 8384 9137 8412
rect 2222 8344 2228 8356
rect 1872 8316 2228 8344
rect 1872 8288 1900 8316
rect 2222 8304 2228 8316
rect 2280 8304 2286 8356
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8344 2927 8347
rect 3510 8344 3516 8356
rect 2915 8316 3516 8344
rect 2915 8313 2927 8316
rect 2869 8307 2927 8313
rect 3510 8304 3516 8316
rect 3568 8304 3574 8356
rect 3970 8344 3976 8356
rect 3931 8316 3976 8344
rect 3970 8304 3976 8316
rect 4028 8304 4034 8356
rect 4338 8304 4344 8356
rect 4396 8304 4402 8356
rect 4430 8304 4436 8356
rect 4488 8344 4494 8356
rect 6181 8347 6239 8353
rect 4488 8316 4844 8344
rect 4488 8304 4494 8316
rect 1854 8236 1860 8288
rect 1912 8236 1918 8288
rect 4816 8276 4844 8316
rect 6181 8313 6193 8347
rect 6227 8344 6239 8347
rect 6638 8344 6644 8356
rect 6227 8316 6644 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 6730 8304 6736 8356
rect 6788 8344 6794 8356
rect 6932 8344 6960 8375
rect 6788 8316 6960 8344
rect 6788 8304 6794 8316
rect 6546 8276 6552 8288
rect 4816 8248 6552 8276
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 6822 8236 6828 8288
rect 6880 8276 6886 8288
rect 7116 8276 7144 8384
rect 6880 8248 7144 8276
rect 6880 8236 6886 8248
rect 8846 8236 8852 8288
rect 8904 8276 8910 8288
rect 8956 8285 8984 8384
rect 9125 8381 9137 8384
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 12989 8415 13047 8421
rect 12989 8381 13001 8415
rect 13035 8412 13047 8415
rect 13357 8415 13415 8421
rect 13357 8412 13369 8415
rect 13035 8384 13369 8412
rect 13035 8381 13047 8384
rect 12989 8375 13047 8381
rect 13357 8381 13369 8384
rect 13403 8412 13415 8415
rect 13446 8412 13452 8424
rect 13403 8384 13452 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 16301 8415 16359 8421
rect 16301 8381 16313 8415
rect 16347 8412 16359 8415
rect 16390 8412 16396 8424
rect 16347 8384 16396 8412
rect 16347 8381 16359 8384
rect 16301 8375 16359 8381
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 16482 8372 16488 8424
rect 16540 8412 16546 8424
rect 17236 8421 17264 8452
rect 17865 8449 17877 8483
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 18138 8440 18144 8492
rect 18196 8480 18202 8492
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 18196 8452 18245 8480
rect 18196 8440 18202 8452
rect 18233 8449 18245 8452
rect 18279 8449 18291 8483
rect 18233 8443 18291 8449
rect 17129 8415 17187 8421
rect 17129 8412 17141 8415
rect 16540 8384 17141 8412
rect 16540 8372 16546 8384
rect 17129 8381 17141 8384
rect 17175 8381 17187 8415
rect 17129 8375 17187 8381
rect 17221 8415 17279 8421
rect 17221 8381 17233 8415
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 14918 8344 14924 8356
rect 14879 8316 14924 8344
rect 14918 8304 14924 8316
rect 14976 8304 14982 8356
rect 16942 8344 16948 8356
rect 16316 8316 16948 8344
rect 8941 8279 8999 8285
rect 8941 8276 8953 8279
rect 8904 8248 8953 8276
rect 8904 8236 8910 8248
rect 8941 8245 8953 8248
rect 8987 8245 8999 8279
rect 8941 8239 8999 8245
rect 10689 8279 10747 8285
rect 10689 8245 10701 8279
rect 10735 8276 10747 8279
rect 10962 8276 10968 8288
rect 10735 8248 10968 8276
rect 10735 8245 10747 8248
rect 10689 8239 10747 8245
rect 10962 8236 10968 8248
rect 11020 8276 11026 8288
rect 11241 8279 11299 8285
rect 11241 8276 11253 8279
rect 11020 8248 11253 8276
rect 11020 8236 11026 8248
rect 11241 8245 11253 8248
rect 11287 8245 11299 8279
rect 11241 8239 11299 8245
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 16316 8276 16344 8316
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 17497 8347 17555 8353
rect 17497 8344 17509 8347
rect 17144 8316 17509 8344
rect 17144 8288 17172 8316
rect 17497 8313 17509 8316
rect 17543 8344 17555 8347
rect 17862 8344 17868 8356
rect 17543 8316 17868 8344
rect 17543 8313 17555 8316
rect 17497 8307 17555 8313
rect 17862 8304 17868 8316
rect 17920 8304 17926 8356
rect 18046 8344 18052 8356
rect 18007 8316 18052 8344
rect 18046 8304 18052 8316
rect 18104 8304 18110 8356
rect 18417 8347 18475 8353
rect 18417 8313 18429 8347
rect 18463 8344 18475 8347
rect 18506 8344 18512 8356
rect 18463 8316 18512 8344
rect 18463 8313 18475 8316
rect 18417 8307 18475 8313
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 15344 8248 16344 8276
rect 15344 8236 15350 8248
rect 17126 8236 17132 8288
rect 17184 8236 17190 8288
rect 1104 8186 18860 8208
rect 1104 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 3430 8186
rect 3482 8134 7622 8186
rect 7674 8134 7686 8186
rect 7738 8134 7750 8186
rect 7802 8134 7814 8186
rect 7866 8134 7878 8186
rect 7930 8134 12070 8186
rect 12122 8134 12134 8186
rect 12186 8134 12198 8186
rect 12250 8134 12262 8186
rect 12314 8134 12326 8186
rect 12378 8134 16518 8186
rect 16570 8134 16582 8186
rect 16634 8134 16646 8186
rect 16698 8134 16710 8186
rect 16762 8134 16774 8186
rect 16826 8134 18860 8186
rect 1104 8112 18860 8134
rect 2222 8072 2228 8084
rect 2183 8044 2228 8072
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2593 8075 2651 8081
rect 2593 8041 2605 8075
rect 2639 8072 2651 8075
rect 3418 8072 3424 8084
rect 2639 8044 3424 8072
rect 2639 8041 2651 8044
rect 2593 8035 2651 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 4338 8032 4344 8084
rect 4396 8072 4402 8084
rect 4709 8075 4767 8081
rect 4709 8072 4721 8075
rect 4396 8044 4721 8072
rect 4396 8032 4402 8044
rect 4709 8041 4721 8044
rect 4755 8041 4767 8075
rect 4709 8035 4767 8041
rect 5537 8075 5595 8081
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 5718 8072 5724 8084
rect 5583 8044 5724 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 7282 8072 7288 8084
rect 7243 8044 7288 8072
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 7392 8044 9597 8072
rect 2682 8004 2688 8016
rect 2643 7976 2688 8004
rect 2682 7964 2688 7976
rect 2740 8004 2746 8016
rect 3326 8004 3332 8016
rect 2740 7976 3332 8004
rect 2740 7964 2746 7976
rect 3326 7964 3332 7976
rect 3384 7964 3390 8016
rect 5626 8004 5632 8016
rect 3528 7976 4936 8004
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 1719 7908 2268 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 2240 7880 2268 7908
rect 3142 7896 3148 7948
rect 3200 7936 3206 7948
rect 3528 7945 3556 7976
rect 3513 7939 3571 7945
rect 3513 7936 3525 7939
rect 3200 7908 3525 7936
rect 3200 7896 3206 7908
rect 3513 7905 3525 7908
rect 3559 7905 3571 7939
rect 4154 7936 4160 7948
rect 4067 7908 4160 7936
rect 3513 7899 3571 7905
rect 4154 7896 4160 7908
rect 4212 7936 4218 7948
rect 4522 7936 4528 7948
rect 4212 7908 4528 7936
rect 4212 7896 4218 7908
rect 4522 7896 4528 7908
rect 4580 7896 4586 7948
rect 1489 7871 1547 7877
rect 1489 7837 1501 7871
rect 1535 7868 1547 7871
rect 2041 7871 2099 7877
rect 2041 7868 2053 7871
rect 1535 7840 2053 7868
rect 1535 7837 1547 7840
rect 1489 7831 1547 7837
rect 2041 7837 2053 7840
rect 2087 7868 2099 7871
rect 2130 7868 2136 7880
rect 2087 7840 2136 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 2409 7871 2467 7877
rect 2409 7868 2421 7871
rect 2280 7840 2421 7868
rect 2280 7828 2286 7840
rect 2409 7837 2421 7840
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 3384 7840 4200 7868
rect 3384 7828 3390 7840
rect 3418 7800 3424 7812
rect 3252 7772 3424 7800
rect 1578 7692 1584 7744
rect 1636 7732 1642 7744
rect 1857 7735 1915 7741
rect 1857 7732 1869 7735
rect 1636 7704 1869 7732
rect 1636 7692 1642 7704
rect 1857 7701 1869 7704
rect 1903 7701 1915 7735
rect 1857 7695 1915 7701
rect 2682 7692 2688 7744
rect 2740 7732 2746 7744
rect 3252 7741 3280 7772
rect 3418 7760 3424 7772
rect 3476 7760 3482 7812
rect 4172 7800 4200 7840
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4341 7871 4399 7877
rect 4341 7868 4353 7871
rect 4304 7840 4353 7868
rect 4304 7828 4310 7840
rect 4341 7837 4353 7840
rect 4387 7837 4399 7871
rect 4908 7868 4936 7976
rect 5000 7976 5632 8004
rect 5000 7945 5028 7976
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 7190 7964 7196 8016
rect 7248 8004 7254 8016
rect 7392 8004 7420 8044
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 9585 8035 9643 8041
rect 12713 8075 12771 8081
rect 12713 8041 12725 8075
rect 12759 8072 12771 8075
rect 14090 8072 14096 8084
rect 12759 8044 14096 8072
rect 12759 8041 12771 8044
rect 12713 8035 12771 8041
rect 14090 8032 14096 8044
rect 14148 8032 14154 8084
rect 15565 8075 15623 8081
rect 15565 8072 15577 8075
rect 14200 8044 15577 8072
rect 7248 7976 7420 8004
rect 7248 7964 7254 7976
rect 13906 7964 13912 8016
rect 13964 8004 13970 8016
rect 14200 8004 14228 8044
rect 15565 8041 15577 8044
rect 15611 8041 15623 8075
rect 15565 8035 15623 8041
rect 15746 8032 15752 8084
rect 15804 8072 15810 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 15804 8044 17049 8072
rect 15804 8032 15810 8044
rect 17037 8041 17049 8044
rect 17083 8041 17095 8075
rect 17037 8035 17095 8041
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 18233 8075 18291 8081
rect 18233 8072 18245 8075
rect 17552 8044 18245 8072
rect 17552 8032 17558 8044
rect 18233 8041 18245 8044
rect 18279 8072 18291 8075
rect 18322 8072 18328 8084
rect 18279 8044 18328 8072
rect 18279 8041 18291 8044
rect 18233 8035 18291 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 13964 7976 14228 8004
rect 13964 7964 13970 7976
rect 16942 7964 16948 8016
rect 17000 8004 17006 8016
rect 17126 8004 17132 8016
rect 17000 7976 17132 8004
rect 17000 7964 17006 7976
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 18046 8004 18052 8016
rect 18007 7976 18052 8004
rect 18046 7964 18052 7976
rect 18104 7964 18110 8016
rect 4985 7939 5043 7945
rect 4985 7905 4997 7939
rect 5031 7905 5043 7939
rect 4985 7899 5043 7905
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7936 5135 7939
rect 5166 7936 5172 7948
rect 5123 7908 5172 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 9306 7936 9312 7948
rect 5276 7908 6040 7936
rect 5276 7868 5304 7908
rect 4908 7840 5304 7868
rect 5905 7871 5963 7877
rect 4341 7831 4399 7837
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 5074 7800 5080 7812
rect 4172 7772 5080 7800
rect 5074 7760 5080 7772
rect 5132 7760 5138 7812
rect 5169 7803 5227 7809
rect 5169 7769 5181 7803
rect 5215 7800 5227 7803
rect 5258 7800 5264 7812
rect 5215 7772 5264 7800
rect 5215 7769 5227 7772
rect 5169 7763 5227 7769
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 5920 7744 5948 7831
rect 6012 7800 6040 7908
rect 8680 7908 9312 7936
rect 6172 7871 6230 7877
rect 6172 7837 6184 7871
rect 6218 7868 6230 7871
rect 7466 7868 7472 7880
rect 6218 7840 7472 7868
rect 6218 7837 6230 7840
rect 6172 7831 6230 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 8680 7868 8708 7908
rect 9306 7896 9312 7908
rect 9364 7896 9370 7948
rect 17310 7896 17316 7948
rect 17368 7936 17374 7948
rect 17589 7939 17647 7945
rect 17589 7936 17601 7939
rect 17368 7908 17601 7936
rect 17368 7896 17374 7908
rect 17589 7905 17601 7908
rect 17635 7905 17647 7939
rect 17589 7899 17647 7905
rect 7576 7840 8708 7868
rect 8757 7871 8815 7877
rect 7576 7800 7604 7840
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 8846 7868 8852 7880
rect 8803 7840 8852 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 8846 7828 8852 7840
rect 8904 7868 8910 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8904 7840 8953 7868
rect 8904 7828 8910 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9490 7868 9496 7880
rect 9088 7840 9496 7868
rect 9088 7828 9094 7840
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 10226 7828 10232 7880
rect 10284 7868 10290 7880
rect 10698 7871 10756 7877
rect 10698 7868 10710 7871
rect 10284 7840 10710 7868
rect 10284 7828 10290 7840
rect 10698 7837 10710 7840
rect 10744 7868 10756 7871
rect 10744 7840 10916 7868
rect 10744 7837 10756 7840
rect 10698 7831 10756 7837
rect 6012 7772 7604 7800
rect 8512 7803 8570 7809
rect 8512 7769 8524 7803
rect 8558 7800 8570 7803
rect 9766 7800 9772 7812
rect 8558 7772 9772 7800
rect 8558 7769 8570 7772
rect 8512 7763 8570 7769
rect 9766 7760 9772 7772
rect 9824 7800 9830 7812
rect 10778 7800 10784 7812
rect 9824 7772 10784 7800
rect 9824 7760 9830 7772
rect 10778 7760 10784 7772
rect 10836 7760 10842 7812
rect 10888 7800 10916 7840
rect 10962 7828 10968 7880
rect 11020 7868 11026 7880
rect 11149 7871 11207 7877
rect 11149 7868 11161 7871
rect 11020 7840 11161 7868
rect 11020 7828 11026 7840
rect 11149 7837 11161 7840
rect 11195 7868 11207 7871
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 11195 7840 11345 7868
rect 11195 7837 11207 7840
rect 11149 7831 11207 7837
rect 11333 7837 11345 7840
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11422 7828 11428 7880
rect 11480 7868 11486 7880
rect 11589 7871 11647 7877
rect 11589 7868 11601 7871
rect 11480 7840 11601 7868
rect 11480 7828 11486 7840
rect 11589 7837 11601 7840
rect 11635 7837 11647 7871
rect 11589 7831 11647 7837
rect 13446 7828 13452 7880
rect 13504 7868 13510 7880
rect 13817 7871 13875 7877
rect 13817 7868 13829 7871
rect 13504 7840 13829 7868
rect 13504 7828 13510 7840
rect 13817 7837 13829 7840
rect 13863 7868 13875 7871
rect 15470 7868 15476 7880
rect 13863 7840 15476 7868
rect 13863 7837 13875 7840
rect 13817 7831 13875 7837
rect 15470 7828 15476 7840
rect 15528 7868 15534 7880
rect 16390 7868 16396 7880
rect 15528 7840 16396 7868
rect 15528 7828 15534 7840
rect 16390 7828 16396 7840
rect 16448 7868 16454 7880
rect 16945 7871 17003 7877
rect 16945 7868 16957 7871
rect 16448 7840 16957 7868
rect 16448 7828 16454 7840
rect 16945 7837 16957 7840
rect 16991 7837 17003 7871
rect 16945 7831 17003 7837
rect 17218 7828 17224 7880
rect 17276 7868 17282 7880
rect 17405 7871 17463 7877
rect 17405 7868 17417 7871
rect 17276 7840 17417 7868
rect 17276 7828 17282 7840
rect 17405 7837 17417 7840
rect 17451 7837 17463 7871
rect 17862 7868 17868 7880
rect 17823 7840 17868 7868
rect 17405 7831 17463 7837
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 11238 7800 11244 7812
rect 10888 7772 11244 7800
rect 11238 7760 11244 7772
rect 11296 7760 11302 7812
rect 15206 7803 15264 7809
rect 15206 7800 15218 7803
rect 12406 7772 15218 7800
rect 2869 7735 2927 7741
rect 2869 7732 2881 7735
rect 2740 7704 2881 7732
rect 2740 7692 2746 7704
rect 2869 7701 2881 7704
rect 2915 7701 2927 7735
rect 2869 7695 2927 7701
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7701 3295 7735
rect 3237 7695 3295 7701
rect 3326 7692 3332 7744
rect 3384 7732 3390 7744
rect 3789 7735 3847 7741
rect 3789 7732 3801 7735
rect 3384 7704 3801 7732
rect 3384 7692 3390 7704
rect 3789 7701 3801 7704
rect 3835 7701 3847 7735
rect 4246 7732 4252 7744
rect 4207 7704 4252 7732
rect 3789 7695 3847 7701
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7732 5871 7735
rect 5902 7732 5908 7744
rect 5859 7704 5908 7732
rect 5859 7701 5871 7704
rect 5813 7695 5871 7701
rect 5902 7692 5908 7704
rect 5960 7692 5966 7744
rect 7282 7692 7288 7744
rect 7340 7732 7346 7744
rect 7377 7735 7435 7741
rect 7377 7732 7389 7735
rect 7340 7704 7389 7732
rect 7340 7692 7346 7704
rect 7377 7701 7389 7704
rect 7423 7732 7435 7735
rect 9122 7732 9128 7744
rect 7423 7704 9128 7732
rect 7423 7701 7435 7704
rect 7377 7695 7435 7701
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 10502 7692 10508 7744
rect 10560 7732 10566 7744
rect 12406 7732 12434 7772
rect 15206 7769 15218 7772
rect 15252 7769 15264 7803
rect 15206 7763 15264 7769
rect 16700 7803 16758 7809
rect 16700 7769 16712 7803
rect 16746 7800 16758 7803
rect 17034 7800 17040 7812
rect 16746 7772 17040 7800
rect 16746 7769 16758 7772
rect 16700 7763 16758 7769
rect 17034 7760 17040 7772
rect 17092 7760 17098 7812
rect 17126 7760 17132 7812
rect 17184 7800 17190 7812
rect 17497 7803 17555 7809
rect 17497 7800 17509 7803
rect 17184 7772 17509 7800
rect 17184 7760 17190 7772
rect 17497 7769 17509 7772
rect 17543 7769 17555 7803
rect 17497 7763 17555 7769
rect 17678 7760 17684 7812
rect 17736 7800 17742 7812
rect 18417 7803 18475 7809
rect 18417 7800 18429 7803
rect 17736 7772 18429 7800
rect 17736 7760 17742 7772
rect 18417 7769 18429 7772
rect 18463 7769 18475 7803
rect 18417 7763 18475 7769
rect 10560 7704 12434 7732
rect 10560 7692 10566 7704
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 13633 7735 13691 7741
rect 13633 7732 13645 7735
rect 13596 7704 13645 7732
rect 13596 7692 13602 7704
rect 13633 7701 13645 7704
rect 13679 7701 13691 7735
rect 13633 7695 13691 7701
rect 13906 7692 13912 7744
rect 13964 7732 13970 7744
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 13964 7704 14105 7732
rect 13964 7692 13970 7704
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 14093 7695 14151 7701
rect 1104 7642 18860 7664
rect 1104 7590 5398 7642
rect 5450 7590 5462 7642
rect 5514 7590 5526 7642
rect 5578 7590 5590 7642
rect 5642 7590 5654 7642
rect 5706 7590 9846 7642
rect 9898 7590 9910 7642
rect 9962 7590 9974 7642
rect 10026 7590 10038 7642
rect 10090 7590 10102 7642
rect 10154 7590 14294 7642
rect 14346 7590 14358 7642
rect 14410 7590 14422 7642
rect 14474 7590 14486 7642
rect 14538 7590 14550 7642
rect 14602 7590 18860 7642
rect 1104 7568 18860 7590
rect 2961 7531 3019 7537
rect 2961 7497 2973 7531
rect 3007 7528 3019 7531
rect 3050 7528 3056 7540
rect 3007 7500 3056 7528
rect 3007 7497 3019 7500
rect 2961 7491 3019 7497
rect 3050 7488 3056 7500
rect 3108 7528 3114 7540
rect 3329 7531 3387 7537
rect 3108 7500 3280 7528
rect 3108 7488 3114 7500
rect 3252 7460 3280 7500
rect 3329 7497 3341 7531
rect 3375 7528 3387 7531
rect 3418 7528 3424 7540
rect 3375 7500 3424 7528
rect 3375 7497 3387 7500
rect 3329 7491 3387 7497
rect 3418 7488 3424 7500
rect 3476 7488 3482 7540
rect 3878 7528 3884 7540
rect 3839 7500 3884 7528
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 4617 7531 4675 7537
rect 4617 7497 4629 7531
rect 4663 7528 4675 7531
rect 4798 7528 4804 7540
rect 4663 7500 4804 7528
rect 4663 7497 4675 7500
rect 4617 7491 4675 7497
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 5077 7531 5135 7537
rect 5077 7497 5089 7531
rect 5123 7528 5135 7531
rect 5166 7528 5172 7540
rect 5123 7500 5172 7528
rect 5123 7497 5135 7500
rect 5077 7491 5135 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 6457 7531 6515 7537
rect 5316 7500 6132 7528
rect 5316 7488 5322 7500
rect 3602 7460 3608 7472
rect 3252 7432 3608 7460
rect 3602 7420 3608 7432
rect 3660 7420 3666 7472
rect 4522 7460 4528 7472
rect 4483 7432 4528 7460
rect 4522 7420 4528 7432
rect 4580 7420 4586 7472
rect 4985 7463 5043 7469
rect 4985 7429 4997 7463
rect 5031 7460 5043 7463
rect 5994 7460 6000 7472
rect 5031 7432 6000 7460
rect 5031 7429 5043 7432
rect 4985 7423 5043 7429
rect 5994 7420 6000 7432
rect 6052 7420 6058 7472
rect 6104 7460 6132 7500
rect 6457 7497 6469 7531
rect 6503 7528 6515 7531
rect 6822 7528 6828 7540
rect 6503 7500 6828 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7466 7488 7472 7540
rect 7524 7528 7530 7540
rect 7650 7528 7656 7540
rect 7524 7500 7656 7528
rect 7524 7488 7530 7500
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 8294 7528 8300 7540
rect 7975 7500 8300 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8294 7488 8300 7500
rect 8352 7528 8358 7540
rect 8570 7528 8576 7540
rect 8352 7500 8576 7528
rect 8352 7488 8358 7500
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 12894 7528 12900 7540
rect 12855 7500 12900 7528
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 13354 7528 13360 7540
rect 13315 7500 13360 7528
rect 13354 7488 13360 7500
rect 13412 7488 13418 7540
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 13541 7531 13599 7537
rect 13541 7528 13553 7531
rect 13504 7500 13553 7528
rect 13504 7488 13510 7500
rect 13541 7497 13553 7500
rect 13587 7497 13599 7531
rect 13541 7491 13599 7497
rect 13725 7531 13783 7537
rect 13725 7497 13737 7531
rect 13771 7528 13783 7531
rect 13814 7528 13820 7540
rect 13771 7500 13820 7528
rect 13771 7497 13783 7500
rect 13725 7491 13783 7497
rect 13814 7488 13820 7500
rect 13872 7528 13878 7540
rect 14182 7528 14188 7540
rect 13872 7500 14188 7528
rect 13872 7488 13878 7500
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 15286 7528 15292 7540
rect 15247 7500 15292 7528
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 15470 7528 15476 7540
rect 15431 7500 15476 7528
rect 15470 7488 15476 7500
rect 15528 7528 15534 7540
rect 15565 7531 15623 7537
rect 15565 7528 15577 7531
rect 15528 7500 15577 7528
rect 15528 7488 15534 7500
rect 15565 7497 15577 7500
rect 15611 7497 15623 7531
rect 15565 7491 15623 7497
rect 16209 7531 16267 7537
rect 16209 7497 16221 7531
rect 16255 7528 16267 7531
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 16255 7500 16681 7528
rect 16255 7497 16267 7500
rect 16209 7491 16267 7497
rect 16669 7497 16681 7500
rect 16715 7497 16727 7531
rect 16669 7491 16727 7497
rect 17129 7531 17187 7537
rect 17129 7497 17141 7531
rect 17175 7528 17187 7531
rect 17862 7528 17868 7540
rect 17175 7500 17724 7528
rect 17823 7500 17868 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 6104 7432 7604 7460
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 2130 7392 2136 7404
rect 2091 7364 2136 7392
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 3142 7392 3148 7404
rect 2792 7364 3148 7392
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7293 2007 7327
rect 1949 7287 2007 7293
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7324 2099 7327
rect 2314 7324 2320 7336
rect 2087 7296 2320 7324
rect 2087 7293 2099 7296
rect 2041 7287 2099 7293
rect 1486 7256 1492 7268
rect 1447 7228 1492 7256
rect 1486 7216 1492 7228
rect 1544 7216 1550 7268
rect 1964 7256 1992 7287
rect 2314 7284 2320 7296
rect 2372 7284 2378 7336
rect 2792 7333 2820 7364
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7392 3847 7395
rect 3835 7364 4200 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 2777 7327 2835 7333
rect 2777 7293 2789 7327
rect 2823 7293 2835 7327
rect 2777 7287 2835 7293
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7293 2927 7327
rect 2869 7287 2927 7293
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7293 4031 7327
rect 3973 7287 4031 7293
rect 2792 7256 2820 7287
rect 1964 7228 2820 7256
rect 2498 7188 2504 7200
rect 2459 7160 2504 7188
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 2884 7188 2912 7287
rect 2958 7216 2964 7268
rect 3016 7256 3022 7268
rect 3016 7228 3464 7256
rect 3016 7216 3022 7228
rect 3050 7188 3056 7200
rect 2884 7160 3056 7188
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 3436 7197 3464 7228
rect 3786 7216 3792 7268
rect 3844 7256 3850 7268
rect 3988 7256 4016 7287
rect 4172 7256 4200 7364
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 5626 7392 5632 7404
rect 4304 7364 5632 7392
rect 4304 7352 4310 7364
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 6816 7395 6874 7401
rect 6816 7361 6828 7395
rect 6862 7392 6874 7395
rect 7282 7392 7288 7404
rect 6862 7364 7288 7392
rect 6862 7361 6874 7364
rect 6816 7355 6874 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 4338 7284 4344 7336
rect 4396 7324 4402 7336
rect 5261 7327 5319 7333
rect 5261 7324 5273 7327
rect 4396 7296 5273 7324
rect 4396 7284 4402 7296
rect 5261 7293 5273 7296
rect 5307 7293 5319 7327
rect 5261 7287 5319 7293
rect 4246 7256 4252 7268
rect 3844 7228 4016 7256
rect 4159 7228 4252 7256
rect 3844 7216 3850 7228
rect 4246 7216 4252 7228
rect 4304 7256 4310 7268
rect 5276 7256 5304 7287
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 6549 7327 6607 7333
rect 6549 7324 6561 7327
rect 5960 7296 6561 7324
rect 5960 7284 5966 7296
rect 6549 7293 6561 7296
rect 6595 7293 6607 7327
rect 7576 7324 7604 7432
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 9398 7469 9404 7472
rect 9392 7460 9404 7469
rect 8168 7432 9260 7460
rect 9359 7432 9404 7460
rect 8168 7420 8174 7432
rect 8846 7352 8852 7404
rect 8904 7392 8910 7404
rect 9232 7392 9260 7432
rect 9392 7423 9404 7432
rect 9398 7420 9404 7423
rect 9456 7420 9462 7472
rect 11606 7420 11612 7472
rect 11664 7460 11670 7472
rect 11762 7463 11820 7469
rect 11762 7460 11774 7463
rect 11664 7432 11774 7460
rect 11664 7420 11670 7432
rect 11762 7429 11774 7432
rect 11808 7429 11820 7463
rect 11762 7423 11820 7429
rect 8904 7364 9168 7392
rect 9232 7364 10548 7392
rect 8904 7352 8910 7364
rect 9140 7336 9168 7364
rect 8938 7324 8944 7336
rect 7576 7296 8944 7324
rect 6549 7287 6607 7293
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 9122 7324 9128 7336
rect 9083 7296 9128 7324
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 8021 7259 8079 7265
rect 4304 7228 4384 7256
rect 5276 7228 6040 7256
rect 4304 7216 4310 7228
rect 4356 7197 4384 7228
rect 3421 7191 3479 7197
rect 3421 7157 3433 7191
rect 3467 7157 3479 7191
rect 3421 7151 3479 7157
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 5258 7188 5264 7200
rect 4387 7160 5264 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 5534 7188 5540 7200
rect 5495 7160 5540 7188
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 5902 7188 5908 7200
rect 5863 7160 5908 7188
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 6012 7188 6040 7228
rect 8021 7225 8033 7259
rect 8067 7256 8079 7259
rect 8205 7259 8263 7265
rect 8205 7256 8217 7259
rect 8067 7228 8217 7256
rect 8067 7225 8079 7228
rect 8021 7219 8079 7225
rect 8205 7225 8217 7228
rect 8251 7256 8263 7259
rect 9140 7256 9168 7284
rect 10520 7265 10548 7364
rect 10962 7352 10968 7404
rect 11020 7392 11026 7404
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 11020 7364 11529 7392
rect 11020 7352 11026 7364
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 14838 7395 14896 7401
rect 14838 7392 14850 7395
rect 13872 7364 14850 7392
rect 13872 7352 13878 7364
rect 14838 7361 14850 7364
rect 14884 7392 14896 7395
rect 15105 7395 15163 7401
rect 14884 7364 15056 7392
rect 14884 7361 14896 7364
rect 14838 7355 14896 7361
rect 11330 7324 11336 7336
rect 11291 7296 11336 7324
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 15028 7324 15056 7364
rect 15105 7361 15117 7395
rect 15151 7392 15163 7395
rect 15488 7392 15516 7488
rect 15746 7420 15752 7472
rect 15804 7460 15810 7472
rect 17144 7460 17172 7491
rect 15804 7432 17172 7460
rect 15804 7420 15810 7432
rect 17586 7420 17592 7472
rect 17644 7420 17650 7472
rect 16114 7392 16120 7404
rect 15151 7364 15516 7392
rect 16075 7364 16120 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 16850 7352 16856 7404
rect 16908 7392 16914 7404
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 16908 7364 17049 7392
rect 16908 7352 16914 7364
rect 17037 7361 17049 7364
rect 17083 7392 17095 7395
rect 17604 7392 17632 7420
rect 17083 7364 17632 7392
rect 17696 7392 17724 7500
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 17957 7395 18015 7401
rect 17957 7392 17969 7395
rect 17696 7364 17969 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17957 7361 17969 7364
rect 18003 7392 18015 7395
rect 19334 7392 19340 7404
rect 18003 7364 19340 7392
rect 18003 7361 18015 7364
rect 17957 7355 18015 7361
rect 19334 7352 19340 7364
rect 19392 7352 19398 7404
rect 15838 7324 15844 7336
rect 15028 7296 15844 7324
rect 15838 7284 15844 7296
rect 15896 7284 15902 7336
rect 16206 7284 16212 7336
rect 16264 7324 16270 7336
rect 16301 7327 16359 7333
rect 16301 7324 16313 7327
rect 16264 7296 16313 7324
rect 16264 7284 16270 7296
rect 16301 7293 16313 7296
rect 16347 7293 16359 7327
rect 16301 7287 16359 7293
rect 17313 7327 17371 7333
rect 17313 7293 17325 7327
rect 17359 7324 17371 7327
rect 17586 7324 17592 7336
rect 17359 7296 17592 7324
rect 17359 7293 17371 7296
rect 17313 7287 17371 7293
rect 17586 7284 17592 7296
rect 17644 7284 17650 7336
rect 17862 7284 17868 7336
rect 17920 7324 17926 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17920 7296 18061 7324
rect 17920 7284 17926 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18322 7324 18328 7336
rect 18283 7296 18328 7324
rect 18049 7287 18107 7293
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 8251 7228 9168 7256
rect 10505 7259 10563 7265
rect 8251 7225 8263 7228
rect 8205 7219 8263 7225
rect 10505 7225 10517 7259
rect 10551 7256 10563 7259
rect 10551 7228 11376 7256
rect 10551 7225 10563 7228
rect 10505 7219 10563 7225
rect 9490 7188 9496 7200
rect 6012 7160 9496 7188
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 10689 7191 10747 7197
rect 10689 7157 10701 7191
rect 10735 7188 10747 7191
rect 10962 7188 10968 7200
rect 10735 7160 10968 7188
rect 10735 7157 10747 7160
rect 10689 7151 10747 7157
rect 10962 7148 10968 7160
rect 11020 7188 11026 7200
rect 11057 7191 11115 7197
rect 11057 7188 11069 7191
rect 11020 7160 11069 7188
rect 11020 7148 11026 7160
rect 11057 7157 11069 7160
rect 11103 7157 11115 7191
rect 11348 7188 11376 7228
rect 12802 7188 12808 7200
rect 11348 7160 12808 7188
rect 11057 7151 11115 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 15746 7188 15752 7200
rect 15707 7160 15752 7188
rect 15746 7148 15752 7160
rect 15804 7148 15810 7200
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 17497 7191 17555 7197
rect 17497 7188 17509 7191
rect 16356 7160 17509 7188
rect 16356 7148 16362 7160
rect 17497 7157 17509 7160
rect 17543 7157 17555 7191
rect 17497 7151 17555 7157
rect 1104 7098 18860 7120
rect 1104 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 3430 7098
rect 3482 7046 7622 7098
rect 7674 7046 7686 7098
rect 7738 7046 7750 7098
rect 7802 7046 7814 7098
rect 7866 7046 7878 7098
rect 7930 7046 12070 7098
rect 12122 7046 12134 7098
rect 12186 7046 12198 7098
rect 12250 7046 12262 7098
rect 12314 7046 12326 7098
rect 12378 7046 16518 7098
rect 16570 7046 16582 7098
rect 16634 7046 16646 7098
rect 16698 7046 16710 7098
rect 16762 7046 16774 7098
rect 16826 7046 18860 7098
rect 1104 7024 18860 7046
rect 1670 6984 1676 6996
rect 1631 6956 1676 6984
rect 1670 6944 1676 6956
rect 1728 6944 1734 6996
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 2590 6984 2596 6996
rect 2372 6956 2596 6984
rect 2372 6944 2378 6956
rect 2590 6944 2596 6956
rect 2648 6944 2654 6996
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 3050 6984 3056 6996
rect 2924 6956 3056 6984
rect 2924 6944 2930 6956
rect 3050 6944 3056 6956
rect 3108 6944 3114 6996
rect 3878 6984 3884 6996
rect 3839 6956 3884 6984
rect 3878 6944 3884 6956
rect 3936 6944 3942 6996
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 7190 6984 7196 6996
rect 4120 6956 7196 6984
rect 4120 6944 4126 6956
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 7285 6987 7343 6993
rect 7285 6953 7297 6987
rect 7331 6984 7343 6987
rect 7466 6984 7472 6996
rect 7331 6956 7472 6984
rect 7331 6953 7343 6956
rect 7285 6947 7343 6953
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 9766 6944 9772 6996
rect 9824 6984 9830 6996
rect 9953 6987 10011 6993
rect 9953 6984 9965 6987
rect 9824 6956 9965 6984
rect 9824 6944 9830 6956
rect 9953 6953 9965 6956
rect 9999 6953 10011 6987
rect 11422 6984 11428 6996
rect 11383 6956 11428 6984
rect 9953 6947 10011 6953
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 13817 6987 13875 6993
rect 13817 6984 13829 6987
rect 13504 6956 13829 6984
rect 13504 6944 13510 6956
rect 13817 6953 13829 6956
rect 13863 6953 13875 6987
rect 18046 6984 18052 6996
rect 13817 6947 13875 6953
rect 14016 6956 17080 6984
rect 18007 6956 18052 6984
rect 2498 6876 2504 6928
rect 2556 6916 2562 6928
rect 4338 6916 4344 6928
rect 2556 6888 2774 6916
rect 2556 6876 2562 6888
rect 2130 6848 2136 6860
rect 2091 6820 2136 6848
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6780 1547 6783
rect 2041 6783 2099 6789
rect 2041 6780 2053 6783
rect 1535 6752 2053 6780
rect 1535 6749 1547 6752
rect 1489 6743 1547 6749
rect 2041 6749 2053 6752
rect 2087 6780 2099 6783
rect 2314 6780 2320 6792
rect 2087 6752 2320 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 2746 6780 2774 6888
rect 2976 6888 4344 6916
rect 2976 6857 3004 6888
rect 4338 6876 4344 6888
rect 4396 6876 4402 6928
rect 5626 6876 5632 6928
rect 5684 6916 5690 6928
rect 5813 6919 5871 6925
rect 5813 6916 5825 6919
rect 5684 6888 5825 6916
rect 5684 6876 5690 6888
rect 5813 6885 5825 6888
rect 5859 6885 5871 6919
rect 7374 6916 7380 6928
rect 7335 6888 7380 6916
rect 5813 6879 5871 6885
rect 7374 6876 7380 6888
rect 7432 6876 7438 6928
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6817 3019 6851
rect 2961 6811 3019 6817
rect 3050 6808 3056 6860
rect 3108 6848 3114 6860
rect 3145 6851 3203 6857
rect 3145 6848 3157 6851
rect 3108 6820 3157 6848
rect 3108 6808 3114 6820
rect 3145 6817 3157 6820
rect 3191 6817 3203 6851
rect 3145 6811 3203 6817
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 13081 6851 13139 6857
rect 13081 6848 13093 6851
rect 12952 6820 13093 6848
rect 12952 6808 12958 6820
rect 13081 6817 13093 6820
rect 13127 6817 13139 6851
rect 13081 6811 13139 6817
rect 13464 6848 13492 6944
rect 13538 6876 13544 6928
rect 13596 6916 13602 6928
rect 13725 6919 13783 6925
rect 13725 6916 13737 6919
rect 13596 6888 13737 6916
rect 13596 6876 13602 6888
rect 13725 6885 13737 6888
rect 13771 6916 13783 6919
rect 14016 6916 14044 6956
rect 17052 6928 17080 6956
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 13771 6888 14044 6916
rect 13771 6885 13783 6888
rect 13725 6879 13783 6885
rect 17034 6876 17040 6928
rect 17092 6916 17098 6928
rect 17218 6916 17224 6928
rect 17092 6888 17224 6916
rect 17092 6876 17098 6888
rect 17218 6876 17224 6888
rect 17276 6876 17282 6928
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 13464 6820 14105 6848
rect 3237 6783 3295 6789
rect 3237 6780 3249 6783
rect 2746 6752 3249 6780
rect 3237 6749 3249 6752
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 3602 6740 3608 6792
rect 3660 6740 3666 6792
rect 4062 6780 4068 6792
rect 4023 6752 4068 6780
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 4338 6780 4344 6792
rect 4295 6752 4344 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 4338 6740 4344 6752
rect 4396 6740 4402 6792
rect 4433 6783 4491 6789
rect 4433 6749 4445 6783
rect 4479 6780 4491 6783
rect 5902 6780 5908 6792
rect 4479 6752 5908 6780
rect 4479 6749 4491 6752
rect 4433 6743 4491 6749
rect 2501 6715 2559 6721
rect 2501 6681 2513 6715
rect 2547 6712 2559 6715
rect 3620 6712 3648 6740
rect 4816 6724 4844 6752
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 7098 6780 7104 6792
rect 6052 6752 7104 6780
rect 6052 6740 6058 6752
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 8757 6783 8815 6789
rect 8757 6749 8769 6783
rect 8803 6780 8815 6783
rect 8803 6752 9076 6780
rect 8803 6749 8815 6752
rect 8757 6743 8815 6749
rect 2547 6684 3648 6712
rect 4700 6715 4758 6721
rect 2547 6681 2559 6684
rect 2501 6675 2559 6681
rect 4700 6681 4712 6715
rect 4746 6681 4758 6715
rect 4700 6675 4758 6681
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 1857 6647 1915 6653
rect 1857 6644 1869 6647
rect 1544 6616 1869 6644
rect 1544 6604 1550 6616
rect 1857 6613 1869 6616
rect 1903 6613 1915 6647
rect 1857 6607 1915 6613
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 3050 6644 3056 6656
rect 2740 6616 3056 6644
rect 2740 6604 2746 6616
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3602 6644 3608 6656
rect 3563 6616 3608 6644
rect 3602 6604 3608 6616
rect 3660 6604 3666 6656
rect 4724 6644 4752 6675
rect 4798 6672 4804 6724
rect 4856 6672 4862 6724
rect 5074 6672 5080 6724
rect 5132 6712 5138 6724
rect 6172 6715 6230 6721
rect 5132 6684 6132 6712
rect 5132 6672 5138 6684
rect 5718 6644 5724 6656
rect 4724 6616 5724 6644
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 6104 6644 6132 6684
rect 6172 6681 6184 6715
rect 6218 6712 6230 6715
rect 7374 6712 7380 6724
rect 6218 6684 7380 6712
rect 6218 6681 6230 6684
rect 6172 6675 6230 6681
rect 7374 6672 7380 6684
rect 7432 6672 7438 6724
rect 8512 6715 8570 6721
rect 8512 6681 8524 6715
rect 8558 6712 8570 6715
rect 8662 6712 8668 6724
rect 8558 6684 8668 6712
rect 8558 6681 8570 6684
rect 8512 6675 8570 6681
rect 8662 6672 8668 6684
rect 8720 6672 8726 6724
rect 8846 6644 8852 6656
rect 6104 6616 8852 6644
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 9048 6653 9076 6752
rect 11054 6740 11060 6792
rect 11112 6789 11118 6792
rect 11112 6780 11124 6789
rect 11333 6783 11391 6789
rect 11112 6752 11157 6780
rect 11112 6743 11124 6752
rect 11333 6749 11345 6783
rect 11379 6749 11391 6783
rect 11333 6743 11391 6749
rect 11112 6740 11118 6743
rect 10962 6672 10968 6724
rect 11020 6712 11026 6724
rect 11348 6712 11376 6743
rect 12066 6740 12072 6792
rect 12124 6780 12130 6792
rect 12805 6783 12863 6789
rect 12124 6752 12756 6780
rect 12124 6740 12130 6752
rect 11020 6684 11376 6712
rect 11020 6672 11026 6684
rect 11698 6672 11704 6724
rect 11756 6712 11762 6724
rect 11974 6712 11980 6724
rect 11756 6684 11980 6712
rect 11756 6672 11762 6684
rect 11974 6672 11980 6684
rect 12032 6712 12038 6724
rect 12538 6715 12596 6721
rect 12538 6712 12550 6715
rect 12032 6684 12550 6712
rect 12032 6672 12038 6684
rect 12538 6681 12550 6684
rect 12584 6681 12596 6715
rect 12728 6712 12756 6752
rect 12805 6749 12817 6783
rect 12851 6780 12863 6783
rect 13464 6780 13492 6820
rect 14093 6817 14105 6820
rect 14139 6817 14151 6851
rect 17586 6848 17592 6860
rect 17547 6820 17592 6848
rect 14093 6811 14151 6817
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 18414 6808 18420 6860
rect 18472 6808 18478 6860
rect 12851 6752 13492 6780
rect 12851 6749 12863 6752
rect 12805 6743 12863 6749
rect 13630 6740 13636 6792
rect 13688 6780 13694 6792
rect 14349 6783 14407 6789
rect 14349 6780 14361 6783
rect 13688 6752 14361 6780
rect 13688 6740 13694 6752
rect 14349 6749 14361 6752
rect 14395 6749 14407 6783
rect 14349 6743 14407 6749
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 16945 6783 17003 6789
rect 16945 6780 16957 6783
rect 16448 6752 16957 6780
rect 16448 6740 16454 6752
rect 16945 6749 16957 6752
rect 16991 6749 17003 6783
rect 16945 6743 17003 6749
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17497 6783 17555 6789
rect 17497 6780 17509 6783
rect 17276 6752 17509 6780
rect 17276 6740 17282 6752
rect 17497 6749 17509 6752
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 17865 6783 17923 6789
rect 17865 6749 17877 6783
rect 17911 6749 17923 6783
rect 17865 6743 17923 6749
rect 18233 6783 18291 6789
rect 18233 6749 18245 6783
rect 18279 6780 18291 6783
rect 18432 6780 18460 6808
rect 19150 6780 19156 6792
rect 18279 6752 19156 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 13357 6715 13415 6721
rect 13357 6712 13369 6715
rect 12728 6684 13369 6712
rect 12538 6675 12596 6681
rect 13357 6681 13369 6684
rect 13403 6712 13415 6715
rect 13541 6715 13599 6721
rect 13541 6712 13553 6715
rect 13403 6684 13553 6712
rect 13403 6681 13415 6684
rect 13357 6675 13415 6681
rect 13541 6681 13553 6684
rect 13587 6712 13599 6715
rect 16574 6712 16580 6724
rect 13587 6684 16580 6712
rect 13587 6681 13599 6684
rect 13541 6675 13599 6681
rect 16574 6672 16580 6684
rect 16632 6672 16638 6724
rect 16700 6715 16758 6721
rect 16700 6681 16712 6715
rect 16746 6712 16758 6715
rect 16850 6712 16856 6724
rect 16746 6684 16856 6712
rect 16746 6681 16758 6684
rect 16700 6675 16758 6681
rect 16850 6672 16856 6684
rect 16908 6712 16914 6724
rect 17310 6712 17316 6724
rect 16908 6684 17316 6712
rect 16908 6672 16914 6684
rect 17310 6672 17316 6684
rect 17368 6672 17374 6724
rect 17880 6712 17908 6743
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 17880 6684 18920 6712
rect 9033 6647 9091 6653
rect 9033 6613 9045 6647
rect 9079 6644 9091 6647
rect 9122 6644 9128 6656
rect 9079 6616 9128 6644
rect 9079 6613 9091 6616
rect 9033 6607 9091 6613
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 12986 6644 12992 6656
rect 12947 6616 12992 6644
rect 12986 6604 12992 6616
rect 13044 6604 13050 6656
rect 13722 6604 13728 6656
rect 13780 6644 13786 6656
rect 15378 6644 15384 6656
rect 13780 6616 15384 6644
rect 13780 6604 13786 6616
rect 15378 6604 15384 6616
rect 15436 6644 15442 6656
rect 15473 6647 15531 6653
rect 15473 6644 15485 6647
rect 15436 6616 15485 6644
rect 15436 6604 15442 6616
rect 15473 6613 15485 6616
rect 15519 6613 15531 6647
rect 15473 6607 15531 6613
rect 15562 6604 15568 6656
rect 15620 6644 15626 6656
rect 15620 6616 15665 6644
rect 15620 6604 15626 6616
rect 16114 6604 16120 6656
rect 16172 6644 16178 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 16172 6616 17049 6644
rect 16172 6604 16178 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 17037 6607 17095 6613
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17405 6647 17463 6653
rect 17405 6644 17417 6647
rect 17276 6616 17417 6644
rect 17276 6604 17282 6616
rect 17405 6613 17417 6616
rect 17451 6613 17463 6647
rect 18414 6644 18420 6656
rect 18375 6616 18420 6644
rect 17405 6607 17463 6613
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 1104 6554 18860 6576
rect 1104 6502 5398 6554
rect 5450 6502 5462 6554
rect 5514 6502 5526 6554
rect 5578 6502 5590 6554
rect 5642 6502 5654 6554
rect 5706 6502 9846 6554
rect 9898 6502 9910 6554
rect 9962 6502 9974 6554
rect 10026 6502 10038 6554
rect 10090 6502 10102 6554
rect 10154 6502 14294 6554
rect 14346 6502 14358 6554
rect 14410 6502 14422 6554
rect 14474 6502 14486 6554
rect 14538 6502 14550 6554
rect 14602 6502 18860 6554
rect 1104 6480 18860 6502
rect 1118 6400 1124 6452
rect 1176 6440 1182 6452
rect 2777 6443 2835 6449
rect 2777 6440 2789 6443
rect 1176 6412 2789 6440
rect 1176 6400 1182 6412
rect 2777 6409 2789 6412
rect 2823 6409 2835 6443
rect 2777 6403 2835 6409
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 4341 6443 4399 6449
rect 4341 6440 4353 6443
rect 3660 6412 4353 6440
rect 3660 6400 3666 6412
rect 4341 6409 4353 6412
rect 4387 6409 4399 6443
rect 4341 6403 4399 6409
rect 4433 6443 4491 6449
rect 4433 6409 4445 6443
rect 4479 6440 4491 6443
rect 4614 6440 4620 6452
rect 4479 6412 4620 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 9582 6400 9588 6452
rect 9640 6400 9646 6452
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6409 10655 6443
rect 10597 6403 10655 6409
rect 10781 6443 10839 6449
rect 10781 6409 10793 6443
rect 10827 6440 10839 6443
rect 10962 6440 10968 6452
rect 10827 6412 10968 6440
rect 10827 6409 10839 6412
rect 10781 6403 10839 6409
rect 3789 6375 3847 6381
rect 3789 6372 3801 6375
rect 1688 6344 3801 6372
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 1688 6313 1716 6344
rect 3789 6341 3801 6344
rect 3835 6341 3847 6375
rect 3789 6335 3847 6341
rect 1673 6307 1731 6313
rect 1673 6304 1685 6307
rect 1544 6276 1685 6304
rect 1544 6264 1550 6276
rect 1673 6273 1685 6276
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6273 2099 6307
rect 2406 6304 2412 6316
rect 2367 6276 2412 6304
rect 2041 6267 2099 6273
rect 1302 6196 1308 6248
rect 1360 6236 1366 6248
rect 2056 6236 2084 6267
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6304 3203 6307
rect 3602 6304 3608 6316
rect 3191 6276 3608 6304
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 1360 6208 2084 6236
rect 1360 6196 1366 6208
rect 2130 6196 2136 6248
rect 2188 6236 2194 6248
rect 2314 6236 2320 6248
rect 2188 6208 2320 6236
rect 2188 6196 2194 6208
rect 2314 6196 2320 6208
rect 2372 6236 2378 6248
rect 3160 6236 3188 6267
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 3804 6304 3832 6335
rect 5718 6332 5724 6384
rect 5776 6372 5782 6384
rect 8386 6372 8392 6384
rect 5776 6344 8392 6372
rect 5776 6332 5782 6344
rect 8386 6332 8392 6344
rect 8444 6332 8450 6384
rect 9306 6332 9312 6384
rect 9364 6372 9370 6384
rect 9484 6375 9542 6381
rect 9484 6372 9496 6375
rect 9364 6344 9496 6372
rect 9364 6332 9370 6344
rect 9484 6341 9496 6344
rect 9530 6341 9542 6375
rect 9600 6372 9628 6400
rect 10612 6372 10640 6403
rect 10962 6400 10968 6412
rect 11020 6440 11026 6452
rect 11333 6443 11391 6449
rect 11333 6440 11345 6443
rect 11020 6412 11345 6440
rect 11020 6400 11026 6412
rect 11333 6409 11345 6412
rect 11379 6440 11391 6443
rect 11609 6443 11667 6449
rect 11609 6440 11621 6443
rect 11379 6412 11621 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 11609 6409 11621 6412
rect 11655 6440 11667 6443
rect 11977 6443 12035 6449
rect 11977 6440 11989 6443
rect 11655 6412 11989 6440
rect 11655 6409 11667 6412
rect 11609 6403 11667 6409
rect 11977 6409 11989 6412
rect 12023 6440 12035 6443
rect 12161 6443 12219 6449
rect 12161 6440 12173 6443
rect 12023 6412 12173 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 12161 6409 12173 6412
rect 12207 6440 12219 6443
rect 13357 6443 13415 6449
rect 13357 6440 13369 6443
rect 12207 6412 13369 6440
rect 12207 6409 12219 6412
rect 12161 6403 12219 6409
rect 13357 6409 13369 6412
rect 13403 6440 13415 6443
rect 13446 6440 13452 6452
rect 13403 6412 13452 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 14921 6443 14979 6449
rect 14921 6440 14933 6443
rect 14752 6412 14933 6440
rect 10686 6372 10692 6384
rect 9600 6344 10692 6372
rect 9484 6335 9542 6341
rect 10686 6332 10692 6344
rect 10744 6332 10750 6384
rect 12621 6375 12679 6381
rect 12621 6341 12633 6375
rect 12667 6372 12679 6375
rect 13538 6372 13544 6384
rect 12667 6344 13544 6372
rect 12667 6341 12679 6344
rect 12621 6335 12679 6341
rect 13538 6332 13544 6344
rect 13596 6332 13602 6384
rect 14584 6375 14642 6381
rect 14584 6341 14596 6375
rect 14630 6372 14642 6375
rect 14752 6372 14780 6412
rect 14921 6409 14933 6412
rect 14967 6440 14979 6443
rect 15102 6440 15108 6452
rect 14967 6412 15108 6440
rect 14967 6409 14979 6412
rect 14921 6403 14979 6409
rect 15102 6400 15108 6412
rect 15160 6400 15166 6452
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 16393 6443 16451 6449
rect 16393 6440 16405 6443
rect 15988 6412 16405 6440
rect 15988 6400 15994 6412
rect 16393 6409 16405 6412
rect 16439 6409 16451 6443
rect 17218 6440 17224 6452
rect 17179 6412 17224 6440
rect 16393 6403 16451 6409
rect 17218 6400 17224 6412
rect 17276 6400 17282 6452
rect 17681 6443 17739 6449
rect 17681 6409 17693 6443
rect 17727 6440 17739 6443
rect 18322 6440 18328 6452
rect 17727 6412 18328 6440
rect 17727 6409 17739 6412
rect 17681 6403 17739 6409
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 18414 6400 18420 6452
rect 18472 6440 18478 6452
rect 18892 6440 18920 6684
rect 18472 6412 18920 6440
rect 18472 6400 18478 6412
rect 15562 6372 15568 6384
rect 14630 6344 14780 6372
rect 14844 6344 15568 6372
rect 14630 6341 14642 6344
rect 14584 6335 14642 6341
rect 14844 6316 14872 6344
rect 15562 6332 15568 6344
rect 15620 6372 15626 6384
rect 17773 6375 17831 6381
rect 15620 6344 16344 6372
rect 15620 6332 15626 6344
rect 3804 6276 4292 6304
rect 2372 6208 3188 6236
rect 3237 6239 3295 6245
rect 2372 6196 2378 6208
rect 3237 6205 3249 6239
rect 3283 6205 3295 6239
rect 3418 6236 3424 6248
rect 3379 6208 3424 6236
rect 3237 6199 3295 6205
rect 2225 6171 2283 6177
rect 2225 6137 2237 6171
rect 2271 6168 2283 6171
rect 2958 6168 2964 6180
rect 2271 6140 2964 6168
rect 2271 6137 2283 6140
rect 2225 6131 2283 6137
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 3050 6128 3056 6180
rect 3108 6168 3114 6180
rect 3252 6168 3280 6199
rect 3418 6196 3424 6208
rect 3476 6196 3482 6248
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 4062 6236 4068 6248
rect 3936 6208 4068 6236
rect 3936 6196 3942 6208
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 3108 6140 3280 6168
rect 4264 6168 4292 6276
rect 4430 6264 4436 6316
rect 4488 6304 4494 6316
rect 5068 6307 5126 6313
rect 5068 6304 5080 6307
rect 4488 6276 5080 6304
rect 4488 6264 4494 6276
rect 5068 6273 5080 6276
rect 5114 6304 5126 6307
rect 6086 6304 6092 6316
rect 5114 6276 6092 6304
rect 5114 6273 5126 6276
rect 5068 6267 5126 6273
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 7357 6307 7415 6313
rect 7357 6304 7369 6307
rect 6196 6276 7369 6304
rect 4614 6236 4620 6248
rect 4575 6208 4620 6236
rect 4614 6196 4620 6208
rect 4672 6196 4678 6248
rect 4798 6236 4804 6248
rect 4759 6208 4804 6236
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 4522 6168 4528 6180
rect 4264 6140 4528 6168
rect 3108 6128 3114 6140
rect 4522 6128 4528 6140
rect 4580 6128 4586 6180
rect 5994 6128 6000 6180
rect 6052 6168 6058 6180
rect 6196 6177 6224 6276
rect 7357 6273 7369 6276
rect 7403 6273 7415 6307
rect 7357 6267 7415 6273
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 9122 6304 9128 6316
rect 8711 6276 9128 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 9122 6264 9128 6276
rect 9180 6304 9186 6316
rect 9217 6307 9275 6313
rect 9217 6304 9229 6307
rect 9180 6276 9229 6304
rect 9180 6264 9186 6276
rect 9217 6273 9229 6276
rect 9263 6273 9275 6307
rect 12894 6304 12900 6316
rect 9217 6267 9275 6273
rect 9324 6276 12900 6304
rect 7101 6239 7159 6245
rect 7101 6236 7113 6239
rect 6380 6208 7113 6236
rect 6181 6171 6239 6177
rect 6181 6168 6193 6171
rect 6052 6140 6193 6168
rect 6052 6128 6058 6140
rect 6181 6137 6193 6140
rect 6227 6137 6239 6171
rect 6181 6131 6239 6137
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1489 6103 1547 6109
rect 1489 6100 1501 6103
rect 1452 6072 1501 6100
rect 1452 6060 1458 6072
rect 1489 6069 1501 6072
rect 1535 6069 1547 6103
rect 1489 6063 1547 6069
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 1857 6103 1915 6109
rect 1857 6100 1869 6103
rect 1728 6072 1869 6100
rect 1728 6060 1734 6072
rect 1857 6069 1869 6072
rect 1903 6069 1915 6103
rect 1857 6063 1915 6069
rect 2685 6103 2743 6109
rect 2685 6069 2697 6103
rect 2731 6100 2743 6103
rect 3068 6100 3096 6128
rect 6380 6112 6408 6208
rect 7101 6205 7113 6208
rect 7147 6205 7159 6239
rect 7101 6199 7159 6205
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 9324 6236 9352 6276
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 14090 6304 14096 6316
rect 13044 6276 14096 6304
rect 13044 6264 13050 6276
rect 14090 6264 14096 6276
rect 14148 6304 14154 6316
rect 14148 6276 14780 6304
rect 14148 6264 14154 6276
rect 8996 6208 9352 6236
rect 14752 6236 14780 6276
rect 14826 6264 14832 6316
rect 14884 6304 14890 6316
rect 14884 6276 14977 6304
rect 14884 6264 14890 6276
rect 16022 6264 16028 6316
rect 16080 6313 16086 6316
rect 16316 6313 16344 6344
rect 17773 6341 17785 6375
rect 17819 6372 17831 6375
rect 18046 6372 18052 6384
rect 17819 6344 18052 6372
rect 17819 6341 17831 6344
rect 17773 6335 17831 6341
rect 18046 6332 18052 6344
rect 18104 6332 18110 6384
rect 16080 6304 16092 6313
rect 16301 6307 16359 6313
rect 16080 6276 16125 6304
rect 16080 6267 16092 6276
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 16390 6304 16396 6316
rect 16347 6276 16396 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 16080 6264 16086 6267
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 17494 6264 17500 6316
rect 17552 6304 17558 6316
rect 18141 6307 18199 6313
rect 18141 6304 18153 6307
rect 17552 6276 18153 6304
rect 17552 6264 17558 6276
rect 18141 6273 18153 6276
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 18230 6264 18236 6316
rect 18288 6304 18294 6316
rect 18325 6307 18383 6313
rect 18325 6304 18337 6307
rect 18288 6276 18337 6304
rect 18288 6264 18294 6276
rect 18325 6273 18337 6276
rect 18371 6273 18383 6307
rect 18325 6267 18383 6273
rect 14918 6236 14924 6248
rect 14752 6208 14924 6236
rect 8996 6196 9002 6208
rect 14918 6196 14924 6208
rect 14976 6196 14982 6248
rect 16758 6236 16764 6248
rect 16671 6208 16764 6236
rect 16758 6196 16764 6208
rect 16816 6236 16822 6248
rect 17862 6236 17868 6248
rect 16816 6208 17080 6236
rect 17823 6208 17868 6236
rect 16816 6196 16822 6208
rect 8110 6128 8116 6180
rect 8168 6168 8174 6180
rect 8481 6171 8539 6177
rect 8168 6140 8423 6168
rect 8168 6128 8174 6140
rect 2731 6072 3096 6100
rect 2731 6069 2743 6072
rect 2685 6063 2743 6069
rect 3878 6060 3884 6112
rect 3936 6100 3942 6112
rect 3973 6103 4031 6109
rect 3973 6100 3985 6103
rect 3936 6072 3985 6100
rect 3936 6060 3942 6072
rect 3973 6069 3985 6072
rect 4019 6069 4031 6103
rect 6362 6100 6368 6112
rect 6323 6072 6368 6100
rect 3973 6063 4031 6069
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6641 6103 6699 6109
rect 6641 6069 6653 6103
rect 6687 6100 6699 6103
rect 8294 6100 8300 6112
rect 6687 6072 8300 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 8395 6100 8423 6140
rect 8481 6137 8493 6171
rect 8527 6168 8539 6171
rect 9214 6168 9220 6180
rect 8527 6140 9220 6168
rect 8527 6137 8539 6140
rect 8481 6131 8539 6137
rect 9214 6128 9220 6140
rect 9272 6128 9278 6180
rect 10226 6128 10232 6180
rect 10284 6168 10290 6180
rect 13449 6171 13507 6177
rect 10284 6140 13032 6168
rect 10284 6128 10290 6140
rect 11698 6100 11704 6112
rect 8395 6072 11704 6100
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12805 6103 12863 6109
rect 12492 6072 12537 6100
rect 12492 6060 12498 6072
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 12894 6100 12900 6112
rect 12851 6072 12900 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13004 6109 13032 6140
rect 13449 6137 13461 6171
rect 13495 6168 13507 6171
rect 13814 6168 13820 6180
rect 13495 6140 13820 6168
rect 13495 6137 13507 6140
rect 13449 6131 13507 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 16574 6128 16580 6180
rect 16632 6168 16638 6180
rect 17052 6168 17080 6208
rect 17862 6196 17868 6208
rect 17920 6196 17926 6248
rect 18414 6168 18420 6180
rect 16632 6140 16988 6168
rect 17052 6140 18420 6168
rect 16632 6128 16638 6140
rect 12989 6103 13047 6109
rect 12989 6069 13001 6103
rect 13035 6100 13047 6103
rect 13170 6100 13176 6112
rect 13035 6072 13176 6100
rect 13035 6069 13047 6072
rect 12989 6063 13047 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 16960 6109 16988 6140
rect 18414 6128 18420 6140
rect 18472 6128 18478 6180
rect 16945 6103 17003 6109
rect 16945 6069 16957 6103
rect 16991 6100 17003 6103
rect 17126 6100 17132 6112
rect 16991 6072 17132 6100
rect 16991 6069 17003 6072
rect 16945 6063 17003 6069
rect 17126 6060 17132 6072
rect 17184 6060 17190 6112
rect 17310 6100 17316 6112
rect 17271 6072 17316 6100
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 1104 6010 18860 6032
rect 1104 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 3430 6010
rect 3482 5958 7622 6010
rect 7674 5958 7686 6010
rect 7738 5958 7750 6010
rect 7802 5958 7814 6010
rect 7866 5958 7878 6010
rect 7930 5958 12070 6010
rect 12122 5958 12134 6010
rect 12186 5958 12198 6010
rect 12250 5958 12262 6010
rect 12314 5958 12326 6010
rect 12378 5958 16518 6010
rect 16570 5958 16582 6010
rect 16634 5958 16646 6010
rect 16698 5958 16710 6010
rect 16762 5958 16774 6010
rect 16826 5958 18860 6010
rect 1104 5936 18860 5958
rect 1486 5896 1492 5908
rect 1447 5868 1492 5896
rect 1486 5856 1492 5868
rect 1544 5856 1550 5908
rect 2317 5899 2375 5905
rect 2317 5865 2329 5899
rect 2363 5896 2375 5899
rect 2406 5896 2412 5908
rect 2363 5868 2412 5896
rect 2363 5865 2375 5868
rect 2317 5859 2375 5865
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3145 5899 3203 5905
rect 3145 5896 3157 5899
rect 2924 5868 3157 5896
rect 2924 5856 2930 5868
rect 3145 5865 3157 5868
rect 3191 5865 3203 5899
rect 3602 5896 3608 5908
rect 3563 5868 3608 5896
rect 3145 5859 3203 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 11977 5899 12035 5905
rect 11977 5896 11989 5899
rect 4672 5868 11989 5896
rect 4672 5856 4678 5868
rect 11977 5865 11989 5868
rect 12023 5865 12035 5899
rect 11977 5859 12035 5865
rect 1504 5624 1532 5856
rect 2608 5800 4568 5828
rect 1946 5720 1952 5772
rect 2004 5760 2010 5772
rect 2608 5769 2636 5800
rect 2593 5763 2651 5769
rect 2004 5732 2544 5760
rect 2004 5720 2010 5732
rect 1854 5652 1860 5704
rect 1912 5692 1918 5704
rect 2041 5695 2099 5701
rect 2041 5692 2053 5695
rect 1912 5664 2053 5692
rect 1912 5652 1918 5664
rect 2041 5661 2053 5664
rect 2087 5661 2099 5695
rect 2516 5692 2544 5732
rect 2593 5729 2605 5763
rect 2639 5729 2651 5763
rect 2593 5723 2651 5729
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5760 2743 5763
rect 2774 5760 2780 5772
rect 2731 5732 2780 5760
rect 2731 5729 2743 5732
rect 2685 5723 2743 5729
rect 2774 5720 2780 5732
rect 2832 5720 2838 5772
rect 3973 5763 4031 5769
rect 3973 5729 3985 5763
rect 4019 5760 4031 5763
rect 4154 5760 4160 5772
rect 4019 5732 4160 5760
rect 4019 5729 4031 5732
rect 3973 5723 4031 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 3329 5695 3387 5701
rect 3329 5692 3341 5695
rect 2516 5664 3341 5692
rect 2041 5655 2099 5661
rect 3329 5661 3341 5664
rect 3375 5661 3387 5695
rect 3329 5655 3387 5661
rect 2777 5627 2835 5633
rect 2777 5624 2789 5627
rect 1504 5596 2789 5624
rect 2777 5593 2789 5596
rect 2823 5593 2835 5627
rect 3344 5624 3372 5655
rect 3602 5652 3608 5704
rect 3660 5692 3666 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3660 5664 4077 5692
rect 3660 5652 3666 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4157 5627 4215 5633
rect 4157 5624 4169 5627
rect 3344 5596 4169 5624
rect 2777 5587 2835 5593
rect 4157 5593 4169 5596
rect 4203 5624 4215 5627
rect 4430 5624 4436 5636
rect 4203 5596 4436 5624
rect 4203 5593 4215 5596
rect 4157 5587 4215 5593
rect 4430 5584 4436 5596
rect 4488 5584 4494 5636
rect 4540 5624 4568 5800
rect 5810 5788 5816 5840
rect 5868 5828 5874 5840
rect 5997 5831 6055 5837
rect 5997 5828 6009 5831
rect 5868 5800 6009 5828
rect 5868 5788 5874 5800
rect 5997 5797 6009 5800
rect 6043 5797 6055 5831
rect 5997 5791 6055 5797
rect 6086 5788 6092 5840
rect 6144 5828 6150 5840
rect 6144 5800 6189 5828
rect 6144 5788 6150 5800
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5760 4675 5763
rect 4663 5732 4752 5760
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 4724 5704 4752 5732
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 6362 5652 6368 5704
rect 6420 5692 6426 5704
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 6420 5664 7481 5692
rect 6420 5652 6426 5664
rect 7469 5661 7481 5664
rect 7515 5692 7527 5695
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 7515 5664 7573 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 7561 5661 7573 5664
rect 7607 5692 7619 5695
rect 7745 5695 7803 5701
rect 7745 5692 7757 5695
rect 7607 5664 7757 5692
rect 7607 5661 7619 5664
rect 7561 5655 7619 5661
rect 7745 5661 7757 5664
rect 7791 5692 7803 5695
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7791 5664 8125 5692
rect 7791 5661 7803 5664
rect 7745 5655 7803 5661
rect 8113 5661 8125 5664
rect 8159 5692 8171 5695
rect 9122 5692 9128 5704
rect 8159 5664 9128 5692
rect 8159 5661 8171 5664
rect 8113 5655 8171 5661
rect 9122 5652 9128 5664
rect 9180 5692 9186 5704
rect 10597 5695 10655 5701
rect 10597 5692 10609 5695
rect 9180 5664 10609 5692
rect 9180 5652 9186 5664
rect 10597 5661 10609 5664
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 4884 5627 4942 5633
rect 4540 5596 4743 5624
rect 1302 5516 1308 5568
rect 1360 5556 1366 5568
rect 1581 5559 1639 5565
rect 1581 5556 1593 5559
rect 1360 5528 1593 5556
rect 1360 5516 1366 5528
rect 1581 5525 1593 5528
rect 1627 5525 1639 5559
rect 1581 5519 1639 5525
rect 1762 5516 1768 5568
rect 1820 5556 1826 5568
rect 1857 5559 1915 5565
rect 1857 5556 1869 5559
rect 1820 5528 1869 5556
rect 1820 5516 1826 5528
rect 1857 5525 1869 5528
rect 1903 5525 1915 5559
rect 4522 5556 4528 5568
rect 4483 5528 4528 5556
rect 1857 5519 1915 5525
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 4715 5556 4743 5596
rect 4884 5593 4896 5627
rect 4930 5624 4942 5627
rect 5902 5624 5908 5636
rect 4930 5596 5908 5624
rect 4930 5593 4942 5596
rect 4884 5587 4942 5593
rect 5902 5584 5908 5596
rect 5960 5584 5966 5636
rect 7190 5584 7196 5636
rect 7248 5633 7254 5636
rect 7248 5624 7260 5633
rect 7248 5596 7293 5624
rect 7248 5587 7260 5596
rect 7248 5584 7254 5587
rect 8018 5584 8024 5636
rect 8076 5624 8082 5636
rect 9370 5627 9428 5633
rect 9370 5624 9382 5627
rect 8076 5596 9382 5624
rect 8076 5584 8082 5596
rect 9370 5593 9382 5596
rect 9416 5624 9428 5627
rect 9674 5624 9680 5636
rect 9416 5596 9680 5624
rect 9416 5593 9428 5596
rect 9370 5587 9428 5593
rect 9674 5584 9680 5596
rect 9732 5584 9738 5636
rect 10612 5624 10640 5655
rect 10686 5652 10692 5704
rect 10744 5692 10750 5704
rect 10864 5695 10922 5701
rect 10864 5692 10876 5695
rect 10744 5664 10876 5692
rect 10744 5652 10750 5664
rect 10864 5661 10876 5664
rect 10910 5661 10922 5695
rect 10864 5655 10922 5661
rect 10962 5624 10968 5636
rect 10612 5596 10968 5624
rect 10962 5584 10968 5596
rect 11020 5584 11026 5636
rect 11992 5624 12020 5859
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 12124 5868 12169 5896
rect 12124 5856 12130 5868
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 13725 5899 13783 5905
rect 13725 5896 13737 5899
rect 13504 5868 13737 5896
rect 13504 5856 13510 5868
rect 13725 5865 13737 5868
rect 13771 5896 13783 5899
rect 15562 5896 15568 5908
rect 13771 5868 15240 5896
rect 15523 5868 15568 5896
rect 13771 5865 13783 5868
rect 13725 5859 13783 5865
rect 15212 5828 15240 5868
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15712 5868 15761 5896
rect 15712 5856 15718 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 15749 5859 15807 5865
rect 15838 5856 15844 5908
rect 15896 5896 15902 5908
rect 15933 5899 15991 5905
rect 15933 5896 15945 5899
rect 15896 5868 15945 5896
rect 15896 5856 15902 5868
rect 15933 5865 15945 5868
rect 15979 5865 15991 5899
rect 17218 5896 17224 5908
rect 15933 5859 15991 5865
rect 16040 5868 17224 5896
rect 16040 5828 16068 5868
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 15212 5800 16068 5828
rect 16298 5720 16304 5772
rect 16356 5760 16362 5772
rect 16577 5763 16635 5769
rect 16577 5760 16589 5763
rect 16356 5732 16589 5760
rect 16356 5720 16362 5732
rect 16577 5729 16589 5732
rect 16623 5729 16635 5763
rect 16577 5723 16635 5729
rect 16761 5763 16819 5769
rect 16761 5729 16773 5763
rect 16807 5760 16819 5763
rect 16850 5760 16856 5772
rect 16807 5732 16856 5760
rect 16807 5729 16819 5732
rect 16761 5723 16819 5729
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 17494 5760 17500 5772
rect 17455 5732 17500 5760
rect 17494 5720 17500 5732
rect 17552 5720 17558 5772
rect 18325 5763 18383 5769
rect 18325 5729 18337 5763
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 13182 5695 13240 5701
rect 13182 5692 13194 5695
rect 12124 5664 13194 5692
rect 12124 5652 12130 5664
rect 13182 5661 13194 5664
rect 13228 5661 13240 5695
rect 13446 5692 13452 5704
rect 13359 5664 13452 5692
rect 13182 5655 13240 5661
rect 13446 5652 13452 5664
rect 13504 5692 13510 5704
rect 13909 5695 13967 5701
rect 13909 5692 13921 5695
rect 13504 5664 13921 5692
rect 13504 5652 13510 5664
rect 13909 5661 13921 5664
rect 13955 5692 13967 5695
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13955 5664 14105 5692
rect 13955 5661 13967 5664
rect 13909 5655 13967 5661
rect 14093 5661 14105 5664
rect 14139 5692 14151 5695
rect 14826 5692 14832 5704
rect 14139 5664 14832 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5692 16543 5695
rect 17310 5692 17316 5704
rect 16531 5664 17316 5692
rect 16531 5661 16543 5664
rect 16485 5655 16543 5661
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 13814 5624 13820 5636
rect 11992 5596 13820 5624
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 14360 5627 14418 5633
rect 14360 5593 14372 5627
rect 14406 5624 14418 5627
rect 15102 5624 15108 5636
rect 14406 5596 15108 5624
rect 14406 5593 14418 5596
rect 14360 5587 14418 5593
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 16758 5624 16764 5636
rect 15672 5596 16764 5624
rect 15672 5568 15700 5596
rect 16758 5584 16764 5596
rect 16816 5624 16822 5636
rect 17586 5624 17592 5636
rect 16816 5596 17592 5624
rect 16816 5584 16822 5596
rect 17586 5584 17592 5596
rect 17644 5624 17650 5636
rect 18340 5624 18368 5723
rect 17644 5596 18368 5624
rect 17644 5584 17650 5596
rect 5994 5556 6000 5568
rect 4715 5528 6000 5556
rect 5994 5516 6000 5528
rect 6052 5516 6058 5568
rect 6086 5516 6092 5568
rect 6144 5556 6150 5568
rect 10226 5556 10232 5568
rect 6144 5528 10232 5556
rect 6144 5516 6150 5528
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 10505 5559 10563 5565
rect 10505 5525 10517 5559
rect 10551 5556 10563 5559
rect 11882 5556 11888 5568
rect 10551 5528 11888 5556
rect 10551 5525 10563 5528
rect 10505 5519 10563 5525
rect 11882 5516 11888 5528
rect 11940 5556 11946 5568
rect 12066 5556 12072 5568
rect 11940 5528 12072 5556
rect 11940 5516 11946 5528
rect 12066 5516 12072 5528
rect 12124 5516 12130 5568
rect 15473 5559 15531 5565
rect 15473 5525 15485 5559
rect 15519 5556 15531 5559
rect 15654 5556 15660 5568
rect 15519 5528 15660 5556
rect 15519 5525 15531 5528
rect 15473 5519 15531 5525
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 16114 5556 16120 5568
rect 16075 5528 16120 5556
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 16206 5516 16212 5568
rect 16264 5556 16270 5568
rect 16945 5559 17003 5565
rect 16945 5556 16957 5559
rect 16264 5528 16957 5556
rect 16264 5516 16270 5528
rect 16945 5525 16957 5528
rect 16991 5525 17003 5559
rect 17310 5556 17316 5568
rect 17271 5528 17316 5556
rect 16945 5519 17003 5525
rect 17310 5516 17316 5528
rect 17368 5516 17374 5568
rect 17405 5559 17463 5565
rect 17405 5525 17417 5559
rect 17451 5556 17463 5559
rect 17773 5559 17831 5565
rect 17773 5556 17785 5559
rect 17451 5528 17785 5556
rect 17451 5525 17463 5528
rect 17405 5519 17463 5525
rect 17773 5525 17785 5528
rect 17819 5525 17831 5559
rect 18138 5556 18144 5568
rect 18099 5528 18144 5556
rect 17773 5519 17831 5525
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 18230 5516 18236 5568
rect 18288 5556 18294 5568
rect 18288 5528 18333 5556
rect 18288 5516 18294 5528
rect 1104 5466 18860 5488
rect 1104 5414 5398 5466
rect 5450 5414 5462 5466
rect 5514 5414 5526 5466
rect 5578 5414 5590 5466
rect 5642 5414 5654 5466
rect 5706 5414 9846 5466
rect 9898 5414 9910 5466
rect 9962 5414 9974 5466
rect 10026 5414 10038 5466
rect 10090 5414 10102 5466
rect 10154 5414 14294 5466
rect 14346 5414 14358 5466
rect 14410 5414 14422 5466
rect 14474 5414 14486 5466
rect 14538 5414 14550 5466
rect 14602 5414 18860 5466
rect 1104 5392 18860 5414
rect 2593 5355 2651 5361
rect 2593 5321 2605 5355
rect 2639 5352 2651 5355
rect 2774 5352 2780 5364
rect 2639 5324 2780 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 3970 5352 3976 5364
rect 3931 5324 3976 5352
rect 3970 5312 3976 5324
rect 4028 5312 4034 5364
rect 4065 5355 4123 5361
rect 4065 5321 4077 5355
rect 4111 5352 4123 5355
rect 4433 5355 4491 5361
rect 4433 5352 4445 5355
rect 4111 5324 4445 5352
rect 4111 5321 4123 5324
rect 4065 5315 4123 5321
rect 4433 5321 4445 5324
rect 4479 5321 4491 5355
rect 4433 5315 4491 5321
rect 4798 5312 4804 5364
rect 4856 5352 4862 5364
rect 6089 5355 6147 5361
rect 6089 5352 6101 5355
rect 4856 5324 6101 5352
rect 4856 5312 4862 5324
rect 6089 5321 6101 5324
rect 6135 5352 6147 5355
rect 6362 5352 6368 5364
rect 6135 5324 6368 5352
rect 6135 5321 6147 5324
rect 6089 5315 6147 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 6454 5312 6460 5364
rect 6512 5352 6518 5364
rect 13906 5352 13912 5364
rect 6512 5324 13912 5352
rect 6512 5312 6518 5324
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 14200 5324 15516 5352
rect 4154 5244 4160 5296
rect 4212 5284 4218 5296
rect 4706 5284 4712 5296
rect 4212 5256 4712 5284
rect 4212 5244 4218 5256
rect 4706 5244 4712 5256
rect 4764 5284 4770 5296
rect 4764 5256 5764 5284
rect 4764 5244 4770 5256
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2222 5216 2228 5228
rect 2087 5188 2228 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 1688 5148 1716 5179
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5216 2467 5219
rect 2498 5216 2504 5228
rect 2455 5188 2504 5216
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3145 5219 3203 5225
rect 3145 5216 3157 5219
rect 3108 5188 3157 5216
rect 3108 5176 3114 5188
rect 3145 5185 3157 5188
rect 3191 5216 3203 5219
rect 4338 5216 4344 5228
rect 3191 5188 4344 5216
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 4338 5176 4344 5188
rect 4396 5176 4402 5228
rect 4522 5176 4528 5228
rect 4580 5216 4586 5228
rect 4801 5219 4859 5225
rect 4801 5216 4813 5219
rect 4580 5188 4813 5216
rect 4580 5176 4586 5188
rect 4801 5185 4813 5188
rect 4847 5185 4859 5219
rect 5626 5216 5632 5228
rect 5587 5188 5632 5216
rect 4801 5179 4859 5185
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 5736 5216 5764 5256
rect 6380 5216 6408 5312
rect 9585 5287 9643 5293
rect 9585 5284 9597 5287
rect 6656 5256 9597 5284
rect 6656 5228 6684 5256
rect 6638 5216 6644 5228
rect 5736 5188 5856 5216
rect 6380 5188 6644 5216
rect 2682 5148 2688 5160
rect 1688 5120 2688 5148
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 3237 5151 3295 5157
rect 3237 5148 3249 5151
rect 2924 5120 3249 5148
rect 2924 5108 2930 5120
rect 3237 5117 3249 5120
rect 3283 5117 3295 5151
rect 3237 5111 3295 5117
rect 3421 5151 3479 5157
rect 3421 5117 3433 5151
rect 3467 5117 3479 5151
rect 3421 5111 3479 5117
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 4430 5148 4436 5160
rect 4295 5120 4436 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 3436 5080 3464 5111
rect 4430 5108 4436 5120
rect 4488 5108 4494 5160
rect 4893 5151 4951 5157
rect 4893 5117 4905 5151
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 4522 5080 4528 5092
rect 3436 5052 4528 5080
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 4908 5080 4936 5111
rect 4982 5108 4988 5160
rect 5040 5148 5046 5160
rect 5718 5148 5724 5160
rect 5040 5120 5085 5148
rect 5679 5120 5724 5148
rect 5040 5108 5046 5120
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 5828 5157 5856 5188
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 6914 5225 6920 5228
rect 6908 5216 6920 5225
rect 6875 5188 6920 5216
rect 6908 5179 6920 5188
rect 6914 5176 6920 5179
rect 6972 5176 6978 5228
rect 8128 5225 8156 5256
rect 9585 5253 9597 5256
rect 9631 5253 9643 5287
rect 9585 5247 9643 5253
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 9769 5287 9827 5293
rect 9769 5284 9781 5287
rect 9732 5256 9781 5284
rect 9732 5244 9738 5256
rect 9769 5253 9781 5256
rect 9815 5253 9827 5287
rect 10962 5284 10968 5296
rect 9769 5247 9827 5253
rect 9968 5256 10968 5284
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8380 5219 8438 5225
rect 8380 5185 8392 5219
rect 8426 5216 8438 5219
rect 8662 5216 8668 5228
rect 8426 5188 8668 5216
rect 8426 5185 8438 5188
rect 8380 5179 8438 5185
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5117 5871 5151
rect 9784 5148 9812 5247
rect 9968 5228 9996 5256
rect 10962 5244 10968 5256
rect 11020 5244 11026 5296
rect 11790 5293 11796 5296
rect 11784 5284 11796 5293
rect 11751 5256 11796 5284
rect 11784 5247 11796 5256
rect 11790 5244 11796 5247
rect 11848 5244 11854 5296
rect 13814 5244 13820 5296
rect 13872 5284 13878 5296
rect 14102 5287 14160 5293
rect 14102 5284 14114 5287
rect 13872 5256 14114 5284
rect 13872 5244 13878 5256
rect 14102 5253 14114 5256
rect 14148 5253 14160 5287
rect 14102 5247 14160 5253
rect 9950 5216 9956 5228
rect 9863 5188 9956 5216
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 10209 5219 10267 5225
rect 10209 5216 10221 5219
rect 10060 5188 10221 5216
rect 10060 5148 10088 5188
rect 10209 5185 10221 5188
rect 10255 5185 10267 5219
rect 10209 5179 10267 5185
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5216 11575 5219
rect 11606 5216 11612 5228
rect 11563 5188 11612 5216
rect 11563 5185 11575 5188
rect 11517 5179 11575 5185
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 13170 5176 13176 5228
rect 13228 5216 13234 5228
rect 14200 5216 14228 5324
rect 14826 5284 14832 5296
rect 14476 5256 14832 5284
rect 14476 5225 14504 5256
rect 14826 5244 14832 5256
rect 14884 5244 14890 5296
rect 15488 5284 15516 5324
rect 15562 5312 15568 5364
rect 15620 5352 15626 5364
rect 15933 5355 15991 5361
rect 15933 5352 15945 5355
rect 15620 5324 15945 5352
rect 15620 5312 15626 5324
rect 15933 5321 15945 5324
rect 15979 5321 15991 5355
rect 16390 5352 16396 5364
rect 16351 5324 16396 5352
rect 15933 5315 15991 5321
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 17310 5312 17316 5364
rect 17368 5352 17374 5364
rect 17405 5355 17463 5361
rect 17405 5352 17417 5355
rect 17368 5324 17417 5352
rect 17368 5312 17374 5324
rect 17405 5321 17417 5324
rect 17451 5321 17463 5355
rect 18230 5352 18236 5364
rect 18191 5324 18236 5352
rect 17405 5315 17463 5321
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 18322 5312 18328 5364
rect 18380 5352 18386 5364
rect 18380 5324 18425 5352
rect 18380 5312 18386 5324
rect 15488 5256 15608 5284
rect 13228 5188 14228 5216
rect 14369 5219 14427 5225
rect 13228 5176 13234 5188
rect 14369 5185 14381 5219
rect 14415 5216 14427 5219
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 14415 5188 14473 5216
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 14728 5219 14786 5225
rect 14728 5185 14740 5219
rect 14774 5216 14786 5219
rect 15470 5216 15476 5228
rect 14774 5188 15476 5216
rect 14774 5185 14786 5188
rect 14728 5179 14786 5185
rect 15470 5176 15476 5188
rect 15528 5176 15534 5228
rect 15580 5216 15608 5256
rect 16942 5244 16948 5296
rect 17000 5284 17006 5296
rect 17494 5284 17500 5296
rect 17000 5256 17500 5284
rect 17000 5244 17006 5256
rect 17494 5244 17500 5256
rect 17552 5284 17558 5296
rect 17773 5287 17831 5293
rect 17773 5284 17785 5287
rect 17552 5256 17785 5284
rect 17552 5244 17558 5256
rect 17773 5253 17785 5256
rect 17819 5253 17831 5287
rect 17773 5247 17831 5253
rect 16298 5216 16304 5228
rect 15580 5188 16304 5216
rect 16298 5176 16304 5188
rect 16356 5216 16362 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 16356 5188 17049 5216
rect 16356 5176 16362 5188
rect 17037 5185 17049 5188
rect 17083 5216 17095 5219
rect 17402 5216 17408 5228
rect 17083 5188 17408 5216
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 17865 5219 17923 5225
rect 17865 5216 17877 5219
rect 17696 5188 17877 5216
rect 16758 5148 16764 5160
rect 9784 5120 10088 5148
rect 12820 5120 13400 5148
rect 16719 5120 16764 5148
rect 5813 5111 5871 5117
rect 5261 5083 5319 5089
rect 5261 5080 5273 5083
rect 4908 5052 5273 5080
rect 5261 5049 5273 5052
rect 5307 5049 5319 5083
rect 8018 5080 8024 5092
rect 7979 5052 8024 5080
rect 5261 5043 5319 5049
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 9398 5040 9404 5092
rect 9456 5080 9462 5092
rect 9493 5083 9551 5089
rect 9493 5080 9505 5083
rect 9456 5052 9505 5080
rect 9456 5040 9462 5052
rect 9493 5049 9505 5052
rect 9539 5049 9551 5083
rect 9493 5043 9551 5049
rect 1486 5012 1492 5024
rect 1447 4984 1492 5012
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 1854 5012 1860 5024
rect 1815 4984 1860 5012
rect 1854 4972 1860 4984
rect 1912 4972 1918 5024
rect 2222 5012 2228 5024
rect 2183 4984 2228 5012
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 3605 5015 3663 5021
rect 2832 4984 2877 5012
rect 2832 4972 2838 4984
rect 3605 4981 3617 5015
rect 3651 5012 3663 5015
rect 3786 5012 3792 5024
rect 3651 4984 3792 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 4338 4972 4344 5024
rect 4396 5012 4402 5024
rect 5626 5012 5632 5024
rect 4396 4984 5632 5012
rect 4396 4972 4402 4984
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 11333 5015 11391 5021
rect 11333 4981 11345 5015
rect 11379 5012 11391 5015
rect 12820 5012 12848 5120
rect 12897 5083 12955 5089
rect 12897 5049 12909 5083
rect 12943 5080 12955 5083
rect 13078 5080 13084 5092
rect 12943 5052 13084 5080
rect 12943 5049 12955 5052
rect 12897 5043 12955 5049
rect 13078 5040 13084 5052
rect 13136 5040 13142 5092
rect 11379 4984 12848 5012
rect 11379 4981 11391 4984
rect 11333 4975 11391 4981
rect 12986 4972 12992 5024
rect 13044 5012 13050 5024
rect 13372 5012 13400 5120
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 16942 5148 16948 5160
rect 16903 5120 16948 5148
rect 16942 5108 16948 5120
rect 17000 5108 17006 5160
rect 17310 5108 17316 5160
rect 17368 5148 17374 5160
rect 17589 5151 17647 5157
rect 17589 5148 17601 5151
rect 17368 5120 17601 5148
rect 17368 5108 17374 5120
rect 17589 5117 17601 5120
rect 17635 5117 17647 5151
rect 17589 5111 17647 5117
rect 15841 5083 15899 5089
rect 15841 5049 15853 5083
rect 15887 5080 15899 5083
rect 16022 5080 16028 5092
rect 15887 5052 16028 5080
rect 15887 5049 15899 5052
rect 15841 5043 15899 5049
rect 16022 5040 16028 5052
rect 16080 5040 16086 5092
rect 16666 5080 16672 5092
rect 16132 5052 16672 5080
rect 16132 5012 16160 5052
rect 16666 5040 16672 5052
rect 16724 5040 16730 5092
rect 17218 5040 17224 5092
rect 17276 5080 17282 5092
rect 17696 5080 17724 5188
rect 17865 5185 17877 5188
rect 17911 5216 17923 5219
rect 18322 5216 18328 5228
rect 17911 5188 18328 5216
rect 17911 5185 17923 5188
rect 17865 5179 17923 5185
rect 18322 5176 18328 5188
rect 18380 5176 18386 5228
rect 17276 5052 17724 5080
rect 17276 5040 17282 5052
rect 13044 4984 13089 5012
rect 13372 4984 16160 5012
rect 16301 5015 16359 5021
rect 13044 4972 13050 4984
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 19150 5012 19156 5024
rect 16347 4984 19156 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 1104 4922 18860 4944
rect 1104 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 3430 4922
rect 3482 4870 7622 4922
rect 7674 4870 7686 4922
rect 7738 4870 7750 4922
rect 7802 4870 7814 4922
rect 7866 4870 7878 4922
rect 7930 4870 12070 4922
rect 12122 4870 12134 4922
rect 12186 4870 12198 4922
rect 12250 4870 12262 4922
rect 12314 4870 12326 4922
rect 12378 4870 16518 4922
rect 16570 4870 16582 4922
rect 16634 4870 16646 4922
rect 16698 4870 16710 4922
rect 16762 4870 16774 4922
rect 16826 4870 18860 4922
rect 1104 4848 18860 4870
rect 1765 4811 1823 4817
rect 1765 4777 1777 4811
rect 1811 4808 1823 4811
rect 1946 4808 1952 4820
rect 1811 4780 1952 4808
rect 1811 4777 1823 4780
rect 1765 4771 1823 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2866 4808 2872 4820
rect 2827 4780 2872 4808
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 4338 4808 4344 4820
rect 4299 4780 4344 4808
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 5074 4768 5080 4820
rect 5132 4808 5138 4820
rect 5813 4811 5871 4817
rect 5813 4808 5825 4811
rect 5132 4780 5825 4808
rect 5132 4768 5138 4780
rect 5813 4777 5825 4780
rect 5859 4808 5871 4811
rect 8018 4808 8024 4820
rect 5859 4780 8024 4808
rect 5859 4777 5871 4780
rect 5813 4771 5871 4777
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 8846 4768 8852 4820
rect 8904 4808 8910 4820
rect 9769 4811 9827 4817
rect 9769 4808 9781 4811
rect 8904 4780 9781 4808
rect 8904 4768 8910 4780
rect 9769 4777 9781 4780
rect 9815 4777 9827 4811
rect 9950 4808 9956 4820
rect 9911 4780 9956 4808
rect 9769 4771 9827 4777
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 10226 4768 10232 4820
rect 10284 4808 10290 4820
rect 10410 4808 10416 4820
rect 10284 4780 10416 4808
rect 10284 4768 10290 4780
rect 10410 4768 10416 4780
rect 10468 4808 10474 4820
rect 12986 4808 12992 4820
rect 10468 4780 12992 4808
rect 10468 4768 10474 4780
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 13265 4811 13323 4817
rect 13265 4777 13277 4811
rect 13311 4808 13323 4811
rect 13446 4808 13452 4820
rect 13311 4780 13452 4808
rect 13311 4777 13323 4780
rect 13265 4771 13323 4777
rect 13446 4768 13452 4780
rect 13504 4808 13510 4820
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13504 4780 13645 4808
rect 13504 4768 13510 4780
rect 13633 4777 13645 4780
rect 13679 4808 13691 4811
rect 13817 4811 13875 4817
rect 13817 4808 13829 4811
rect 13679 4780 13829 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 13817 4777 13829 4780
rect 13863 4777 13875 4811
rect 13817 4771 13875 4777
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 14139 4780 16160 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 3050 4740 3056 4752
rect 1627 4712 3056 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 3050 4700 3056 4712
rect 3108 4700 3114 4752
rect 3418 4740 3424 4752
rect 3331 4712 3424 4740
rect 2130 4672 2136 4684
rect 2091 4644 2136 4672
rect 2130 4632 2136 4644
rect 2188 4632 2194 4684
rect 2317 4675 2375 4681
rect 2317 4641 2329 4675
rect 2363 4672 2375 4675
rect 2774 4672 2780 4684
rect 2363 4644 2780 4672
rect 2363 4641 2375 4644
rect 2317 4635 2375 4641
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 3344 4681 3372 4712
rect 3418 4700 3424 4712
rect 3476 4740 3482 4752
rect 4062 4740 4068 4752
rect 3476 4712 4068 4740
rect 3476 4700 3482 4712
rect 4062 4700 4068 4712
rect 4120 4700 4126 4752
rect 5902 4740 5908 4752
rect 5863 4712 5908 4740
rect 5902 4700 5908 4712
rect 5960 4700 5966 4752
rect 8757 4743 8815 4749
rect 8757 4709 8769 4743
rect 8803 4740 8815 4743
rect 9674 4740 9680 4752
rect 8803 4712 9680 4740
rect 8803 4709 8815 4712
rect 8757 4703 8815 4709
rect 9674 4700 9680 4712
rect 9732 4700 9738 4752
rect 10045 4743 10103 4749
rect 10045 4709 10057 4743
rect 10091 4709 10103 4743
rect 10045 4703 10103 4709
rect 3329 4675 3387 4681
rect 3329 4641 3341 4675
rect 3375 4641 3387 4675
rect 3329 4635 3387 4641
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4672 3571 4675
rect 3559 4644 4384 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4604 2007 4607
rect 4065 4607 4123 4613
rect 1995 4576 3280 4604
rect 1995 4573 2007 4576
rect 1949 4567 2007 4573
rect 3252 4548 3280 4576
rect 4065 4573 4077 4607
rect 4111 4604 4123 4607
rect 4246 4604 4252 4616
rect 4111 4576 4252 4604
rect 4111 4573 4123 4576
rect 4065 4567 4123 4573
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 2409 4539 2467 4545
rect 2409 4505 2421 4539
rect 2455 4536 2467 4539
rect 2958 4536 2964 4548
rect 2455 4508 2964 4536
rect 2455 4505 2467 4508
rect 2409 4499 2467 4505
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 3234 4536 3240 4548
rect 3195 4508 3240 4536
rect 3234 4496 3240 4508
rect 3292 4496 3298 4548
rect 2777 4471 2835 4477
rect 2777 4437 2789 4471
rect 2823 4468 2835 4471
rect 3050 4468 3056 4480
rect 2823 4440 3056 4468
rect 2823 4437 2835 4440
rect 2777 4431 2835 4437
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 3881 4471 3939 4477
rect 3881 4437 3893 4471
rect 3927 4468 3939 4471
rect 4062 4468 4068 4480
rect 3927 4440 4068 4468
rect 3927 4437 3939 4440
rect 3881 4431 3939 4437
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 4356 4468 4384 4644
rect 9306 4632 9312 4684
rect 9364 4672 9370 4684
rect 10060 4672 10088 4703
rect 13538 4700 13544 4752
rect 13596 4740 13602 4752
rect 14108 4740 14136 4771
rect 13596 4712 14136 4740
rect 13596 4700 13602 4712
rect 9364 4644 10088 4672
rect 15473 4675 15531 4681
rect 9364 4632 9370 4644
rect 15473 4641 15485 4675
rect 15519 4672 15531 4675
rect 15562 4672 15568 4684
rect 15519 4644 15568 4672
rect 15519 4641 15531 4644
rect 15473 4635 15531 4641
rect 15562 4632 15568 4644
rect 15620 4632 15626 4684
rect 16132 4681 16160 4780
rect 17034 4768 17040 4820
rect 17092 4808 17098 4820
rect 17586 4808 17592 4820
rect 17092 4780 17592 4808
rect 17092 4768 17098 4780
rect 17586 4768 17592 4780
rect 17644 4768 17650 4820
rect 17957 4811 18015 4817
rect 17957 4777 17969 4811
rect 18003 4808 18015 4811
rect 18138 4808 18144 4820
rect 18003 4780 18144 4808
rect 18003 4777 18015 4780
rect 17957 4771 18015 4777
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 18414 4808 18420 4820
rect 18375 4780 18420 4808
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 16117 4675 16175 4681
rect 15672 4644 16068 4672
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4479 4576 4844 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 4816 4548 4844 4576
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 6696 4576 7297 4604
rect 6696 4564 6702 4576
rect 7285 4573 7297 4576
rect 7331 4604 7343 4607
rect 7377 4607 7435 4613
rect 7377 4604 7389 4607
rect 7331 4576 7389 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 7377 4573 7389 4576
rect 7423 4573 7435 4607
rect 7377 4567 7435 4573
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 7644 4607 7702 4613
rect 7644 4604 7656 4607
rect 7524 4576 7656 4604
rect 7524 4564 7530 4576
rect 7644 4573 7656 4576
rect 7690 4604 7702 4607
rect 8478 4604 8484 4616
rect 7690 4576 8484 4604
rect 7690 4573 7702 4576
rect 7644 4567 7702 4573
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 9398 4604 9404 4616
rect 9359 4576 9404 4604
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4604 9643 4607
rect 9766 4604 9772 4616
rect 9631 4576 9772 4604
rect 9631 4573 9643 4576
rect 9585 4567 9643 4573
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4604 11483 4607
rect 11701 4607 11759 4613
rect 11701 4604 11713 4607
rect 11471 4576 11713 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 4706 4545 4712 4548
rect 4700 4536 4712 4545
rect 4667 4508 4712 4536
rect 4700 4499 4712 4508
rect 4706 4496 4712 4499
rect 4764 4496 4770 4548
rect 4798 4496 4804 4548
rect 4856 4496 4862 4548
rect 6914 4536 6920 4548
rect 5920 4508 6920 4536
rect 5920 4468 5948 4508
rect 6914 4496 6920 4508
rect 6972 4496 6978 4548
rect 7006 4496 7012 4548
rect 7064 4545 7070 4548
rect 7064 4536 7076 4545
rect 9125 4539 9183 4545
rect 7064 4508 7109 4536
rect 7064 4499 7076 4508
rect 9125 4505 9137 4539
rect 9171 4536 9183 4539
rect 9490 4536 9496 4548
rect 9171 4508 9496 4536
rect 9171 4505 9183 4508
rect 9125 4499 9183 4505
rect 7064 4496 7070 4499
rect 9490 4496 9496 4508
rect 9548 4496 9554 4548
rect 10410 4536 10416 4548
rect 9646 4508 10416 4536
rect 4356 4440 5948 4468
rect 5994 4428 6000 4480
rect 6052 4468 6058 4480
rect 9646 4468 9674 4508
rect 10410 4496 10416 4508
rect 10468 4536 10474 4548
rect 11158 4539 11216 4545
rect 11158 4536 11170 4539
rect 10468 4508 11170 4536
rect 10468 4496 10474 4508
rect 11158 4505 11170 4508
rect 11204 4505 11216 4539
rect 11158 4499 11216 4505
rect 11624 4480 11652 4576
rect 11701 4573 11713 4576
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 12894 4564 12900 4616
rect 12952 4604 12958 4616
rect 15672 4604 15700 4644
rect 12952 4576 15700 4604
rect 12952 4564 12958 4576
rect 15746 4564 15752 4616
rect 15804 4604 15810 4616
rect 15933 4607 15991 4613
rect 15933 4604 15945 4607
rect 15804 4576 15945 4604
rect 15804 4564 15810 4576
rect 15933 4573 15945 4576
rect 15979 4573 15991 4607
rect 16040 4604 16068 4644
rect 16117 4641 16129 4675
rect 16163 4641 16175 4675
rect 16117 4635 16175 4641
rect 16666 4632 16672 4684
rect 16724 4672 16730 4684
rect 16850 4672 16856 4684
rect 16724 4644 16856 4672
rect 16724 4632 16730 4644
rect 16850 4632 16856 4644
rect 16908 4672 16914 4684
rect 16945 4675 17003 4681
rect 16945 4672 16957 4675
rect 16908 4644 16957 4672
rect 16908 4632 16914 4644
rect 16945 4641 16957 4644
rect 16991 4672 17003 4675
rect 17034 4672 17040 4684
rect 16991 4644 17040 4672
rect 16991 4641 17003 4644
rect 16945 4635 17003 4641
rect 17034 4632 17040 4644
rect 17092 4632 17098 4684
rect 17310 4672 17316 4684
rect 17271 4644 17316 4672
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 17586 4604 17592 4616
rect 16040 4576 17356 4604
rect 17547 4576 17592 4604
rect 15933 4567 15991 4573
rect 11968 4539 12026 4545
rect 11968 4505 11980 4539
rect 12014 4536 12026 4539
rect 14090 4536 14096 4548
rect 12014 4508 14096 4536
rect 12014 4505 12026 4508
rect 11968 4499 12026 4505
rect 14090 4496 14096 4508
rect 14148 4496 14154 4548
rect 15194 4496 15200 4548
rect 15252 4545 15258 4548
rect 15252 4536 15264 4545
rect 16666 4536 16672 4548
rect 15252 4508 15297 4536
rect 15488 4508 16672 4536
rect 15252 4499 15264 4508
rect 15252 4496 15258 4499
rect 11606 4468 11612 4480
rect 6052 4440 9674 4468
rect 11567 4440 11612 4468
rect 6052 4428 6058 4440
rect 11606 4428 11612 4440
rect 11664 4428 11670 4480
rect 13081 4471 13139 4477
rect 13081 4437 13093 4471
rect 13127 4468 13139 4471
rect 15488 4468 15516 4508
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 16761 4539 16819 4545
rect 16761 4505 16773 4539
rect 16807 4536 16819 4539
rect 17218 4536 17224 4548
rect 16807 4508 17224 4536
rect 16807 4505 16819 4508
rect 16761 4499 16819 4505
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 17328 4536 17356 4576
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4604 18107 4607
rect 18506 4604 18512 4616
rect 18095 4576 18512 4604
rect 18095 4573 18107 4576
rect 18049 4567 18107 4573
rect 18506 4564 18512 4576
rect 18564 4604 18570 4616
rect 19242 4604 19248 4616
rect 18564 4576 19248 4604
rect 18564 4564 18570 4576
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 17770 4536 17776 4548
rect 17328 4508 17776 4536
rect 17770 4496 17776 4508
rect 17828 4496 17834 4548
rect 13127 4440 15516 4468
rect 15565 4471 15623 4477
rect 13127 4437 13139 4440
rect 13081 4431 13139 4437
rect 15565 4437 15577 4471
rect 15611 4468 15623 4471
rect 15930 4468 15936 4480
rect 15611 4440 15936 4468
rect 15611 4437 15623 4440
rect 15565 4431 15623 4437
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 16025 4471 16083 4477
rect 16025 4437 16037 4471
rect 16071 4468 16083 4471
rect 16206 4468 16212 4480
rect 16071 4440 16212 4468
rect 16071 4437 16083 4440
rect 16025 4431 16083 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 16390 4468 16396 4480
rect 16351 4440 16396 4468
rect 16390 4428 16396 4440
rect 16448 4428 16454 4480
rect 16850 4428 16856 4480
rect 16908 4468 16914 4480
rect 16908 4440 16953 4468
rect 16908 4428 16914 4440
rect 17126 4428 17132 4480
rect 17184 4468 17190 4480
rect 17497 4471 17555 4477
rect 17497 4468 17509 4471
rect 17184 4440 17509 4468
rect 17184 4428 17190 4440
rect 17497 4437 17509 4440
rect 17543 4437 17555 4471
rect 18230 4468 18236 4480
rect 18191 4440 18236 4468
rect 17497 4431 17555 4437
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 1104 4378 18860 4400
rect 1104 4326 5398 4378
rect 5450 4326 5462 4378
rect 5514 4326 5526 4378
rect 5578 4326 5590 4378
rect 5642 4326 5654 4378
rect 5706 4326 9846 4378
rect 9898 4326 9910 4378
rect 9962 4326 9974 4378
rect 10026 4326 10038 4378
rect 10090 4326 10102 4378
rect 10154 4326 14294 4378
rect 14346 4326 14358 4378
rect 14410 4326 14422 4378
rect 14474 4326 14486 4378
rect 14538 4326 14550 4378
rect 14602 4326 18860 4378
rect 1104 4304 18860 4326
rect 2685 4267 2743 4273
rect 2685 4233 2697 4267
rect 2731 4264 2743 4267
rect 2869 4267 2927 4273
rect 2869 4264 2881 4267
rect 2731 4236 2881 4264
rect 2731 4233 2743 4236
rect 2685 4227 2743 4233
rect 2869 4233 2881 4236
rect 2915 4264 2927 4267
rect 3053 4267 3111 4273
rect 3053 4264 3065 4267
rect 2915 4236 3065 4264
rect 2915 4233 2927 4236
rect 2869 4227 2927 4233
rect 3053 4233 3065 4236
rect 3099 4264 3111 4267
rect 3234 4264 3240 4276
rect 3099 4236 3240 4264
rect 3099 4233 3111 4236
rect 3053 4227 3111 4233
rect 3234 4224 3240 4236
rect 3292 4264 3298 4276
rect 4246 4264 4252 4276
rect 3292 4236 4252 4264
rect 3292 4224 3298 4236
rect 1489 4199 1547 4205
rect 1489 4165 1501 4199
rect 1535 4196 1547 4199
rect 1578 4196 1584 4208
rect 1535 4168 1584 4196
rect 1535 4165 1547 4168
rect 1489 4159 1547 4165
rect 1578 4156 1584 4168
rect 1636 4196 1642 4208
rect 1673 4199 1731 4205
rect 1673 4196 1685 4199
rect 1636 4168 1685 4196
rect 1636 4156 1642 4168
rect 1673 4165 1685 4168
rect 1719 4196 1731 4199
rect 3418 4196 3424 4208
rect 1719 4168 3424 4196
rect 1719 4165 1731 4168
rect 1673 4159 1731 4165
rect 3418 4156 3424 4168
rect 3476 4156 3482 4208
rect 3528 4205 3556 4236
rect 4246 4224 4252 4236
rect 4304 4264 4310 4276
rect 4341 4267 4399 4273
rect 4341 4264 4353 4267
rect 4304 4236 4353 4264
rect 4304 4224 4310 4236
rect 4341 4233 4353 4236
rect 4387 4233 4399 4267
rect 4341 4227 4399 4233
rect 6730 4224 6736 4276
rect 6788 4264 6794 4276
rect 8389 4267 8447 4273
rect 8389 4264 8401 4267
rect 6788 4236 8401 4264
rect 6788 4224 6794 4236
rect 8389 4233 8401 4236
rect 8435 4264 8447 4267
rect 9306 4264 9312 4276
rect 8435 4236 9312 4264
rect 8435 4233 8447 4236
rect 8389 4227 8447 4233
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 11606 4264 11612 4276
rect 11519 4236 11612 4264
rect 11606 4224 11612 4236
rect 11664 4264 11670 4276
rect 11793 4267 11851 4273
rect 11793 4264 11805 4267
rect 11664 4236 11805 4264
rect 11664 4224 11670 4236
rect 11793 4233 11805 4236
rect 11839 4264 11851 4267
rect 11977 4267 12035 4273
rect 11977 4264 11989 4267
rect 11839 4236 11989 4264
rect 11839 4233 11851 4236
rect 11793 4227 11851 4233
rect 11977 4233 11989 4236
rect 12023 4264 12035 4267
rect 13446 4264 13452 4276
rect 12023 4236 13452 4264
rect 12023 4233 12035 4236
rect 11977 4227 12035 4233
rect 13446 4224 13452 4236
rect 13504 4264 13510 4276
rect 13633 4267 13691 4273
rect 13633 4264 13645 4267
rect 13504 4236 13645 4264
rect 13504 4224 13510 4236
rect 3513 4199 3571 4205
rect 3513 4165 3525 4199
rect 3559 4165 3571 4199
rect 3513 4159 3571 4165
rect 4154 4156 4160 4208
rect 4212 4196 4218 4208
rect 9582 4205 9588 4208
rect 9524 4199 9588 4205
rect 4212 4168 4292 4196
rect 4212 4156 4218 4168
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2590 4128 2596 4140
rect 2455 4100 2596 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 4264 4137 4292 4168
rect 9524 4165 9536 4199
rect 9570 4165 9588 4199
rect 9524 4159 9588 4165
rect 9582 4156 9588 4159
rect 9640 4156 9646 4208
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 5068 4131 5126 4137
rect 5068 4128 5080 4131
rect 4488 4100 5080 4128
rect 4488 4088 4494 4100
rect 5068 4097 5080 4100
rect 5114 4128 5126 4131
rect 5114 4100 5856 4128
rect 5114 4097 5126 4100
rect 5068 4091 5126 4097
rect 3329 4063 3387 4069
rect 3329 4029 3341 4063
rect 3375 4029 3387 4063
rect 4154 4060 4160 4072
rect 4115 4032 4160 4060
rect 3329 4023 3387 4029
rect 3344 3992 3372 4023
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 4798 4060 4804 4072
rect 4759 4032 4804 4060
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 4614 3992 4620 4004
rect 3344 3964 4620 3992
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 5828 3992 5856 4100
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 6236 4100 6377 4128
rect 6236 4088 6242 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 8018 4088 8024 4140
rect 8076 4137 8082 4140
rect 8076 4128 8088 4137
rect 9766 4128 9772 4140
rect 8076 4100 8121 4128
rect 9727 4100 9772 4128
rect 8076 4091 8088 4100
rect 8076 4088 8082 4091
rect 9766 4088 9772 4100
rect 9824 4128 9830 4140
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 9824 4100 9873 4128
rect 9824 4088 9830 4100
rect 9861 4097 9873 4100
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 10117 4131 10175 4137
rect 10117 4128 10129 4131
rect 10008 4100 10129 4128
rect 10008 4088 10014 4100
rect 10117 4097 10129 4100
rect 10163 4097 10175 4131
rect 10117 4091 10175 4097
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 13556 4137 13584 4236
rect 13633 4233 13645 4236
rect 13679 4233 13691 4267
rect 13633 4227 13691 4233
rect 16025 4267 16083 4273
rect 16025 4233 16037 4267
rect 16071 4264 16083 4267
rect 16390 4264 16396 4276
rect 16071 4236 16396 4264
rect 16071 4233 16083 4236
rect 16025 4227 16083 4233
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 16942 4224 16948 4276
rect 17000 4264 17006 4276
rect 17129 4267 17187 4273
rect 17129 4264 17141 4267
rect 17000 4236 17141 4264
rect 17000 4224 17006 4236
rect 17129 4233 17141 4236
rect 17175 4233 17187 4267
rect 17129 4227 17187 4233
rect 17497 4267 17555 4273
rect 17497 4233 17509 4267
rect 17543 4264 17555 4267
rect 17770 4264 17776 4276
rect 17543 4236 17776 4264
rect 17543 4233 17555 4236
rect 17497 4227 17555 4233
rect 17770 4224 17776 4236
rect 17828 4224 17834 4276
rect 18138 4264 18144 4276
rect 18099 4236 18144 4264
rect 18138 4224 18144 4236
rect 18196 4224 18202 4276
rect 15933 4199 15991 4205
rect 15933 4165 15945 4199
rect 15979 4196 15991 4199
rect 16114 4196 16120 4208
rect 15979 4168 16120 4196
rect 15979 4165 15991 4168
rect 15933 4159 15991 4165
rect 16114 4156 16120 4168
rect 16172 4156 16178 4208
rect 16408 4168 17632 4196
rect 13274 4131 13332 4137
rect 13274 4128 13286 4131
rect 12860 4100 13286 4128
rect 12860 4088 12866 4100
rect 13274 4097 13286 4100
rect 13320 4128 13332 4131
rect 13541 4131 13599 4137
rect 13320 4100 13492 4128
rect 13320 4097 13332 4100
rect 13274 4091 13332 4097
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 8297 4063 8355 4069
rect 6687 4032 7328 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 6917 3995 6975 4001
rect 6917 3992 6929 3995
rect 5828 3964 6929 3992
rect 6917 3961 6929 3964
rect 6963 3961 6975 3995
rect 6917 3955 6975 3961
rect 1670 3884 1676 3936
rect 1728 3924 1734 3936
rect 1857 3927 1915 3933
rect 1857 3924 1869 3927
rect 1728 3896 1869 3924
rect 1728 3884 1734 3896
rect 1857 3893 1869 3896
rect 1903 3893 1915 3927
rect 1857 3887 1915 3893
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 2225 3927 2283 3933
rect 2225 3924 2237 3927
rect 2004 3896 2237 3924
rect 2004 3884 2010 3896
rect 2225 3893 2237 3896
rect 2271 3893 2283 3927
rect 2225 3887 2283 3893
rect 3881 3927 3939 3933
rect 3881 3893 3893 3927
rect 3927 3924 3939 3927
rect 4246 3924 4252 3936
rect 3927 3896 4252 3924
rect 3927 3893 3939 3896
rect 3881 3887 3939 3893
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 4709 3927 4767 3933
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 5718 3924 5724 3936
rect 4755 3896 5724 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6181 3927 6239 3933
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 7006 3924 7012 3936
rect 6227 3896 7012 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 7300 3924 7328 4032
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8386 4060 8392 4072
rect 8343 4032 8392 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 13464 4060 13492 4100
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 14093 4131 14151 4137
rect 14093 4128 14105 4131
rect 13587 4100 14105 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 14093 4097 14105 4100
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 14182 4088 14188 4140
rect 14240 4128 14246 4140
rect 14349 4131 14407 4137
rect 14349 4128 14361 4131
rect 14240 4100 14361 4128
rect 14240 4088 14246 4100
rect 14349 4097 14361 4100
rect 14395 4097 14407 4131
rect 14349 4091 14407 4097
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 16408 4137 16436 4168
rect 16393 4131 16451 4137
rect 16393 4128 16405 4131
rect 16356 4100 16405 4128
rect 16356 4088 16362 4100
rect 16393 4097 16405 4100
rect 16439 4097 16451 4131
rect 16393 4091 16451 4097
rect 16761 4131 16819 4137
rect 16761 4097 16773 4131
rect 16807 4128 16819 4131
rect 17494 4128 17500 4140
rect 16807 4100 17500 4128
rect 16807 4097 16819 4100
rect 16761 4091 16819 4097
rect 17494 4088 17500 4100
rect 17552 4088 17558 4140
rect 17604 4128 17632 4168
rect 17954 4128 17960 4140
rect 17604 4100 17960 4128
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 18417 4131 18475 4137
rect 18417 4097 18429 4131
rect 18463 4128 18475 4131
rect 19334 4128 19340 4140
rect 18463 4100 19340 4128
rect 18463 4097 18475 4100
rect 18417 4091 18475 4097
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 13817 4063 13875 4069
rect 13817 4060 13829 4063
rect 13464 4032 13829 4060
rect 13817 4029 13829 4032
rect 13863 4029 13875 4063
rect 13817 4023 13875 4029
rect 15470 4020 15476 4072
rect 15528 4060 15534 4072
rect 16117 4063 16175 4069
rect 16117 4060 16129 4063
rect 15528 4032 16129 4060
rect 15528 4020 15534 4032
rect 16117 4029 16129 4032
rect 16163 4029 16175 4063
rect 17310 4060 17316 4072
rect 16117 4023 16175 4029
rect 16224 4032 17316 4060
rect 11238 3992 11244 4004
rect 8312 3964 8892 3992
rect 11199 3964 11244 3992
rect 8312 3924 8340 3964
rect 7300 3896 8340 3924
rect 8864 3924 8892 3964
rect 11238 3952 11244 3964
rect 11296 3992 11302 4004
rect 12526 3992 12532 4004
rect 11296 3964 12532 3992
rect 11296 3952 11302 3964
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 16224 3992 16252 4032
rect 17310 4020 17316 4032
rect 17368 4020 17374 4072
rect 17402 4020 17408 4072
rect 17460 4060 17466 4072
rect 17589 4063 17647 4069
rect 17589 4060 17601 4063
rect 17460 4032 17601 4060
rect 17460 4020 17466 4032
rect 17589 4029 17601 4032
rect 17635 4029 17647 4063
rect 17589 4023 17647 4029
rect 17681 4063 17739 4069
rect 17681 4029 17693 4063
rect 17727 4029 17739 4063
rect 17681 4023 17739 4029
rect 15488 3964 16252 3992
rect 10226 3924 10232 3936
rect 8864 3896 10232 3924
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 10836 3896 12173 3924
rect 10836 3884 10842 3896
rect 12161 3893 12173 3896
rect 12207 3893 12219 3927
rect 12161 3887 12219 3893
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15488 3933 15516 3964
rect 16298 3952 16304 4004
rect 16356 3992 16362 4004
rect 16945 3995 17003 4001
rect 16945 3992 16957 3995
rect 16356 3964 16957 3992
rect 16356 3952 16362 3964
rect 16945 3961 16957 3964
rect 16991 3961 17003 3995
rect 17328 3992 17356 4020
rect 17696 3992 17724 4023
rect 17770 4020 17776 4072
rect 17828 4060 17834 4072
rect 19058 4060 19064 4072
rect 17828 4032 19064 4060
rect 17828 4020 17834 4032
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 17328 3964 17724 3992
rect 16945 3955 17003 3961
rect 15473 3927 15531 3933
rect 15473 3924 15485 3927
rect 15160 3896 15485 3924
rect 15160 3884 15166 3896
rect 15473 3893 15485 3896
rect 15519 3893 15531 3927
rect 15473 3887 15531 3893
rect 15565 3927 15623 3933
rect 15565 3893 15577 3927
rect 15611 3924 15623 3927
rect 15746 3924 15752 3936
rect 15611 3896 15752 3924
rect 15611 3893 15623 3896
rect 15565 3887 15623 3893
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 1104 3834 18860 3856
rect 1104 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 3430 3834
rect 3482 3782 7622 3834
rect 7674 3782 7686 3834
rect 7738 3782 7750 3834
rect 7802 3782 7814 3834
rect 7866 3782 7878 3834
rect 7930 3782 12070 3834
rect 12122 3782 12134 3834
rect 12186 3782 12198 3834
rect 12250 3782 12262 3834
rect 12314 3782 12326 3834
rect 12378 3782 16518 3834
rect 16570 3782 16582 3834
rect 16634 3782 16646 3834
rect 16698 3782 16710 3834
rect 16762 3782 16774 3834
rect 16826 3782 18860 3834
rect 1104 3760 18860 3782
rect 1489 3723 1547 3729
rect 1489 3689 1501 3723
rect 1535 3720 1547 3723
rect 1578 3720 1584 3732
rect 1535 3692 1584 3720
rect 1535 3689 1547 3692
rect 1489 3683 1547 3689
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 1673 3723 1731 3729
rect 1673 3689 1685 3723
rect 1719 3720 1731 3723
rect 2314 3720 2320 3732
rect 1719 3692 2320 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 3881 3723 3939 3729
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 4798 3720 4804 3732
rect 3927 3692 4804 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4798 3680 4804 3692
rect 4856 3720 4862 3732
rect 4985 3723 5043 3729
rect 4985 3720 4997 3723
rect 4856 3692 4997 3720
rect 4856 3680 4862 3692
rect 4985 3689 4997 3692
rect 5031 3689 5043 3723
rect 6362 3720 6368 3732
rect 4985 3683 5043 3689
rect 5460 3692 6368 3720
rect 1210 3612 1216 3664
rect 1268 3652 1274 3664
rect 1765 3655 1823 3661
rect 1765 3652 1777 3655
rect 1268 3624 1777 3652
rect 1268 3612 1274 3624
rect 1765 3621 1777 3624
rect 1811 3621 1823 3655
rect 1765 3615 1823 3621
rect 2041 3655 2099 3661
rect 2041 3621 2053 3655
rect 2087 3652 2099 3655
rect 2498 3652 2504 3664
rect 2087 3624 2504 3652
rect 2087 3621 2099 3624
rect 2041 3615 2099 3621
rect 1780 3516 1808 3615
rect 2498 3612 2504 3624
rect 2556 3612 2562 3664
rect 2590 3612 2596 3664
rect 2648 3652 2654 3664
rect 2869 3655 2927 3661
rect 2869 3652 2881 3655
rect 2648 3624 2881 3652
rect 2648 3612 2654 3624
rect 2869 3621 2881 3624
rect 2915 3621 2927 3655
rect 2869 3615 2927 3621
rect 2958 3612 2964 3664
rect 3016 3652 3022 3664
rect 3973 3655 4031 3661
rect 3973 3652 3985 3655
rect 3016 3624 3985 3652
rect 3016 3612 3022 3624
rect 3973 3621 3985 3624
rect 4019 3621 4031 3655
rect 3973 3615 4031 3621
rect 4706 3612 4712 3664
rect 4764 3652 4770 3664
rect 5169 3655 5227 3661
rect 5169 3652 5181 3655
rect 4764 3624 5181 3652
rect 4764 3612 4770 3624
rect 5169 3621 5181 3624
rect 5215 3621 5227 3655
rect 5169 3615 5227 3621
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3584 2283 3587
rect 2406 3584 2412 3596
rect 2271 3556 2412 3584
rect 2271 3553 2283 3556
rect 2225 3547 2283 3553
rect 2406 3544 2412 3556
rect 2464 3584 2470 3596
rect 2464 3556 3004 3584
rect 2464 3544 2470 3556
rect 1780 3488 2728 3516
rect 2038 3408 2044 3460
rect 2096 3448 2102 3460
rect 2501 3451 2559 3457
rect 2501 3448 2513 3451
rect 2096 3420 2513 3448
rect 2096 3408 2102 3420
rect 2501 3417 2513 3420
rect 2547 3417 2559 3451
rect 2700 3448 2728 3488
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 2832 3488 2877 3516
rect 2832 3476 2838 3488
rect 2976 3448 3004 3556
rect 3050 3544 3056 3596
rect 3108 3584 3114 3596
rect 3329 3587 3387 3593
rect 3329 3584 3341 3587
rect 3108 3556 3341 3584
rect 3108 3544 3114 3556
rect 3329 3553 3341 3556
rect 3375 3553 3387 3587
rect 3329 3547 3387 3553
rect 3421 3587 3479 3593
rect 3421 3553 3433 3587
rect 3467 3584 3479 3587
rect 3467 3556 4476 3584
rect 3467 3553 3479 3556
rect 3421 3547 3479 3553
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3510 3516 3516 3528
rect 3283 3488 3516 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 4448 3516 4476 3556
rect 4522 3544 4528 3596
rect 4580 3584 4586 3596
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 4580 3556 4629 3584
rect 4580 3544 4586 3556
rect 4617 3553 4629 3556
rect 4663 3584 4675 3587
rect 5460 3584 5488 3692
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 11146 3720 11152 3732
rect 7024 3692 11152 3720
rect 7024 3584 7052 3692
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 11422 3680 11428 3732
rect 11480 3720 11486 3732
rect 11885 3723 11943 3729
rect 11885 3720 11897 3723
rect 11480 3692 11897 3720
rect 11480 3680 11486 3692
rect 11885 3689 11897 3692
rect 11931 3689 11943 3723
rect 13446 3720 13452 3732
rect 13407 3692 13452 3720
rect 11885 3683 11943 3689
rect 13446 3680 13452 3692
rect 13504 3720 13510 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 13504 3692 13645 3720
rect 13504 3680 13510 3692
rect 13633 3689 13645 3692
rect 13679 3720 13691 3723
rect 13817 3723 13875 3729
rect 13817 3720 13829 3723
rect 13679 3692 13829 3720
rect 13679 3689 13691 3692
rect 13633 3683 13691 3689
rect 13817 3689 13829 3692
rect 13863 3689 13875 3723
rect 13817 3683 13875 3689
rect 14093 3723 14151 3729
rect 14093 3689 14105 3723
rect 14139 3720 14151 3723
rect 15194 3720 15200 3732
rect 14139 3692 15200 3720
rect 14139 3689 14151 3692
rect 14093 3683 14151 3689
rect 15194 3680 15200 3692
rect 15252 3680 15258 3732
rect 15470 3680 15476 3732
rect 15528 3720 15534 3732
rect 15565 3723 15623 3729
rect 15565 3720 15577 3723
rect 15528 3692 15577 3720
rect 15528 3680 15534 3692
rect 15565 3689 15577 3692
rect 15611 3689 15623 3723
rect 15565 3683 15623 3689
rect 17218 3680 17224 3732
rect 17276 3720 17282 3732
rect 17497 3723 17555 3729
rect 17497 3720 17509 3723
rect 17276 3692 17509 3720
rect 17276 3680 17282 3692
rect 17497 3689 17509 3692
rect 17543 3689 17555 3723
rect 17497 3683 17555 3689
rect 18046 3680 18052 3732
rect 18104 3720 18110 3732
rect 18325 3723 18383 3729
rect 18325 3720 18337 3723
rect 18104 3692 18337 3720
rect 18104 3680 18110 3692
rect 18325 3689 18337 3692
rect 18371 3689 18383 3723
rect 18325 3683 18383 3689
rect 8018 3612 8024 3664
rect 8076 3652 8082 3664
rect 8076 3624 8791 3652
rect 8076 3612 8082 3624
rect 8386 3584 8392 3596
rect 4663 3556 5488 3584
rect 6472 3556 7052 3584
rect 8128 3556 8392 3584
rect 4663 3553 4675 3556
rect 4617 3547 4675 3553
rect 6472 3516 6500 3556
rect 4448 3488 6500 3516
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3516 6607 3519
rect 6638 3516 6644 3528
rect 6595 3488 6644 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 6638 3476 6644 3488
rect 6696 3516 6702 3528
rect 8128 3525 8156 3556
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 6696 3488 8033 3516
rect 6696 3476 6702 3488
rect 8021 3485 8033 3488
rect 8067 3516 8079 3519
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 8067 3488 8125 3516
rect 8067 3485 8079 3488
rect 8021 3479 8079 3485
rect 8113 3485 8125 3488
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3516 8355 3519
rect 8478 3516 8484 3528
rect 8343 3488 8484 3516
rect 8343 3485 8355 3488
rect 8297 3479 8355 3485
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 3050 3448 3056 3460
rect 2700 3420 2912 3448
rect 2976 3420 3056 3448
rect 2501 3411 2559 3417
rect 2884 3380 2912 3420
rect 3050 3408 3056 3420
rect 3108 3448 3114 3460
rect 4430 3448 4436 3460
rect 3108 3420 4436 3448
rect 3108 3408 3114 3420
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 4614 3408 4620 3460
rect 4672 3448 4678 3460
rect 6304 3451 6362 3457
rect 4672 3420 6224 3448
rect 4672 3408 4678 3420
rect 4341 3383 4399 3389
rect 4341 3380 4353 3383
rect 2884 3352 4353 3380
rect 4341 3349 4353 3352
rect 4387 3380 4399 3383
rect 4706 3380 4712 3392
rect 4387 3352 4712 3380
rect 4387 3349 4399 3352
rect 4341 3343 4399 3349
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 6196 3380 6224 3420
rect 6304 3417 6316 3451
rect 6350 3448 6362 3451
rect 6454 3448 6460 3460
rect 6350 3420 6460 3448
rect 6350 3417 6362 3420
rect 6304 3411 6362 3417
rect 6454 3408 6460 3420
rect 6512 3408 6518 3460
rect 7776 3451 7834 3457
rect 7776 3417 7788 3451
rect 7822 3448 7834 3451
rect 8202 3448 8208 3460
rect 7822 3420 8208 3448
rect 7822 3417 7834 3420
rect 7776 3411 7834 3417
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 8573 3451 8631 3457
rect 8573 3417 8585 3451
rect 8619 3448 8631 3451
rect 8662 3448 8668 3460
rect 8619 3420 8668 3448
rect 8619 3417 8631 3420
rect 8573 3411 8631 3417
rect 8662 3408 8668 3420
rect 8720 3408 8726 3460
rect 8763 3448 8791 3624
rect 8846 3612 8852 3664
rect 8904 3652 8910 3664
rect 9033 3655 9091 3661
rect 9033 3652 9045 3655
rect 8904 3624 9045 3652
rect 8904 3612 8910 3624
rect 9033 3621 9045 3624
rect 9079 3621 9091 3655
rect 9033 3615 9091 3621
rect 9048 3516 9076 3615
rect 13357 3587 13415 3593
rect 13357 3553 13369 3587
rect 13403 3584 13415 3587
rect 13464 3584 13492 3680
rect 13403 3556 13492 3584
rect 15473 3587 15531 3593
rect 13403 3553 13415 3556
rect 13357 3547 13415 3553
rect 15473 3553 15485 3587
rect 15519 3584 15531 3587
rect 15562 3584 15568 3596
rect 15519 3556 15568 3584
rect 15519 3553 15531 3556
rect 15473 3547 15531 3553
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 17862 3544 17868 3596
rect 17920 3584 17926 3596
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 17920 3556 18061 3584
rect 17920 3544 17926 3556
rect 18049 3553 18061 3556
rect 18095 3553 18107 3587
rect 18049 3547 18107 3553
rect 10413 3519 10471 3525
rect 9048 3488 10272 3516
rect 9950 3448 9956 3460
rect 8763 3420 9956 3448
rect 9950 3408 9956 3420
rect 10008 3408 10014 3460
rect 10134 3448 10140 3460
rect 10192 3457 10198 3460
rect 10104 3420 10140 3448
rect 10134 3408 10140 3420
rect 10192 3411 10204 3457
rect 10244 3448 10272 3488
rect 10413 3485 10425 3519
rect 10459 3516 10471 3519
rect 10505 3519 10563 3525
rect 10505 3516 10517 3519
rect 10459 3488 10517 3516
rect 10459 3485 10471 3488
rect 10413 3479 10471 3485
rect 10505 3485 10517 3488
rect 10551 3516 10563 3519
rect 11606 3516 11612 3528
rect 10551 3488 11612 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 11698 3476 11704 3528
rect 11756 3516 11762 3528
rect 13101 3519 13159 3525
rect 11756 3488 12434 3516
rect 11756 3476 11762 3488
rect 10750 3451 10808 3457
rect 10750 3448 10762 3451
rect 10244 3420 10762 3448
rect 10750 3417 10762 3420
rect 10796 3417 10808 3451
rect 10750 3411 10808 3417
rect 10192 3408 10198 3411
rect 10870 3408 10876 3460
rect 10928 3448 10934 3460
rect 10928 3420 12020 3448
rect 10928 3408 10934 3420
rect 6641 3383 6699 3389
rect 6641 3380 6653 3383
rect 6196 3352 6653 3380
rect 6641 3349 6653 3352
rect 6687 3380 6699 3383
rect 8754 3380 8760 3392
rect 6687 3352 8760 3380
rect 6687 3349 6699 3352
rect 6641 3343 6699 3349
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 10502 3380 10508 3392
rect 9732 3352 10508 3380
rect 9732 3340 9738 3352
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 11992 3389 12020 3420
rect 11977 3383 12035 3389
rect 11977 3349 11989 3383
rect 12023 3349 12035 3383
rect 12406 3380 12434 3488
rect 13101 3485 13113 3519
rect 13147 3516 13159 3519
rect 13538 3516 13544 3528
rect 13147 3488 13544 3516
rect 13147 3485 13159 3488
rect 13101 3479 13159 3485
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 15580 3516 15608 3544
rect 15838 3516 15844 3528
rect 15580 3488 15844 3516
rect 15838 3476 15844 3488
rect 15896 3516 15902 3528
rect 16945 3519 17003 3525
rect 16945 3516 16957 3519
rect 15896 3488 16957 3516
rect 15896 3476 15902 3488
rect 16945 3485 16957 3488
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 17129 3519 17187 3525
rect 17129 3485 17141 3519
rect 17175 3516 17187 3519
rect 17218 3516 17224 3528
rect 17175 3488 17224 3516
rect 17175 3485 17187 3488
rect 17129 3479 17187 3485
rect 17218 3476 17224 3488
rect 17276 3516 17282 3528
rect 17678 3516 17684 3528
rect 17276 3488 17684 3516
rect 17276 3476 17282 3488
rect 17678 3476 17684 3488
rect 17736 3476 17742 3528
rect 17954 3516 17960 3528
rect 17880 3488 17960 3516
rect 15228 3451 15286 3457
rect 15228 3417 15240 3451
rect 15274 3448 15286 3451
rect 15654 3448 15660 3460
rect 15274 3420 15660 3448
rect 15274 3417 15286 3420
rect 15228 3411 15286 3417
rect 15654 3408 15660 3420
rect 15712 3408 15718 3460
rect 16700 3451 16758 3457
rect 16700 3417 16712 3451
rect 16746 3448 16758 3451
rect 17034 3448 17040 3460
rect 16746 3420 17040 3448
rect 16746 3417 16758 3420
rect 16700 3411 16758 3417
rect 17034 3408 17040 3420
rect 17092 3408 17098 3460
rect 17880 3457 17908 3488
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 17865 3451 17923 3457
rect 17865 3417 17877 3451
rect 17911 3417 17923 3451
rect 17865 3411 17923 3417
rect 16574 3380 16580 3392
rect 12406 3352 16580 3380
rect 11977 3343 12035 3349
rect 16574 3340 16580 3352
rect 16632 3340 16638 3392
rect 17313 3383 17371 3389
rect 17313 3349 17325 3383
rect 17359 3380 17371 3383
rect 17402 3380 17408 3392
rect 17359 3352 17408 3380
rect 17359 3349 17371 3352
rect 17313 3343 17371 3349
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 17586 3340 17592 3392
rect 17644 3380 17650 3392
rect 17957 3383 18015 3389
rect 17957 3380 17969 3383
rect 17644 3352 17969 3380
rect 17644 3340 17650 3352
rect 17957 3349 17969 3352
rect 18003 3349 18015 3383
rect 17957 3343 18015 3349
rect 1104 3290 18860 3312
rect 1104 3238 5398 3290
rect 5450 3238 5462 3290
rect 5514 3238 5526 3290
rect 5578 3238 5590 3290
rect 5642 3238 5654 3290
rect 5706 3238 9846 3290
rect 9898 3238 9910 3290
rect 9962 3238 9974 3290
rect 10026 3238 10038 3290
rect 10090 3238 10102 3290
rect 10154 3238 14294 3290
rect 14346 3238 14358 3290
rect 14410 3238 14422 3290
rect 14474 3238 14486 3290
rect 14538 3238 14550 3290
rect 14602 3238 18860 3290
rect 1104 3216 18860 3238
rect 3694 3176 3700 3188
rect 2792 3148 3700 3176
rect 2406 3108 2412 3120
rect 1688 3080 2412 3108
rect 1688 3049 1716 3080
rect 2406 3068 2412 3080
rect 2464 3068 2470 3120
rect 2590 3068 2596 3120
rect 2648 3068 2654 3120
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2608 3040 2636 3068
rect 2792 3049 2820 3148
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 4246 3176 4252 3188
rect 4207 3148 4252 3176
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4338 3136 4344 3188
rect 4396 3176 4402 3188
rect 4709 3179 4767 3185
rect 4396 3148 4441 3176
rect 4396 3136 4402 3148
rect 4709 3145 4721 3179
rect 4755 3176 4767 3179
rect 5626 3176 5632 3188
rect 4755 3148 5632 3176
rect 4755 3145 4767 3148
rect 4709 3139 4767 3145
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 5736 3148 7880 3176
rect 3053 3111 3111 3117
rect 3053 3077 3065 3111
rect 3099 3108 3111 3111
rect 5258 3108 5264 3120
rect 3099 3080 5264 3108
rect 3099 3077 3111 3080
rect 3053 3071 3111 3077
rect 5258 3068 5264 3080
rect 5316 3068 5322 3120
rect 2271 3012 2636 3040
rect 2777 3043 2835 3049
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 3326 3040 3332 3052
rect 3287 3012 3332 3040
rect 2777 3003 2835 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3602 3000 3608 3052
rect 3660 3040 3666 3052
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3660 3012 3893 3040
rect 3660 3000 3666 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 5736 3040 5764 3148
rect 6638 3068 6644 3120
rect 6696 3108 6702 3120
rect 7852 3108 7880 3148
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8168 3148 9076 3176
rect 8168 3136 8174 3148
rect 8570 3108 8576 3120
rect 6696 3080 7788 3108
rect 7852 3080 8576 3108
rect 6696 3068 6702 3080
rect 3881 3003 3939 3009
rect 3988 3012 4660 3040
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2941 2099 2975
rect 2041 2935 2099 2941
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2972 2651 2975
rect 3697 2975 3755 2981
rect 2639 2944 3096 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 2056 2904 2084 2935
rect 2866 2904 2872 2916
rect 2056 2876 2872 2904
rect 2866 2864 2872 2876
rect 2924 2864 2930 2916
rect 3068 2904 3096 2944
rect 3697 2941 3709 2975
rect 3743 2972 3755 2975
rect 3988 2972 4016 3012
rect 4154 2972 4160 2984
rect 3743 2944 4016 2972
rect 4115 2944 4160 2972
rect 3743 2941 3755 2944
rect 3697 2935 3755 2941
rect 4154 2932 4160 2944
rect 4212 2932 4218 2984
rect 4522 2904 4528 2916
rect 3068 2876 4528 2904
rect 4522 2864 4528 2876
rect 4580 2864 4586 2916
rect 1486 2836 1492 2848
rect 1447 2808 1492 2836
rect 1486 2796 1492 2808
rect 1544 2796 1550 2848
rect 4632 2836 4660 3012
rect 5184 3012 5764 3040
rect 5914 3043 5972 3049
rect 4801 2907 4859 2913
rect 4801 2873 4813 2907
rect 4847 2904 4859 2907
rect 4890 2904 4896 2916
rect 4847 2876 4896 2904
rect 4847 2873 4859 2876
rect 4801 2867 4859 2873
rect 4890 2864 4896 2876
rect 4948 2904 4954 2916
rect 5184 2904 5212 3012
rect 5914 3009 5926 3043
rect 5960 3040 5972 3043
rect 6086 3040 6092 3052
rect 5960 3012 6092 3040
rect 5960 3009 5972 3012
rect 5914 3003 5972 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7760 3049 7788 3080
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 8754 3117 8760 3120
rect 8748 3108 8760 3117
rect 8715 3080 8760 3108
rect 8748 3071 8760 3080
rect 8754 3068 8760 3071
rect 8812 3068 8818 3120
rect 9048 3108 9076 3148
rect 9214 3136 9220 3188
rect 9272 3176 9278 3188
rect 9861 3179 9919 3185
rect 9861 3176 9873 3179
rect 9272 3148 9873 3176
rect 9272 3136 9278 3148
rect 9861 3145 9873 3148
rect 9907 3176 9919 3179
rect 10318 3176 10324 3188
rect 9907 3148 10324 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 11517 3179 11575 3185
rect 11517 3176 11529 3179
rect 10428 3148 11529 3176
rect 9048 3080 9536 3108
rect 7478 3043 7536 3049
rect 7478 3040 7490 3043
rect 6972 3012 7490 3040
rect 6972 3000 6978 3012
rect 7478 3009 7490 3012
rect 7524 3040 7536 3043
rect 7745 3043 7803 3049
rect 7524 3012 7696 3040
rect 7524 3009 7536 3012
rect 7478 3003 7536 3009
rect 6178 2932 6184 2984
rect 6236 2972 6242 2984
rect 6638 2972 6644 2984
rect 6236 2944 6644 2972
rect 6236 2932 6242 2944
rect 6638 2932 6644 2944
rect 6696 2932 6702 2984
rect 7668 2972 7696 3012
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3040 8447 3043
rect 9030 3040 9036 3052
rect 8435 3012 9036 3040
rect 8435 3009 8447 3012
rect 8389 3003 8447 3009
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 9508 3040 9536 3080
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 10428 3108 10456 3148
rect 11517 3145 11529 3148
rect 11563 3145 11575 3179
rect 14458 3176 14464 3188
rect 11517 3139 11575 3145
rect 13657 3148 14136 3176
rect 14419 3148 14464 3176
rect 9640 3080 10456 3108
rect 9640 3068 9646 3080
rect 10502 3068 10508 3120
rect 10560 3108 10566 3120
rect 11606 3108 11612 3120
rect 10560 3080 11284 3108
rect 10560 3068 10566 3080
rect 10778 3040 10784 3052
rect 9508 3012 10784 3040
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11054 3000 11060 3052
rect 11112 3049 11118 3052
rect 11112 3040 11124 3049
rect 11112 3012 11157 3040
rect 11112 3003 11124 3012
rect 11112 3000 11118 3003
rect 8110 2972 8116 2984
rect 7668 2944 8116 2972
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 8205 2975 8263 2981
rect 8205 2941 8217 2975
rect 8251 2941 8263 2975
rect 8478 2972 8484 2984
rect 8439 2944 8484 2972
rect 8205 2935 8263 2941
rect 6730 2904 6736 2916
rect 4948 2876 5212 2904
rect 6288 2876 6736 2904
rect 4948 2864 4954 2876
rect 6288 2836 6316 2876
rect 6730 2864 6736 2876
rect 6788 2864 6794 2916
rect 4632 2808 6316 2836
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 8018 2836 8024 2848
rect 6420 2808 8024 2836
rect 6420 2796 6426 2808
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 8220 2836 8248 2935
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 11256 2972 11284 3080
rect 11348 3080 11612 3108
rect 11348 3049 11376 3080
rect 11606 3068 11612 3080
rect 11664 3068 11670 3120
rect 13446 3108 13452 3120
rect 13004 3080 13452 3108
rect 13004 3049 13032 3080
rect 13446 3068 13452 3080
rect 13504 3068 13510 3120
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3009 11391 3043
rect 12630 3043 12688 3049
rect 12630 3040 12642 3043
rect 11333 3003 11391 3009
rect 11440 3012 12642 3040
rect 11440 2972 11468 3012
rect 12630 3009 12642 3012
rect 12676 3009 12688 3043
rect 12630 3003 12688 3009
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3040 12955 3043
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12943 3012 13001 3040
rect 12943 3009 12955 3012
rect 12897 3003 12955 3009
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 13078 3000 13084 3052
rect 13136 3040 13142 3052
rect 13256 3043 13314 3049
rect 13256 3040 13268 3043
rect 13136 3012 13268 3040
rect 13136 3000 13142 3012
rect 13256 3009 13268 3012
rect 13302 3040 13314 3043
rect 13657 3040 13685 3148
rect 14108 3108 14136 3148
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 14568 3148 16344 3176
rect 14568 3108 14596 3148
rect 14108 3080 14596 3108
rect 15562 3068 15568 3120
rect 15620 3117 15626 3120
rect 15620 3108 15632 3117
rect 16316 3108 16344 3148
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 16945 3179 17003 3185
rect 16945 3176 16957 3179
rect 16908 3148 16957 3176
rect 16908 3136 16914 3148
rect 16945 3145 16957 3148
rect 16991 3145 17003 3179
rect 16945 3139 17003 3145
rect 17405 3179 17463 3185
rect 17405 3145 17417 3179
rect 17451 3176 17463 3179
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 17451 3148 17785 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 17773 3145 17785 3148
rect 17819 3145 17831 3179
rect 17773 3139 17831 3145
rect 18141 3179 18199 3185
rect 18141 3145 18153 3179
rect 18187 3176 18199 3179
rect 18322 3176 18328 3188
rect 18187 3148 18328 3176
rect 18187 3145 18199 3148
rect 18141 3139 18199 3145
rect 18322 3136 18328 3148
rect 18380 3136 18386 3188
rect 15620 3080 15665 3108
rect 16316 3080 18368 3108
rect 15620 3071 15632 3080
rect 15620 3068 15626 3071
rect 15838 3040 15844 3052
rect 13302 3012 13685 3040
rect 15799 3012 15844 3040
rect 13302 3009 13314 3012
rect 13256 3003 13314 3009
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 15930 3000 15936 3052
rect 15988 3040 15994 3052
rect 15988 3012 16033 3040
rect 15988 3000 15994 3012
rect 16574 3000 16580 3052
rect 16632 3040 16638 3052
rect 17034 3040 17040 3052
rect 16632 3012 17040 3040
rect 16632 3000 16638 3012
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 17313 3043 17371 3049
rect 17313 3040 17325 3043
rect 17184 3012 17325 3040
rect 17184 3000 17190 3012
rect 17313 3009 17325 3012
rect 17359 3009 17371 3043
rect 17313 3003 17371 3009
rect 11256 2944 11468 2972
rect 16022 2932 16028 2984
rect 16080 2972 16086 2984
rect 16117 2975 16175 2981
rect 16117 2972 16129 2975
rect 16080 2944 16129 2972
rect 16080 2932 16086 2944
rect 16117 2941 16129 2944
rect 16163 2941 16175 2975
rect 16117 2935 16175 2941
rect 17589 2975 17647 2981
rect 17589 2941 17601 2975
rect 17635 2972 17647 2975
rect 17862 2972 17868 2984
rect 17635 2944 17868 2972
rect 17635 2941 17647 2944
rect 17589 2935 17647 2941
rect 17862 2932 17868 2944
rect 17920 2932 17926 2984
rect 18340 2981 18368 3080
rect 18233 2975 18291 2981
rect 18233 2941 18245 2975
rect 18279 2941 18291 2975
rect 18233 2935 18291 2941
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2941 18383 2975
rect 18325 2935 18383 2941
rect 9876 2876 10456 2904
rect 9876 2836 9904 2876
rect 8220 2808 9904 2836
rect 9953 2839 10011 2845
rect 9953 2805 9965 2839
rect 9999 2836 10011 2839
rect 10318 2836 10324 2848
rect 9999 2808 10324 2836
rect 9999 2805 10011 2808
rect 9953 2799 10011 2805
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 10428 2836 10456 2876
rect 14090 2864 14096 2916
rect 14148 2904 14154 2916
rect 14366 2904 14372 2916
rect 14148 2876 14372 2904
rect 14148 2864 14154 2876
rect 14366 2864 14372 2876
rect 14424 2864 14430 2916
rect 16850 2904 16856 2916
rect 16763 2876 16856 2904
rect 16850 2864 16856 2876
rect 16908 2904 16914 2916
rect 17494 2904 17500 2916
rect 16908 2876 17500 2904
rect 16908 2864 16914 2876
rect 17494 2864 17500 2876
rect 17552 2904 17558 2916
rect 18248 2904 18276 2935
rect 17552 2876 18276 2904
rect 17552 2864 17558 2876
rect 11146 2836 11152 2848
rect 10428 2808 11152 2836
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 12894 2796 12900 2848
rect 12952 2836 12958 2848
rect 15470 2836 15476 2848
rect 12952 2808 15476 2836
rect 12952 2796 12958 2808
rect 15470 2796 15476 2808
rect 15528 2796 15534 2848
rect 17034 2796 17040 2848
rect 17092 2836 17098 2848
rect 17310 2836 17316 2848
rect 17092 2808 17316 2836
rect 17092 2796 17098 2808
rect 17310 2796 17316 2808
rect 17368 2836 17374 2848
rect 18138 2836 18144 2848
rect 17368 2808 18144 2836
rect 17368 2796 17374 2808
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 1104 2746 18860 2768
rect 1104 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 3430 2746
rect 3482 2694 7622 2746
rect 7674 2694 7686 2746
rect 7738 2694 7750 2746
rect 7802 2694 7814 2746
rect 7866 2694 7878 2746
rect 7930 2694 12070 2746
rect 12122 2694 12134 2746
rect 12186 2694 12198 2746
rect 12250 2694 12262 2746
rect 12314 2694 12326 2746
rect 12378 2694 16518 2746
rect 16570 2694 16582 2746
rect 16634 2694 16646 2746
rect 16698 2694 16710 2746
rect 16762 2694 16774 2746
rect 16826 2694 18860 2746
rect 1104 2672 18860 2694
rect 1302 2592 1308 2644
rect 1360 2632 1366 2644
rect 1489 2635 1547 2641
rect 1489 2632 1501 2635
rect 1360 2604 1501 2632
rect 1360 2592 1366 2604
rect 1489 2601 1501 2604
rect 1535 2601 1547 2635
rect 2682 2632 2688 2644
rect 2643 2604 2688 2632
rect 1489 2595 1547 2601
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 3050 2632 3056 2644
rect 3011 2604 3056 2632
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 5994 2632 6000 2644
rect 4080 2604 6000 2632
rect 1210 2524 1216 2576
rect 1268 2564 1274 2576
rect 2317 2567 2375 2573
rect 2317 2564 2329 2567
rect 1268 2536 2329 2564
rect 1268 2524 1274 2536
rect 2317 2533 2329 2536
rect 2363 2533 2375 2567
rect 2317 2527 2375 2533
rect 2869 2567 2927 2573
rect 2869 2533 2881 2567
rect 2915 2564 2927 2567
rect 2915 2536 4016 2564
rect 2915 2533 2927 2536
rect 2869 2527 2927 2533
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 2774 2496 2780 2508
rect 1995 2468 2780 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 3878 2496 3884 2508
rect 3620 2468 3884 2496
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2397 2191 2431
rect 2498 2428 2504 2440
rect 2459 2400 2504 2428
rect 2133 2391 2191 2397
rect 2148 2360 2176 2391
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 3620 2437 3648 2468
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2397 3663 2431
rect 3786 2428 3792 2440
rect 3747 2400 3792 2428
rect 3605 2391 3663 2397
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 3988 2428 4016 2536
rect 4080 2505 4108 2604
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 6178 2632 6184 2644
rect 6139 2604 6184 2632
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 7009 2635 7067 2641
rect 7009 2601 7021 2635
rect 7055 2632 7067 2635
rect 7466 2632 7472 2644
rect 7055 2604 7472 2632
rect 7055 2601 7067 2604
rect 7009 2595 7067 2601
rect 5077 2567 5135 2573
rect 5077 2533 5089 2567
rect 5123 2533 5135 2567
rect 7024 2564 7052 2595
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 8478 2632 8484 2644
rect 8439 2604 8484 2632
rect 8478 2592 8484 2604
rect 8536 2632 8542 2644
rect 8665 2635 8723 2641
rect 8665 2632 8677 2635
rect 8536 2604 8677 2632
rect 8536 2592 8542 2604
rect 8665 2601 8677 2604
rect 8711 2632 8723 2635
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8711 2604 8953 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 9398 2632 9404 2644
rect 9355 2604 9404 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 11606 2632 11612 2644
rect 11567 2604 11612 2632
rect 11606 2592 11612 2604
rect 11664 2632 11670 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 11664 2604 11713 2632
rect 11664 2592 11670 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 11701 2595 11759 2601
rect 14737 2635 14795 2641
rect 14737 2601 14749 2635
rect 14783 2632 14795 2635
rect 14829 2635 14887 2641
rect 14829 2632 14841 2635
rect 14783 2604 14841 2632
rect 14783 2601 14795 2604
rect 14737 2595 14795 2601
rect 14829 2601 14841 2604
rect 14875 2632 14887 2635
rect 15013 2635 15071 2641
rect 15013 2632 15025 2635
rect 14875 2604 15025 2632
rect 14875 2601 14887 2604
rect 14829 2595 14887 2601
rect 15013 2601 15025 2604
rect 15059 2632 15071 2635
rect 15838 2632 15844 2644
rect 15059 2604 15844 2632
rect 15059 2601 15071 2604
rect 15013 2595 15071 2601
rect 5077 2527 5135 2533
rect 5368 2536 7052 2564
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4154 2456 4160 2508
rect 4212 2496 4218 2508
rect 4525 2499 4583 2505
rect 4525 2496 4537 2499
rect 4212 2468 4537 2496
rect 4212 2456 4218 2468
rect 4525 2465 4537 2468
rect 4571 2496 4583 2499
rect 4798 2496 4804 2508
rect 4571 2468 4804 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 4338 2428 4344 2440
rect 3988 2400 4344 2428
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4430 2388 4436 2440
rect 4488 2428 4494 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4488 2400 4629 2428
rect 4488 2388 4494 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 5092 2428 5120 2527
rect 5368 2505 5396 2536
rect 5353 2499 5411 2505
rect 5353 2465 5365 2499
rect 5399 2465 5411 2499
rect 5353 2459 5411 2465
rect 5445 2499 5503 2505
rect 5445 2465 5457 2499
rect 5491 2496 5503 2499
rect 5626 2496 5632 2508
rect 5491 2468 5632 2496
rect 5491 2465 5503 2468
rect 5445 2459 5503 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 8389 2499 8447 2505
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 8496 2496 8524 2592
rect 8435 2468 8524 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 9861 2499 9919 2505
rect 9861 2496 9873 2499
rect 9732 2468 9873 2496
rect 9732 2456 9738 2468
rect 9861 2465 9873 2468
rect 9907 2465 9919 2499
rect 9861 2459 9919 2465
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2496 10287 2499
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 10275 2468 11161 2496
rect 10275 2465 10287 2468
rect 10229 2459 10287 2465
rect 11149 2465 11161 2468
rect 11195 2496 11207 2499
rect 11624 2496 11652 2592
rect 11195 2468 11652 2496
rect 13909 2499 13967 2505
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 13909 2465 13921 2499
rect 13955 2496 13967 2499
rect 14752 2496 14780 2595
rect 15838 2592 15844 2604
rect 15896 2592 15902 2644
rect 16117 2635 16175 2641
rect 16117 2601 16129 2635
rect 16163 2632 16175 2635
rect 17037 2635 17095 2641
rect 16163 2604 16988 2632
rect 16163 2601 16175 2604
rect 16117 2595 16175 2601
rect 16301 2567 16359 2573
rect 16301 2533 16313 2567
rect 16347 2564 16359 2567
rect 16666 2564 16672 2576
rect 16347 2536 16672 2564
rect 16347 2533 16359 2536
rect 16301 2527 16359 2533
rect 16666 2524 16672 2536
rect 16724 2524 16730 2576
rect 16761 2567 16819 2573
rect 16761 2533 16773 2567
rect 16807 2564 16819 2567
rect 16850 2564 16856 2576
rect 16807 2536 16856 2564
rect 16807 2533 16819 2536
rect 16761 2527 16819 2533
rect 16850 2524 16856 2536
rect 16908 2524 16914 2576
rect 16960 2564 16988 2604
rect 17037 2601 17049 2635
rect 17083 2632 17095 2635
rect 17126 2632 17132 2644
rect 17083 2604 17132 2632
rect 17083 2601 17095 2604
rect 17037 2595 17095 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 17218 2564 17224 2576
rect 16960 2536 17224 2564
rect 17218 2524 17224 2536
rect 17276 2524 17282 2576
rect 18598 2496 18604 2508
rect 13955 2468 14780 2496
rect 14844 2468 18604 2496
rect 13955 2465 13967 2468
rect 13909 2459 13967 2465
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 4764 2400 4809 2428
rect 5092 2400 5549 2428
rect 4764 2388 4770 2400
rect 5537 2397 5549 2400
rect 5583 2397 5595 2431
rect 6454 2428 6460 2440
rect 6415 2400 6460 2428
rect 5537 2391 5595 2397
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 8294 2428 8300 2440
rect 6656 2400 8300 2428
rect 3329 2363 3387 2369
rect 2148 2332 3280 2360
rect 3252 2292 3280 2332
rect 3329 2329 3341 2363
rect 3375 2360 3387 2363
rect 3694 2360 3700 2372
rect 3375 2332 3700 2360
rect 3375 2329 3387 2332
rect 3329 2323 3387 2329
rect 3694 2320 3700 2332
rect 3752 2320 3758 2372
rect 6656 2360 6684 2400
rect 8294 2388 8300 2400
rect 8352 2428 8358 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8352 2400 9137 2428
rect 8352 2388 8358 2400
rect 9125 2397 9137 2400
rect 9171 2428 9183 2431
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 9171 2400 10333 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 10321 2397 10333 2400
rect 10367 2428 10379 2431
rect 12342 2428 12348 2440
rect 10367 2400 12204 2428
rect 12303 2400 12348 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 4540 2332 6684 2360
rect 6733 2363 6791 2369
rect 4540 2292 4568 2332
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 7834 2360 7840 2372
rect 6779 2332 7840 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 7834 2320 7840 2332
rect 7892 2320 7898 2372
rect 7926 2320 7932 2372
rect 7984 2360 7990 2372
rect 8144 2363 8202 2369
rect 8144 2360 8156 2363
rect 7984 2332 8156 2360
rect 7984 2320 7990 2332
rect 8144 2329 8156 2332
rect 8190 2360 8202 2363
rect 9214 2360 9220 2372
rect 8190 2332 9220 2360
rect 8190 2329 8202 2332
rect 8144 2323 8202 2329
rect 9214 2320 9220 2332
rect 9272 2320 9278 2372
rect 9674 2360 9680 2372
rect 9635 2332 9680 2360
rect 9674 2320 9680 2332
rect 9732 2320 9738 2372
rect 11974 2320 11980 2372
rect 12032 2360 12038 2372
rect 12069 2363 12127 2369
rect 12069 2360 12081 2363
rect 12032 2332 12081 2360
rect 12032 2320 12038 2332
rect 12069 2329 12081 2332
rect 12115 2329 12127 2363
rect 12176 2360 12204 2400
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 12526 2388 12532 2440
rect 12584 2428 12590 2440
rect 13642 2431 13700 2437
rect 13642 2428 13654 2431
rect 12584 2400 13654 2428
rect 12584 2388 12590 2400
rect 13642 2397 13654 2400
rect 13688 2397 13700 2431
rect 13642 2391 13700 2397
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 14056 2400 14105 2428
rect 14056 2388 14062 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 12176 2332 12664 2360
rect 12069 2323 12127 2329
rect 3252 2264 4568 2292
rect 5905 2295 5963 2301
rect 5905 2261 5917 2295
rect 5951 2292 5963 2295
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 5951 2264 9781 2292
rect 5951 2261 5963 2264
rect 5905 2255 5963 2261
rect 9769 2261 9781 2264
rect 9815 2261 9827 2295
rect 9769 2255 9827 2261
rect 11054 2252 11060 2304
rect 11112 2292 11118 2304
rect 12529 2295 12587 2301
rect 12529 2292 12541 2295
rect 11112 2264 12541 2292
rect 11112 2252 11118 2264
rect 12529 2261 12541 2264
rect 12575 2261 12587 2295
rect 12636 2292 12664 2332
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 14369 2363 14427 2369
rect 14369 2360 14381 2363
rect 13872 2332 14381 2360
rect 13872 2320 13878 2332
rect 14369 2329 14381 2332
rect 14415 2329 14427 2363
rect 14369 2323 14427 2329
rect 14844 2292 14872 2468
rect 18598 2456 18604 2468
rect 18656 2456 18662 2508
rect 15470 2428 15476 2440
rect 15431 2400 15476 2428
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 15746 2428 15752 2440
rect 15707 2400 15752 2428
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 17126 2428 17132 2440
rect 17087 2400 17132 2428
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2397 17555 2431
rect 17862 2428 17868 2440
rect 17823 2400 17868 2428
rect 17497 2391 17555 2397
rect 14918 2320 14924 2372
rect 14976 2360 14982 2372
rect 17512 2360 17540 2391
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 18138 2388 18144 2440
rect 18196 2428 18202 2440
rect 18233 2431 18291 2437
rect 18233 2428 18245 2431
rect 18196 2400 18245 2428
rect 18196 2388 18202 2400
rect 18233 2397 18245 2400
rect 18279 2397 18291 2431
rect 18233 2391 18291 2397
rect 14976 2332 17540 2360
rect 14976 2320 14982 2332
rect 12636 2264 14872 2292
rect 16485 2295 16543 2301
rect 12529 2255 12587 2261
rect 16485 2261 16497 2295
rect 16531 2292 16543 2295
rect 17034 2292 17040 2304
rect 16531 2264 17040 2292
rect 16531 2261 16543 2264
rect 16485 2255 16543 2261
rect 17034 2252 17040 2264
rect 17092 2252 17098 2304
rect 17310 2292 17316 2304
rect 17271 2264 17316 2292
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 17678 2292 17684 2304
rect 17639 2264 17684 2292
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 18414 2292 18420 2304
rect 18375 2264 18420 2292
rect 18414 2252 18420 2264
rect 18472 2252 18478 2304
rect 1104 2202 18860 2224
rect 1104 2150 5398 2202
rect 5450 2150 5462 2202
rect 5514 2150 5526 2202
rect 5578 2150 5590 2202
rect 5642 2150 5654 2202
rect 5706 2150 9846 2202
rect 9898 2150 9910 2202
rect 9962 2150 9974 2202
rect 10026 2150 10038 2202
rect 10090 2150 10102 2202
rect 10154 2150 14294 2202
rect 14346 2150 14358 2202
rect 14410 2150 14422 2202
rect 14474 2150 14486 2202
rect 14538 2150 14550 2202
rect 14602 2150 18860 2202
rect 1104 2128 18860 2150
rect 17862 2088 17868 2100
rect 16546 2060 17868 2088
rect 4706 1980 4712 2032
rect 4764 2020 4770 2032
rect 12434 2020 12440 2032
rect 4764 1992 12440 2020
rect 4764 1980 4770 1992
rect 12434 1980 12440 1992
rect 12492 2020 12498 2032
rect 16546 2020 16574 2060
rect 17862 2048 17868 2060
rect 17920 2048 17926 2100
rect 12492 1992 16574 2020
rect 12492 1980 12498 1992
rect 16666 1980 16672 2032
rect 16724 2020 16730 2032
rect 18506 2020 18512 2032
rect 16724 1992 18512 2020
rect 16724 1980 16730 1992
rect 18506 1980 18512 1992
rect 18564 1980 18570 2032
rect 14458 1504 14464 1556
rect 14516 1544 14522 1556
rect 16022 1544 16028 1556
rect 14516 1516 16028 1544
rect 14516 1504 14522 1516
rect 16022 1504 16028 1516
rect 16080 1504 16086 1556
<< via1 >>
rect 6276 15308 6328 15360
rect 15200 15308 15252 15360
rect 3424 15240 3476 15292
rect 11244 15240 11296 15292
rect 3056 15172 3108 15224
rect 3976 15172 4028 15224
rect 7012 15172 7064 15224
rect 13544 15172 13596 15224
rect 15292 15172 15344 15224
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 3302 14662 3354 14714
rect 3366 14662 3418 14714
rect 3430 14662 3482 14714
rect 7622 14662 7674 14714
rect 7686 14662 7738 14714
rect 7750 14662 7802 14714
rect 7814 14662 7866 14714
rect 7878 14662 7930 14714
rect 12070 14662 12122 14714
rect 12134 14662 12186 14714
rect 12198 14662 12250 14714
rect 12262 14662 12314 14714
rect 12326 14662 12378 14714
rect 16518 14662 16570 14714
rect 16582 14662 16634 14714
rect 16646 14662 16698 14714
rect 16710 14662 16762 14714
rect 16774 14662 16826 14714
rect 4160 14560 4212 14612
rect 5724 14560 5776 14612
rect 9772 14492 9824 14544
rect 15292 14492 15344 14544
rect 1124 14424 1176 14476
rect 10324 14424 10376 14476
rect 14372 14424 14424 14476
rect 15108 14424 15160 14476
rect 3424 14356 3476 14408
rect 7380 14356 7432 14408
rect 10600 14356 10652 14408
rect 15200 14356 15252 14408
rect 3608 14288 3660 14340
rect 16672 14356 16724 14408
rect 4988 14263 5040 14272
rect 4988 14229 4997 14263
rect 4997 14229 5031 14263
rect 5031 14229 5040 14263
rect 4988 14220 5040 14229
rect 5540 14220 5592 14272
rect 14740 14220 14792 14272
rect 5398 14118 5450 14170
rect 5462 14118 5514 14170
rect 5526 14118 5578 14170
rect 5590 14118 5642 14170
rect 5654 14118 5706 14170
rect 9846 14118 9898 14170
rect 9910 14118 9962 14170
rect 9974 14118 10026 14170
rect 10038 14118 10090 14170
rect 10102 14118 10154 14170
rect 14294 14118 14346 14170
rect 14358 14118 14410 14170
rect 14422 14118 14474 14170
rect 14486 14118 14538 14170
rect 14550 14118 14602 14170
rect 3608 14016 3660 14068
rect 5080 14016 5132 14068
rect 3516 13948 3568 14000
rect 5908 13948 5960 14000
rect 4252 13880 4304 13932
rect 4620 13855 4672 13864
rect 4620 13821 4629 13855
rect 4629 13821 4663 13855
rect 4663 13821 4672 13855
rect 4620 13812 4672 13821
rect 4344 13744 4396 13796
rect 4988 13812 5040 13864
rect 6460 14016 6512 14068
rect 9772 14016 9824 14068
rect 10324 14059 10376 14068
rect 10324 14025 10333 14059
rect 10333 14025 10367 14059
rect 10367 14025 10376 14059
rect 10324 14016 10376 14025
rect 6092 13948 6144 14000
rect 9680 13948 9732 14000
rect 10416 13880 10468 13932
rect 11980 13948 12032 14000
rect 14280 13991 14332 14000
rect 14280 13957 14289 13991
rect 14289 13957 14323 13991
rect 14323 13957 14332 13991
rect 14280 13948 14332 13957
rect 16856 14016 16908 14068
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 15200 13948 15252 14000
rect 15292 13991 15344 14000
rect 15292 13957 15301 13991
rect 15301 13957 15335 13991
rect 15335 13957 15344 13991
rect 15292 13948 15344 13957
rect 18788 13948 18840 14000
rect 16672 13923 16724 13932
rect 16672 13889 16681 13923
rect 16681 13889 16715 13923
rect 16715 13889 16724 13923
rect 16672 13880 16724 13889
rect 10232 13812 10284 13864
rect 12440 13812 12492 13864
rect 13728 13855 13780 13864
rect 13728 13821 13737 13855
rect 13737 13821 13771 13855
rect 13771 13821 13780 13855
rect 13728 13812 13780 13821
rect 14740 13812 14792 13864
rect 5724 13744 5776 13796
rect 6828 13744 6880 13796
rect 16304 13855 16356 13864
rect 16304 13821 16313 13855
rect 16313 13821 16347 13855
rect 16347 13821 16356 13855
rect 16304 13812 16356 13821
rect 18880 13812 18932 13864
rect 2780 13676 2832 13728
rect 6000 13676 6052 13728
rect 6736 13676 6788 13728
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 3302 13574 3354 13626
rect 3366 13574 3418 13626
rect 3430 13574 3482 13626
rect 7622 13574 7674 13626
rect 7686 13574 7738 13626
rect 7750 13574 7802 13626
rect 7814 13574 7866 13626
rect 7878 13574 7930 13626
rect 12070 13574 12122 13626
rect 12134 13574 12186 13626
rect 12198 13574 12250 13626
rect 12262 13574 12314 13626
rect 12326 13574 12378 13626
rect 16518 13574 16570 13626
rect 16582 13574 16634 13626
rect 16646 13574 16698 13626
rect 16710 13574 16762 13626
rect 16774 13574 16826 13626
rect 2780 13515 2832 13524
rect 2780 13481 2789 13515
rect 2789 13481 2823 13515
rect 2823 13481 2832 13515
rect 2780 13472 2832 13481
rect 4620 13472 4672 13524
rect 5816 13472 5868 13524
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 14280 13472 14332 13524
rect 2412 13200 2464 13252
rect 5172 13379 5224 13388
rect 5172 13345 5181 13379
rect 5181 13345 5215 13379
rect 5215 13345 5224 13379
rect 5172 13336 5224 13345
rect 10968 13404 11020 13456
rect 2780 13268 2832 13320
rect 5724 13311 5776 13320
rect 4252 13200 4304 13252
rect 1308 13132 1360 13184
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 7472 13336 7524 13388
rect 4528 13175 4580 13184
rect 4528 13141 4537 13175
rect 4537 13141 4571 13175
rect 4571 13141 4580 13175
rect 4988 13175 5040 13184
rect 4528 13132 4580 13141
rect 4988 13141 4997 13175
rect 4997 13141 5031 13175
rect 5031 13141 5040 13175
rect 4988 13132 5040 13141
rect 5080 13132 5132 13184
rect 6644 13268 6696 13320
rect 6828 13268 6880 13320
rect 12440 13268 12492 13320
rect 15108 13268 15160 13320
rect 6276 13200 6328 13252
rect 13912 13200 13964 13252
rect 6644 13175 6696 13184
rect 6644 13141 6653 13175
rect 6653 13141 6687 13175
rect 6687 13141 6696 13175
rect 6644 13132 6696 13141
rect 7104 13175 7156 13184
rect 7104 13141 7113 13175
rect 7113 13141 7147 13175
rect 7147 13141 7156 13175
rect 7104 13132 7156 13141
rect 15200 13175 15252 13184
rect 15200 13141 15209 13175
rect 15209 13141 15243 13175
rect 15243 13141 15252 13175
rect 15200 13132 15252 13141
rect 5398 13030 5450 13082
rect 5462 13030 5514 13082
rect 5526 13030 5578 13082
rect 5590 13030 5642 13082
rect 5654 13030 5706 13082
rect 9846 13030 9898 13082
rect 9910 13030 9962 13082
rect 9974 13030 10026 13082
rect 10038 13030 10090 13082
rect 10102 13030 10154 13082
rect 14294 13030 14346 13082
rect 14358 13030 14410 13082
rect 14422 13030 14474 13082
rect 14486 13030 14538 13082
rect 14550 13030 14602 13082
rect 4528 12971 4580 12980
rect 4528 12937 4537 12971
rect 4537 12937 4571 12971
rect 4571 12937 4580 12971
rect 4528 12928 4580 12937
rect 5080 12928 5132 12980
rect 5816 12928 5868 12980
rect 6276 12928 6328 12980
rect 6644 12928 6696 12980
rect 7196 12928 7248 12980
rect 15016 12928 15068 12980
rect 2136 12903 2188 12912
rect 2136 12869 2145 12903
rect 2145 12869 2179 12903
rect 2179 12869 2188 12903
rect 2136 12860 2188 12869
rect 4896 12860 4948 12912
rect 6736 12860 6788 12912
rect 17868 12928 17920 12980
rect 1676 12792 1728 12844
rect 4988 12792 5040 12844
rect 4712 12767 4764 12776
rect 4712 12733 4721 12767
rect 4721 12733 4755 12767
rect 4755 12733 4764 12767
rect 4712 12724 4764 12733
rect 7012 12792 7064 12844
rect 7564 12792 7616 12844
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 13360 12835 13412 12844
rect 13360 12801 13369 12835
rect 13369 12801 13403 12835
rect 13403 12801 13412 12835
rect 13360 12792 13412 12801
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 14464 12792 14516 12844
rect 2044 12656 2096 12708
rect 7196 12724 7248 12776
rect 8208 12724 8260 12776
rect 14832 12724 14884 12776
rect 2964 12588 3016 12640
rect 3516 12588 3568 12640
rect 5908 12588 5960 12640
rect 6828 12588 6880 12640
rect 7012 12588 7064 12640
rect 7380 12588 7432 12640
rect 8116 12588 8168 12640
rect 10508 12588 10560 12640
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 3302 12486 3354 12538
rect 3366 12486 3418 12538
rect 3430 12486 3482 12538
rect 7622 12486 7674 12538
rect 7686 12486 7738 12538
rect 7750 12486 7802 12538
rect 7814 12486 7866 12538
rect 7878 12486 7930 12538
rect 12070 12486 12122 12538
rect 12134 12486 12186 12538
rect 12198 12486 12250 12538
rect 12262 12486 12314 12538
rect 12326 12486 12378 12538
rect 16518 12486 16570 12538
rect 16582 12486 16634 12538
rect 16646 12486 16698 12538
rect 16710 12486 16762 12538
rect 16774 12486 16826 12538
rect 2780 12384 2832 12436
rect 11796 12427 11848 12436
rect 11796 12393 11805 12427
rect 11805 12393 11839 12427
rect 11839 12393 11848 12427
rect 11796 12384 11848 12393
rect 6828 12316 6880 12368
rect 6920 12316 6972 12368
rect 9404 12316 9456 12368
rect 14924 12359 14976 12368
rect 2688 12248 2740 12300
rect 3332 12248 3384 12300
rect 4712 12248 4764 12300
rect 2136 12180 2188 12232
rect 3516 12180 3568 12232
rect 3700 12180 3752 12232
rect 4896 12223 4948 12232
rect 4896 12189 4905 12223
rect 4905 12189 4939 12223
rect 4939 12189 4948 12223
rect 4896 12180 4948 12189
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 2596 12112 2648 12164
rect 940 12044 992 12096
rect 2504 12044 2556 12096
rect 4528 12112 4580 12164
rect 4804 12112 4856 12164
rect 6276 12155 6328 12164
rect 6276 12121 6285 12155
rect 6285 12121 6319 12155
rect 6319 12121 6328 12155
rect 6276 12112 6328 12121
rect 7840 12291 7892 12300
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 10232 12291 10284 12300
rect 10232 12257 10241 12291
rect 10241 12257 10275 12291
rect 10275 12257 10284 12291
rect 10232 12248 10284 12257
rect 10784 12248 10836 12300
rect 12072 12248 12124 12300
rect 7104 12180 7156 12232
rect 8024 12180 8076 12232
rect 8208 12180 8260 12232
rect 11796 12180 11848 12232
rect 13084 12248 13136 12300
rect 13360 12248 13412 12300
rect 12992 12180 13044 12232
rect 14924 12325 14933 12359
rect 14933 12325 14967 12359
rect 14967 12325 14976 12359
rect 14924 12316 14976 12325
rect 15016 12316 15068 12368
rect 18144 12316 18196 12368
rect 14832 12248 14884 12300
rect 17592 12248 17644 12300
rect 17500 12180 17552 12232
rect 17868 12180 17920 12232
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 4068 12044 4120 12096
rect 4252 12087 4304 12096
rect 4252 12053 4261 12087
rect 4261 12053 4295 12087
rect 4295 12053 4304 12087
rect 4252 12044 4304 12053
rect 4436 12044 4488 12096
rect 4988 12087 5040 12096
rect 4988 12053 4997 12087
rect 4997 12053 5031 12087
rect 5031 12053 5040 12087
rect 4988 12044 5040 12053
rect 5264 12044 5316 12096
rect 5724 12044 5776 12096
rect 5816 12087 5868 12096
rect 5816 12053 5825 12087
rect 5825 12053 5859 12087
rect 5859 12053 5868 12087
rect 6460 12087 6512 12096
rect 5816 12044 5868 12053
rect 6460 12053 6469 12087
rect 6469 12053 6503 12087
rect 6503 12053 6512 12087
rect 6460 12044 6512 12053
rect 6920 12087 6972 12096
rect 6920 12053 6929 12087
rect 6929 12053 6963 12087
rect 6963 12053 6972 12087
rect 6920 12044 6972 12053
rect 7104 12044 7156 12096
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 7748 12087 7800 12096
rect 7748 12053 7757 12087
rect 7757 12053 7791 12087
rect 7791 12053 7800 12087
rect 7748 12044 7800 12053
rect 7932 12044 7984 12096
rect 8944 12087 8996 12096
rect 8944 12053 8953 12087
rect 8953 12053 8987 12087
rect 8987 12053 8996 12087
rect 8944 12044 8996 12053
rect 9312 12087 9364 12096
rect 9312 12053 9321 12087
rect 9321 12053 9355 12087
rect 9355 12053 9364 12087
rect 9312 12044 9364 12053
rect 9496 12044 9548 12096
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 10508 12044 10560 12096
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 12348 12087 12400 12096
rect 12348 12053 12357 12087
rect 12357 12053 12391 12087
rect 12391 12053 12400 12087
rect 12348 12044 12400 12053
rect 13544 12087 13596 12096
rect 13544 12053 13553 12087
rect 13553 12053 13587 12087
rect 13587 12053 13596 12087
rect 13544 12044 13596 12053
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 15016 12044 15068 12096
rect 16948 12044 17000 12096
rect 17132 12044 17184 12096
rect 17316 12044 17368 12096
rect 17684 12044 17736 12096
rect 5398 11942 5450 11994
rect 5462 11942 5514 11994
rect 5526 11942 5578 11994
rect 5590 11942 5642 11994
rect 5654 11942 5706 11994
rect 9846 11942 9898 11994
rect 9910 11942 9962 11994
rect 9974 11942 10026 11994
rect 10038 11942 10090 11994
rect 10102 11942 10154 11994
rect 14294 11942 14346 11994
rect 14358 11942 14410 11994
rect 14422 11942 14474 11994
rect 14486 11942 14538 11994
rect 14550 11942 14602 11994
rect 2504 11883 2556 11892
rect 2504 11849 2513 11883
rect 2513 11849 2547 11883
rect 2547 11849 2556 11883
rect 2504 11840 2556 11849
rect 2596 11883 2648 11892
rect 2596 11849 2605 11883
rect 2605 11849 2639 11883
rect 2639 11849 2648 11883
rect 2596 11840 2648 11849
rect 1124 11772 1176 11824
rect 2964 11840 3016 11892
rect 4068 11883 4120 11892
rect 4068 11849 4077 11883
rect 4077 11849 4111 11883
rect 4111 11849 4120 11883
rect 4068 11840 4120 11849
rect 4528 11840 4580 11892
rect 4804 11840 4856 11892
rect 4988 11883 5040 11892
rect 4988 11849 4997 11883
rect 4997 11849 5031 11883
rect 5031 11849 5040 11883
rect 4988 11840 5040 11849
rect 5264 11840 5316 11892
rect 5724 11840 5776 11892
rect 5816 11840 5868 11892
rect 6920 11883 6972 11892
rect 6920 11849 6929 11883
rect 6929 11849 6963 11883
rect 6963 11849 6972 11883
rect 6920 11840 6972 11849
rect 8208 11840 8260 11892
rect 8944 11883 8996 11892
rect 8944 11849 8953 11883
rect 8953 11849 8987 11883
rect 8987 11849 8996 11883
rect 8944 11840 8996 11849
rect 9312 11840 9364 11892
rect 9496 11840 9548 11892
rect 3332 11772 3384 11824
rect 6092 11772 6144 11824
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 2504 11704 2556 11756
rect 3516 11636 3568 11688
rect 4160 11704 4212 11756
rect 5724 11704 5776 11756
rect 6368 11772 6420 11824
rect 6644 11772 6696 11824
rect 9772 11772 9824 11824
rect 11980 11840 12032 11892
rect 12348 11840 12400 11892
rect 15108 11840 15160 11892
rect 17132 11883 17184 11892
rect 17132 11849 17141 11883
rect 17141 11849 17175 11883
rect 17175 11849 17184 11883
rect 17132 11840 17184 11849
rect 17500 11840 17552 11892
rect 17776 11840 17828 11892
rect 17960 11883 18012 11892
rect 17960 11849 17969 11883
rect 17969 11849 18003 11883
rect 18003 11849 18012 11883
rect 17960 11840 18012 11849
rect 15016 11772 15068 11824
rect 6920 11704 6972 11756
rect 7840 11704 7892 11756
rect 8944 11704 8996 11756
rect 9680 11704 9732 11756
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 11612 11704 11664 11756
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 4804 11636 4856 11688
rect 5172 11636 5224 11688
rect 6368 11636 6420 11688
rect 6736 11636 6788 11688
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 7472 11679 7524 11688
rect 7472 11645 7481 11679
rect 7481 11645 7515 11679
rect 7515 11645 7524 11679
rect 7472 11636 7524 11645
rect 8116 11636 8168 11688
rect 9128 11679 9180 11688
rect 9128 11645 9137 11679
rect 9137 11645 9171 11679
rect 9171 11645 9180 11679
rect 9128 11636 9180 11645
rect 10784 11636 10836 11688
rect 11796 11636 11848 11688
rect 12072 11679 12124 11688
rect 12072 11645 12081 11679
rect 12081 11645 12115 11679
rect 12115 11645 12124 11679
rect 12072 11636 12124 11645
rect 4344 11568 4396 11620
rect 5080 11568 5132 11620
rect 1492 11543 1544 11552
rect 1492 11509 1501 11543
rect 1501 11509 1535 11543
rect 1535 11509 1544 11543
rect 1492 11500 1544 11509
rect 3700 11500 3752 11552
rect 3884 11500 3936 11552
rect 3976 11500 4028 11552
rect 5816 11568 5868 11620
rect 7932 11568 7984 11620
rect 9680 11568 9732 11620
rect 11428 11568 11480 11620
rect 13728 11704 13780 11756
rect 14740 11704 14792 11756
rect 18236 11772 18288 11824
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 13268 11636 13320 11688
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 15108 11636 15160 11688
rect 15660 11636 15712 11688
rect 16396 11568 16448 11620
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 8300 11500 8352 11552
rect 10324 11543 10376 11552
rect 10324 11509 10333 11543
rect 10333 11509 10367 11543
rect 10367 11509 10376 11543
rect 10324 11500 10376 11509
rect 10416 11500 10468 11552
rect 11152 11500 11204 11552
rect 11336 11500 11388 11552
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 13268 11500 13320 11552
rect 13452 11500 13504 11552
rect 14740 11543 14792 11552
rect 14740 11509 14749 11543
rect 14749 11509 14783 11543
rect 14783 11509 14792 11543
rect 14740 11500 14792 11509
rect 15476 11500 15528 11552
rect 15936 11500 15988 11552
rect 17868 11500 17920 11552
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 3302 11398 3354 11450
rect 3366 11398 3418 11450
rect 3430 11398 3482 11450
rect 7622 11398 7674 11450
rect 7686 11398 7738 11450
rect 7750 11398 7802 11450
rect 7814 11398 7866 11450
rect 7878 11398 7930 11450
rect 12070 11398 12122 11450
rect 12134 11398 12186 11450
rect 12198 11398 12250 11450
rect 12262 11398 12314 11450
rect 12326 11398 12378 11450
rect 16518 11398 16570 11450
rect 16582 11398 16634 11450
rect 16646 11398 16698 11450
rect 16710 11398 16762 11450
rect 16774 11398 16826 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2780 11296 2832 11348
rect 1400 11228 1452 11280
rect 2688 11160 2740 11212
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 4252 11296 4304 11348
rect 2688 11024 2740 11076
rect 4160 11092 4212 11144
rect 6184 11296 6236 11348
rect 7196 11296 7248 11348
rect 7840 11296 7892 11348
rect 5172 11228 5224 11280
rect 4896 11203 4948 11212
rect 4896 11169 4905 11203
rect 4905 11169 4939 11203
rect 4939 11169 4948 11203
rect 4896 11160 4948 11169
rect 6552 11228 6604 11280
rect 8484 11296 8536 11348
rect 9128 11296 9180 11348
rect 6184 11203 6236 11212
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 6644 11160 6696 11212
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 7104 11160 7156 11212
rect 7748 11203 7800 11212
rect 7748 11169 7757 11203
rect 7757 11169 7791 11203
rect 7791 11169 7800 11203
rect 7748 11160 7800 11169
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 8024 11092 8076 11144
rect 4804 11024 4856 11076
rect 7288 11024 7340 11076
rect 7656 11067 7708 11076
rect 7656 11033 7665 11067
rect 7665 11033 7699 11067
rect 7699 11033 7708 11067
rect 7656 11024 7708 11033
rect 7932 11024 7984 11076
rect 1124 10956 1176 11008
rect 2596 10956 2648 11008
rect 2872 10956 2924 11008
rect 4252 10956 4304 11008
rect 4436 10956 4488 11008
rect 4988 10956 5040 11008
rect 5264 10956 5316 11008
rect 6460 10956 6512 11008
rect 7564 10999 7616 11008
rect 7564 10965 7573 10999
rect 7573 10965 7607 10999
rect 7607 10965 7616 10999
rect 8668 11024 8720 11076
rect 9404 11024 9456 11076
rect 10324 11092 10376 11144
rect 14740 11296 14792 11348
rect 14832 11296 14884 11348
rect 15016 11296 15068 11348
rect 15108 11296 15160 11348
rect 17040 11339 17092 11348
rect 10784 11203 10836 11212
rect 10784 11169 10793 11203
rect 10793 11169 10827 11203
rect 10827 11169 10836 11203
rect 10784 11160 10836 11169
rect 11428 11160 11480 11212
rect 14188 11228 14240 11280
rect 16764 11228 16816 11280
rect 17040 11305 17049 11339
rect 17049 11305 17083 11339
rect 17083 11305 17092 11339
rect 17040 11296 17092 11305
rect 18880 11296 18932 11348
rect 11336 11092 11388 11144
rect 11060 11024 11112 11076
rect 11980 11024 12032 11076
rect 7564 10956 7616 10965
rect 8300 10956 8352 11008
rect 8484 10956 8536 11008
rect 12716 11024 12768 11076
rect 13636 11160 13688 11212
rect 15568 11160 15620 11212
rect 15844 11160 15896 11212
rect 17960 11228 18012 11280
rect 18696 11228 18748 11280
rect 17592 11203 17644 11212
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 17592 11160 17644 11169
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 13176 11092 13228 11144
rect 13636 11024 13688 11076
rect 13820 11092 13872 11144
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 16120 11092 16172 11144
rect 16856 11092 16908 11144
rect 17776 11092 17828 11144
rect 18236 11135 18288 11144
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 16580 11024 16632 11076
rect 13452 10999 13504 11008
rect 13452 10965 13461 10999
rect 13461 10965 13495 10999
rect 13495 10965 13504 10999
rect 13452 10956 13504 10965
rect 13912 10956 13964 11008
rect 15108 10999 15160 11008
rect 15108 10965 15117 10999
rect 15117 10965 15151 10999
rect 15151 10965 15160 10999
rect 15108 10956 15160 10965
rect 15476 10999 15528 11008
rect 15476 10965 15485 10999
rect 15485 10965 15519 10999
rect 15519 10965 15528 10999
rect 15476 10956 15528 10965
rect 16212 10999 16264 11008
rect 16212 10965 16221 10999
rect 16221 10965 16255 10999
rect 16255 10965 16264 10999
rect 16212 10956 16264 10965
rect 16856 10956 16908 11008
rect 17132 10956 17184 11008
rect 17408 10999 17460 11008
rect 17408 10965 17417 10999
rect 17417 10965 17451 10999
rect 17451 10965 17460 10999
rect 17408 10956 17460 10965
rect 5398 10854 5450 10906
rect 5462 10854 5514 10906
rect 5526 10854 5578 10906
rect 5590 10854 5642 10906
rect 5654 10854 5706 10906
rect 9846 10854 9898 10906
rect 9910 10854 9962 10906
rect 9974 10854 10026 10906
rect 10038 10854 10090 10906
rect 10102 10854 10154 10906
rect 14294 10854 14346 10906
rect 14358 10854 14410 10906
rect 14422 10854 14474 10906
rect 14486 10854 14538 10906
rect 14550 10854 14602 10906
rect 2412 10752 2464 10804
rect 2688 10795 2740 10804
rect 2688 10761 2697 10795
rect 2697 10761 2731 10795
rect 2731 10761 2740 10795
rect 2688 10752 2740 10761
rect 3056 10752 3108 10804
rect 3424 10752 3476 10804
rect 4528 10752 4580 10804
rect 4712 10752 4764 10804
rect 4896 10752 4948 10804
rect 5080 10752 5132 10804
rect 5632 10752 5684 10804
rect 5724 10752 5776 10804
rect 7564 10752 7616 10804
rect 7656 10752 7708 10804
rect 8484 10795 8536 10804
rect 8484 10761 8493 10795
rect 8493 10761 8527 10795
rect 8527 10761 8536 10795
rect 8484 10752 8536 10761
rect 8944 10795 8996 10804
rect 8944 10761 8953 10795
rect 8953 10761 8987 10795
rect 8987 10761 8996 10795
rect 8944 10752 8996 10761
rect 9404 10795 9456 10804
rect 9404 10761 9413 10795
rect 9413 10761 9447 10795
rect 9447 10761 9456 10795
rect 9404 10752 9456 10761
rect 10600 10795 10652 10804
rect 10600 10761 10609 10795
rect 10609 10761 10643 10795
rect 10643 10761 10652 10795
rect 10600 10752 10652 10761
rect 11060 10752 11112 10804
rect 11244 10795 11296 10804
rect 11244 10761 11253 10795
rect 11253 10761 11287 10795
rect 11287 10761 11296 10795
rect 11244 10752 11296 10761
rect 2412 10616 2464 10668
rect 2688 10616 2740 10668
rect 4068 10684 4120 10736
rect 3424 10616 3476 10668
rect 4712 10659 4764 10668
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 3516 10548 3568 10600
rect 4712 10625 4721 10659
rect 4721 10625 4755 10659
rect 4755 10625 4764 10659
rect 4712 10616 4764 10625
rect 4436 10548 4488 10600
rect 6552 10684 6604 10736
rect 7288 10684 7340 10736
rect 8208 10684 8260 10736
rect 12624 10684 12676 10736
rect 12808 10752 12860 10804
rect 13452 10752 13504 10804
rect 13728 10795 13780 10804
rect 13728 10761 13737 10795
rect 13737 10761 13771 10795
rect 13771 10761 13780 10795
rect 13728 10752 13780 10761
rect 15108 10752 15160 10804
rect 16580 10752 16632 10804
rect 16764 10752 16816 10804
rect 17408 10752 17460 10804
rect 13820 10684 13872 10736
rect 6000 10659 6052 10668
rect 6000 10625 6009 10659
rect 6009 10625 6043 10659
rect 6043 10625 6052 10659
rect 6736 10659 6788 10668
rect 6000 10616 6052 10625
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 5356 10548 5408 10600
rect 7564 10616 7616 10668
rect 8300 10616 8352 10668
rect 9864 10616 9916 10668
rect 9956 10616 10008 10668
rect 14832 10616 14884 10668
rect 15016 10684 15068 10736
rect 18144 10684 18196 10736
rect 15660 10616 15712 10668
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 17868 10659 17920 10668
rect 17868 10625 17877 10659
rect 17877 10625 17911 10659
rect 17911 10625 17920 10659
rect 17868 10616 17920 10625
rect 7196 10548 7248 10600
rect 7748 10548 7800 10600
rect 8392 10548 8444 10600
rect 9496 10591 9548 10600
rect 3884 10480 3936 10532
rect 7012 10480 7064 10532
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 10324 10591 10376 10600
rect 10324 10557 10333 10591
rect 10333 10557 10367 10591
rect 10367 10557 10376 10591
rect 10324 10548 10376 10557
rect 9404 10480 9456 10532
rect 11060 10480 11112 10532
rect 12992 10548 13044 10600
rect 13728 10548 13780 10600
rect 13820 10548 13872 10600
rect 14924 10548 14976 10600
rect 16212 10591 16264 10600
rect 16212 10557 16221 10591
rect 16221 10557 16255 10591
rect 16255 10557 16264 10591
rect 16212 10548 16264 10557
rect 16304 10591 16356 10600
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 17132 10591 17184 10600
rect 16304 10548 16356 10557
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 15292 10480 15344 10532
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 6920 10412 6972 10464
rect 7564 10412 7616 10464
rect 8208 10412 8260 10464
rect 8484 10412 8536 10464
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 12624 10455 12676 10464
rect 12624 10421 12633 10455
rect 12633 10421 12667 10455
rect 12667 10421 12676 10455
rect 12624 10412 12676 10421
rect 14004 10455 14056 10464
rect 14004 10421 14013 10455
rect 14013 10421 14047 10455
rect 14047 10421 14056 10455
rect 14004 10412 14056 10421
rect 14464 10412 14516 10464
rect 15108 10412 15160 10464
rect 17592 10548 17644 10600
rect 18788 10480 18840 10532
rect 18972 10480 19024 10532
rect 19248 10480 19300 10532
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 3430 10310 3482 10362
rect 7622 10310 7674 10362
rect 7686 10310 7738 10362
rect 7750 10310 7802 10362
rect 7814 10310 7866 10362
rect 7878 10310 7930 10362
rect 12070 10310 12122 10362
rect 12134 10310 12186 10362
rect 12198 10310 12250 10362
rect 12262 10310 12314 10362
rect 12326 10310 12378 10362
rect 16518 10310 16570 10362
rect 16582 10310 16634 10362
rect 16646 10310 16698 10362
rect 16710 10310 16762 10362
rect 16774 10310 16826 10362
rect 2228 10251 2280 10260
rect 2228 10217 2237 10251
rect 2237 10217 2271 10251
rect 2271 10217 2280 10251
rect 2228 10208 2280 10217
rect 2780 10208 2832 10260
rect 4252 10208 4304 10260
rect 5816 10208 5868 10260
rect 3700 10140 3752 10192
rect 6368 10140 6420 10192
rect 7380 10208 7432 10260
rect 7748 10208 7800 10260
rect 8208 10208 8260 10260
rect 9864 10208 9916 10260
rect 10968 10208 11020 10260
rect 11060 10208 11112 10260
rect 3056 10072 3108 10124
rect 2228 10004 2280 10056
rect 4436 10072 4488 10124
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 5264 10072 5316 10081
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 6276 10115 6328 10124
rect 6276 10081 6285 10115
rect 6285 10081 6319 10115
rect 6319 10081 6328 10115
rect 6276 10072 6328 10081
rect 6460 10072 6512 10124
rect 8300 10140 8352 10192
rect 10416 10140 10468 10192
rect 4896 10004 4948 10056
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 5632 10004 5684 10056
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 7380 10072 7432 10124
rect 8116 10072 8168 10124
rect 8392 10072 8444 10124
rect 9312 10072 9364 10124
rect 9956 10115 10008 10124
rect 9956 10081 9965 10115
rect 9965 10081 9999 10115
rect 9999 10081 10008 10115
rect 9956 10072 10008 10081
rect 11796 10140 11848 10192
rect 11520 10072 11572 10124
rect 11704 10115 11756 10124
rect 11704 10081 11713 10115
rect 11713 10081 11747 10115
rect 11747 10081 11756 10115
rect 11704 10072 11756 10081
rect 12992 10072 13044 10124
rect 13912 10072 13964 10124
rect 14924 10072 14976 10124
rect 15568 10072 15620 10124
rect 16580 10115 16632 10124
rect 16580 10081 16589 10115
rect 16589 10081 16623 10115
rect 16623 10081 16632 10115
rect 16580 10072 16632 10081
rect 16764 10072 16816 10124
rect 1768 9868 1820 9920
rect 4528 9936 4580 9988
rect 5540 9936 5592 9988
rect 7196 9936 7248 9988
rect 8392 9936 8444 9988
rect 8668 10004 8720 10056
rect 9220 10004 9272 10056
rect 9680 10004 9732 10056
rect 12348 10004 12400 10056
rect 13544 10004 13596 10056
rect 14464 10047 14516 10056
rect 14464 10013 14473 10047
rect 14473 10013 14507 10047
rect 14507 10013 14516 10047
rect 14464 10004 14516 10013
rect 18972 10140 19024 10192
rect 11244 9936 11296 9988
rect 5080 9868 5132 9920
rect 5724 9868 5776 9920
rect 6460 9911 6512 9920
rect 6460 9877 6469 9911
rect 6469 9877 6503 9911
rect 6503 9877 6512 9911
rect 6460 9868 6512 9877
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 7564 9868 7616 9920
rect 7748 9868 7800 9920
rect 7840 9868 7892 9920
rect 8300 9868 8352 9920
rect 8668 9911 8720 9920
rect 8668 9877 8677 9911
rect 8677 9877 8711 9911
rect 8711 9877 8720 9911
rect 8668 9868 8720 9877
rect 8944 9911 8996 9920
rect 8944 9877 8953 9911
rect 8953 9877 8987 9911
rect 8987 9877 8996 9911
rect 8944 9868 8996 9877
rect 9220 9868 9272 9920
rect 9588 9868 9640 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 11152 9911 11204 9920
rect 11152 9877 11161 9911
rect 11161 9877 11195 9911
rect 11195 9877 11204 9911
rect 11612 9911 11664 9920
rect 11152 9868 11204 9877
rect 11612 9877 11621 9911
rect 11621 9877 11655 9911
rect 11655 9877 11664 9911
rect 11612 9868 11664 9877
rect 12624 9936 12676 9988
rect 16672 9936 16724 9988
rect 18052 10004 18104 10056
rect 18144 10004 18196 10056
rect 12532 9911 12584 9920
rect 12532 9877 12541 9911
rect 12541 9877 12575 9911
rect 12575 9877 12584 9911
rect 12900 9911 12952 9920
rect 12532 9868 12584 9877
rect 12900 9877 12909 9911
rect 12909 9877 12943 9911
rect 12943 9877 12952 9911
rect 12900 9868 12952 9877
rect 15016 9868 15068 9920
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15752 9911 15804 9920
rect 15384 9868 15436 9877
rect 15752 9877 15761 9911
rect 15761 9877 15795 9911
rect 15795 9877 15804 9911
rect 15752 9868 15804 9877
rect 17408 9868 17460 9920
rect 17960 9868 18012 9920
rect 18604 9868 18656 9920
rect 5398 9766 5450 9818
rect 5462 9766 5514 9818
rect 5526 9766 5578 9818
rect 5590 9766 5642 9818
rect 5654 9766 5706 9818
rect 9846 9766 9898 9818
rect 9910 9766 9962 9818
rect 9974 9766 10026 9818
rect 10038 9766 10090 9818
rect 10102 9766 10154 9818
rect 14294 9766 14346 9818
rect 14358 9766 14410 9818
rect 14422 9766 14474 9818
rect 14486 9766 14538 9818
rect 14550 9766 14602 9818
rect 2412 9664 2464 9716
rect 4344 9707 4396 9716
rect 4344 9673 4353 9707
rect 4353 9673 4387 9707
rect 4387 9673 4396 9707
rect 4344 9664 4396 9673
rect 5724 9664 5776 9716
rect 6000 9664 6052 9716
rect 6460 9664 6512 9716
rect 7840 9664 7892 9716
rect 3148 9596 3200 9648
rect 3608 9596 3660 9648
rect 4528 9596 4580 9648
rect 5816 9596 5868 9648
rect 5908 9596 5960 9648
rect 6920 9596 6972 9648
rect 7564 9596 7616 9648
rect 9036 9664 9088 9716
rect 9864 9707 9916 9716
rect 9864 9673 9873 9707
rect 9873 9673 9907 9707
rect 9907 9673 9916 9707
rect 9864 9664 9916 9673
rect 11612 9664 11664 9716
rect 12164 9664 12216 9716
rect 12348 9707 12400 9716
rect 12348 9673 12357 9707
rect 12357 9673 12391 9707
rect 12391 9673 12400 9707
rect 12348 9664 12400 9673
rect 12532 9664 12584 9716
rect 13544 9707 13596 9716
rect 13544 9673 13553 9707
rect 13553 9673 13587 9707
rect 13587 9673 13596 9707
rect 13544 9664 13596 9673
rect 14648 9664 14700 9716
rect 14832 9707 14884 9716
rect 14832 9673 14841 9707
rect 14841 9673 14875 9707
rect 14875 9673 14884 9707
rect 14832 9664 14884 9673
rect 15752 9664 15804 9716
rect 16672 9707 16724 9716
rect 16672 9673 16681 9707
rect 16681 9673 16715 9707
rect 16715 9673 16724 9707
rect 16672 9664 16724 9673
rect 17868 9707 17920 9716
rect 17868 9673 17877 9707
rect 17877 9673 17911 9707
rect 17911 9673 17920 9707
rect 17868 9664 17920 9673
rect 18052 9664 18104 9716
rect 2872 9528 2924 9580
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 9220 9596 9272 9648
rect 2044 9460 2096 9512
rect 4068 9460 4120 9512
rect 4344 9460 4396 9512
rect 6460 9460 6512 9512
rect 6644 9460 6696 9512
rect 2872 9392 2924 9444
rect 2228 9324 2280 9376
rect 3700 9324 3752 9376
rect 4160 9392 4212 9444
rect 4896 9392 4948 9444
rect 5448 9392 5500 9444
rect 5632 9392 5684 9444
rect 10324 9596 10376 9648
rect 9956 9571 10008 9580
rect 8668 9460 8720 9512
rect 9220 9503 9272 9512
rect 5172 9367 5224 9376
rect 5172 9333 5181 9367
rect 5181 9333 5215 9367
rect 5215 9333 5224 9367
rect 5172 9324 5224 9333
rect 6276 9324 6328 9376
rect 6552 9324 6604 9376
rect 7564 9324 7616 9376
rect 8300 9324 8352 9376
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 9956 9537 9965 9571
rect 9965 9537 9999 9571
rect 9999 9537 10008 9571
rect 9956 9528 10008 9537
rect 9772 9503 9824 9512
rect 9772 9469 9781 9503
rect 9781 9469 9815 9503
rect 9815 9469 9824 9503
rect 14372 9639 14424 9648
rect 9772 9460 9824 9469
rect 8760 9324 8812 9333
rect 9496 9324 9548 9376
rect 12716 9571 12768 9580
rect 12716 9537 12725 9571
rect 12725 9537 12759 9571
rect 12759 9537 12768 9571
rect 12716 9528 12768 9537
rect 13268 9528 13320 9580
rect 12072 9503 12124 9512
rect 12072 9469 12081 9503
rect 12081 9469 12115 9503
rect 12115 9469 12124 9503
rect 12900 9503 12952 9512
rect 12072 9460 12124 9469
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 12992 9460 13044 9512
rect 14372 9605 14381 9639
rect 14381 9605 14415 9639
rect 14415 9605 14424 9639
rect 14372 9596 14424 9605
rect 15292 9596 15344 9648
rect 15476 9596 15528 9648
rect 15936 9639 15988 9648
rect 15936 9605 15945 9639
rect 15945 9605 15979 9639
rect 15979 9605 15988 9639
rect 15936 9596 15988 9605
rect 16580 9596 16632 9648
rect 17040 9639 17092 9648
rect 17040 9605 17049 9639
rect 17049 9605 17083 9639
rect 17083 9605 17092 9639
rect 17040 9596 17092 9605
rect 17592 9596 17644 9648
rect 14096 9503 14148 9512
rect 14096 9469 14105 9503
rect 14105 9469 14139 9503
rect 14139 9469 14148 9503
rect 14096 9460 14148 9469
rect 14188 9460 14240 9512
rect 12624 9392 12676 9444
rect 17776 9528 17828 9580
rect 14832 9460 14884 9512
rect 15016 9392 15068 9444
rect 11888 9324 11940 9376
rect 12900 9324 12952 9376
rect 13636 9324 13688 9376
rect 14648 9324 14700 9376
rect 15660 9460 15712 9512
rect 16764 9460 16816 9512
rect 17040 9460 17092 9512
rect 17316 9503 17368 9512
rect 17316 9469 17325 9503
rect 17325 9469 17359 9503
rect 17359 9469 17368 9503
rect 17316 9460 17368 9469
rect 15476 9392 15528 9444
rect 16028 9392 16080 9444
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 3430 9222 3482 9274
rect 7622 9222 7674 9274
rect 7686 9222 7738 9274
rect 7750 9222 7802 9274
rect 7814 9222 7866 9274
rect 7878 9222 7930 9274
rect 12070 9222 12122 9274
rect 12134 9222 12186 9274
rect 12198 9222 12250 9274
rect 12262 9222 12314 9274
rect 12326 9222 12378 9274
rect 16518 9222 16570 9274
rect 16582 9222 16634 9274
rect 16646 9222 16698 9274
rect 16710 9222 16762 9274
rect 16774 9222 16826 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 2964 9120 3016 9172
rect 4988 9120 5040 9172
rect 8392 9120 8444 9172
rect 9680 9120 9732 9172
rect 3976 9052 4028 9104
rect 2320 8984 2372 9036
rect 2596 9027 2648 9036
rect 2596 8993 2605 9027
rect 2605 8993 2639 9027
rect 2639 8993 2648 9027
rect 2596 8984 2648 8993
rect 4712 9052 4764 9104
rect 5908 9052 5960 9104
rect 6184 9052 6236 9104
rect 8668 9052 8720 9104
rect 9956 9120 10008 9172
rect 13452 9120 13504 9172
rect 14740 9120 14792 9172
rect 14832 9120 14884 9172
rect 17040 9163 17092 9172
rect 11520 9052 11572 9104
rect 12440 9095 12492 9104
rect 12440 9061 12449 9095
rect 12449 9061 12483 9095
rect 12483 9061 12492 9095
rect 12440 9052 12492 9061
rect 13360 9052 13412 9104
rect 14372 9095 14424 9104
rect 14372 9061 14381 9095
rect 14381 9061 14415 9095
rect 14415 9061 14424 9095
rect 14372 9052 14424 9061
rect 4528 8984 4580 9036
rect 5540 9027 5592 9036
rect 5540 8993 5549 9027
rect 5549 8993 5583 9027
rect 5583 8993 5592 9027
rect 5540 8984 5592 8993
rect 3148 8916 3200 8968
rect 4620 8916 4672 8968
rect 5448 8916 5500 8968
rect 6552 8959 6604 8968
rect 1676 8823 1728 8832
rect 1676 8789 1685 8823
rect 1685 8789 1719 8823
rect 1719 8789 1728 8823
rect 1676 8780 1728 8789
rect 2964 8780 3016 8832
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 3976 8780 4028 8832
rect 5632 8848 5684 8900
rect 5816 8891 5868 8900
rect 5816 8857 5825 8891
rect 5825 8857 5859 8891
rect 5859 8857 5868 8891
rect 5816 8848 5868 8857
rect 4436 8780 4488 8832
rect 4988 8823 5040 8832
rect 4988 8789 4997 8823
rect 4997 8789 5031 8823
rect 5031 8789 5040 8823
rect 4988 8780 5040 8789
rect 5080 8823 5132 8832
rect 5080 8789 5089 8823
rect 5089 8789 5123 8823
rect 5123 8789 5132 8823
rect 5724 8823 5776 8832
rect 5080 8780 5132 8789
rect 5724 8789 5733 8823
rect 5733 8789 5767 8823
rect 5767 8789 5776 8823
rect 5724 8780 5776 8789
rect 6184 8823 6236 8832
rect 6184 8789 6193 8823
rect 6193 8789 6227 8823
rect 6227 8789 6236 8823
rect 6184 8780 6236 8789
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 6644 8916 6696 8968
rect 8760 8984 8812 9036
rect 9496 9027 9548 9036
rect 9496 8993 9505 9027
rect 9505 8993 9539 9027
rect 9539 8993 9548 9027
rect 11152 9027 11204 9036
rect 9496 8984 9548 8993
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 11428 8984 11480 9036
rect 12716 8984 12768 9036
rect 14096 8984 14148 9036
rect 17040 9129 17049 9163
rect 17049 9129 17083 9163
rect 17083 9129 17092 9163
rect 17040 9120 17092 9129
rect 17132 9120 17184 9172
rect 17500 9052 17552 9104
rect 6736 8780 6788 8832
rect 7288 8780 7340 8832
rect 8484 8916 8536 8968
rect 8944 8848 8996 8900
rect 9864 8916 9916 8968
rect 11060 8959 11112 8968
rect 8484 8780 8536 8832
rect 8760 8823 8812 8832
rect 8760 8789 8769 8823
rect 8769 8789 8803 8823
rect 8803 8789 8812 8823
rect 8760 8780 8812 8789
rect 8852 8780 8904 8832
rect 9588 8780 9640 8832
rect 9956 8780 10008 8832
rect 10416 8780 10468 8832
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 12072 8916 12124 8968
rect 12808 8916 12860 8968
rect 15568 8916 15620 8968
rect 16396 8916 16448 8968
rect 16856 8916 16908 8968
rect 16028 8848 16080 8900
rect 11980 8780 12032 8832
rect 12440 8780 12492 8832
rect 12992 8823 13044 8832
rect 12992 8789 13001 8823
rect 13001 8789 13035 8823
rect 13035 8789 13044 8823
rect 12992 8780 13044 8789
rect 13268 8823 13320 8832
rect 13268 8789 13277 8823
rect 13277 8789 13311 8823
rect 13311 8789 13320 8823
rect 13268 8780 13320 8789
rect 14188 8780 14240 8832
rect 14832 8823 14884 8832
rect 14832 8789 14841 8823
rect 14841 8789 14875 8823
rect 14875 8789 14884 8823
rect 14832 8780 14884 8789
rect 15384 8780 15436 8832
rect 15752 8823 15804 8832
rect 15752 8789 15761 8823
rect 15761 8789 15795 8823
rect 15795 8789 15804 8823
rect 15752 8780 15804 8789
rect 16212 8823 16264 8832
rect 16212 8789 16221 8823
rect 16221 8789 16255 8823
rect 16255 8789 16264 8823
rect 16212 8780 16264 8789
rect 16580 8780 16632 8832
rect 17040 8916 17092 8968
rect 17684 8916 17736 8968
rect 18236 8959 18288 8968
rect 18236 8925 18245 8959
rect 18245 8925 18279 8959
rect 18279 8925 18288 8959
rect 18236 8916 18288 8925
rect 17132 8848 17184 8900
rect 17040 8780 17092 8832
rect 17500 8780 17552 8832
rect 17684 8780 17736 8832
rect 18420 8823 18472 8832
rect 18420 8789 18429 8823
rect 18429 8789 18463 8823
rect 18463 8789 18472 8823
rect 18420 8780 18472 8789
rect 5398 8678 5450 8730
rect 5462 8678 5514 8730
rect 5526 8678 5578 8730
rect 5590 8678 5642 8730
rect 5654 8678 5706 8730
rect 9846 8678 9898 8730
rect 9910 8678 9962 8730
rect 9974 8678 10026 8730
rect 10038 8678 10090 8730
rect 10102 8678 10154 8730
rect 14294 8678 14346 8730
rect 14358 8678 14410 8730
rect 14422 8678 14474 8730
rect 14486 8678 14538 8730
rect 14550 8678 14602 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 2136 8576 2188 8628
rect 3148 8576 3200 8628
rect 3792 8576 3844 8628
rect 3884 8576 3936 8628
rect 4436 8619 4488 8628
rect 4436 8585 4445 8619
rect 4445 8585 4479 8619
rect 4479 8585 4488 8619
rect 4436 8576 4488 8585
rect 5264 8576 5316 8628
rect 6736 8576 6788 8628
rect 10508 8619 10560 8628
rect 1952 8508 2004 8560
rect 2320 8440 2372 8492
rect 4252 8508 4304 8560
rect 4620 8508 4672 8560
rect 1124 8372 1176 8424
rect 2964 8440 3016 8492
rect 5908 8508 5960 8560
rect 6552 8508 6604 8560
rect 2688 8415 2740 8424
rect 2688 8381 2697 8415
rect 2697 8381 2731 8415
rect 2731 8381 2740 8415
rect 2688 8372 2740 8381
rect 3424 8415 3476 8424
rect 3424 8381 3433 8415
rect 3433 8381 3467 8415
rect 3467 8381 3476 8415
rect 3424 8372 3476 8381
rect 4252 8372 4304 8424
rect 4896 8440 4948 8492
rect 5816 8440 5868 8492
rect 6368 8440 6420 8492
rect 7288 8508 7340 8560
rect 8392 8508 8444 8560
rect 8944 8508 8996 8560
rect 9220 8508 9272 8560
rect 6460 8372 6512 8424
rect 8208 8440 8260 8492
rect 10508 8585 10517 8619
rect 10517 8585 10551 8619
rect 10551 8585 10560 8619
rect 10508 8576 10560 8585
rect 11796 8576 11848 8628
rect 14648 8576 14700 8628
rect 16580 8576 16632 8628
rect 16948 8576 17000 8628
rect 13912 8508 13964 8560
rect 11060 8440 11112 8492
rect 11336 8440 11388 8492
rect 15568 8508 15620 8560
rect 15660 8508 15712 8560
rect 14096 8440 14148 8492
rect 16212 8440 16264 8492
rect 16764 8440 16816 8492
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 17592 8508 17644 8560
rect 17776 8508 17828 8560
rect 2228 8304 2280 8356
rect 3516 8304 3568 8356
rect 3976 8347 4028 8356
rect 3976 8313 3985 8347
rect 3985 8313 4019 8347
rect 4019 8313 4028 8347
rect 3976 8304 4028 8313
rect 4344 8304 4396 8356
rect 4436 8304 4488 8356
rect 1860 8236 1912 8288
rect 6644 8304 6696 8356
rect 6736 8304 6788 8356
rect 6552 8236 6604 8288
rect 6828 8236 6880 8288
rect 8852 8236 8904 8288
rect 13452 8415 13504 8424
rect 13452 8381 13461 8415
rect 13461 8381 13495 8415
rect 13495 8381 13504 8415
rect 13452 8372 13504 8381
rect 16396 8415 16448 8424
rect 16396 8381 16405 8415
rect 16405 8381 16439 8415
rect 16439 8381 16448 8415
rect 16396 8372 16448 8381
rect 16488 8372 16540 8424
rect 18144 8440 18196 8492
rect 14924 8347 14976 8356
rect 14924 8313 14933 8347
rect 14933 8313 14967 8347
rect 14967 8313 14976 8347
rect 14924 8304 14976 8313
rect 10968 8236 11020 8288
rect 15292 8236 15344 8288
rect 16948 8304 17000 8356
rect 17868 8304 17920 8356
rect 18052 8347 18104 8356
rect 18052 8313 18061 8347
rect 18061 8313 18095 8347
rect 18095 8313 18104 8347
rect 18052 8304 18104 8313
rect 18512 8304 18564 8356
rect 17132 8236 17184 8288
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 3430 8134 3482 8186
rect 7622 8134 7674 8186
rect 7686 8134 7738 8186
rect 7750 8134 7802 8186
rect 7814 8134 7866 8186
rect 7878 8134 7930 8186
rect 12070 8134 12122 8186
rect 12134 8134 12186 8186
rect 12198 8134 12250 8186
rect 12262 8134 12314 8186
rect 12326 8134 12378 8186
rect 16518 8134 16570 8186
rect 16582 8134 16634 8186
rect 16646 8134 16698 8186
rect 16710 8134 16762 8186
rect 16774 8134 16826 8186
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 3424 8032 3476 8084
rect 4344 8032 4396 8084
rect 5724 8032 5776 8084
rect 7288 8075 7340 8084
rect 7288 8041 7297 8075
rect 7297 8041 7331 8075
rect 7331 8041 7340 8075
rect 7288 8032 7340 8041
rect 2688 8007 2740 8016
rect 2688 7973 2697 8007
rect 2697 7973 2731 8007
rect 2731 7973 2740 8007
rect 2688 7964 2740 7973
rect 3332 7964 3384 8016
rect 3148 7896 3200 7948
rect 4160 7939 4212 7948
rect 4160 7905 4169 7939
rect 4169 7905 4203 7939
rect 4203 7905 4212 7939
rect 4160 7896 4212 7905
rect 4528 7896 4580 7948
rect 2136 7828 2188 7880
rect 2228 7828 2280 7880
rect 3332 7828 3384 7880
rect 1584 7692 1636 7744
rect 2688 7692 2740 7744
rect 3424 7760 3476 7812
rect 4252 7828 4304 7880
rect 5632 7964 5684 8016
rect 7196 7964 7248 8016
rect 14096 8032 14148 8084
rect 13912 7964 13964 8016
rect 15752 8032 15804 8084
rect 17500 8032 17552 8084
rect 18328 8032 18380 8084
rect 16948 7964 17000 8016
rect 17132 7964 17184 8016
rect 18052 8007 18104 8016
rect 18052 7973 18061 8007
rect 18061 7973 18095 8007
rect 18095 7973 18104 8007
rect 18052 7964 18104 7973
rect 5172 7896 5224 7948
rect 5080 7760 5132 7812
rect 5264 7760 5316 7812
rect 7472 7828 7524 7880
rect 9312 7896 9364 7948
rect 17316 7896 17368 7948
rect 8852 7828 8904 7880
rect 9036 7828 9088 7880
rect 9496 7828 9548 7880
rect 10232 7828 10284 7880
rect 9772 7760 9824 7812
rect 10784 7760 10836 7812
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 11428 7828 11480 7880
rect 13452 7828 13504 7880
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 16396 7828 16448 7880
rect 17224 7828 17276 7880
rect 17868 7871 17920 7880
rect 17868 7837 17877 7871
rect 17877 7837 17911 7871
rect 17911 7837 17920 7871
rect 17868 7828 17920 7837
rect 11244 7760 11296 7812
rect 3332 7735 3384 7744
rect 3332 7701 3341 7735
rect 3341 7701 3375 7735
rect 3375 7701 3384 7735
rect 3332 7692 3384 7701
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 5908 7692 5960 7744
rect 7288 7692 7340 7744
rect 9128 7692 9180 7744
rect 10508 7692 10560 7744
rect 17040 7760 17092 7812
rect 17132 7760 17184 7812
rect 17684 7760 17736 7812
rect 13544 7692 13596 7744
rect 13912 7692 13964 7744
rect 5398 7590 5450 7642
rect 5462 7590 5514 7642
rect 5526 7590 5578 7642
rect 5590 7590 5642 7642
rect 5654 7590 5706 7642
rect 9846 7590 9898 7642
rect 9910 7590 9962 7642
rect 9974 7590 10026 7642
rect 10038 7590 10090 7642
rect 10102 7590 10154 7642
rect 14294 7590 14346 7642
rect 14358 7590 14410 7642
rect 14422 7590 14474 7642
rect 14486 7590 14538 7642
rect 14550 7590 14602 7642
rect 3056 7488 3108 7540
rect 3424 7488 3476 7540
rect 3884 7531 3936 7540
rect 3884 7497 3893 7531
rect 3893 7497 3927 7531
rect 3927 7497 3936 7531
rect 3884 7488 3936 7497
rect 4804 7488 4856 7540
rect 5172 7488 5224 7540
rect 5264 7488 5316 7540
rect 3608 7420 3660 7472
rect 4528 7463 4580 7472
rect 4528 7429 4537 7463
rect 4537 7429 4571 7463
rect 4571 7429 4580 7463
rect 4528 7420 4580 7429
rect 6000 7420 6052 7472
rect 6828 7488 6880 7540
rect 7472 7488 7524 7540
rect 7656 7488 7708 7540
rect 8300 7488 8352 7540
rect 8576 7488 8628 7540
rect 12900 7531 12952 7540
rect 12900 7497 12909 7531
rect 12909 7497 12943 7531
rect 12943 7497 12952 7531
rect 12900 7488 12952 7497
rect 13360 7531 13412 7540
rect 13360 7497 13369 7531
rect 13369 7497 13403 7531
rect 13403 7497 13412 7531
rect 13360 7488 13412 7497
rect 13452 7488 13504 7540
rect 13820 7488 13872 7540
rect 14188 7488 14240 7540
rect 15292 7531 15344 7540
rect 15292 7497 15301 7531
rect 15301 7497 15335 7531
rect 15335 7497 15344 7531
rect 15292 7488 15344 7497
rect 15476 7531 15528 7540
rect 15476 7497 15485 7531
rect 15485 7497 15519 7531
rect 15519 7497 15528 7531
rect 15476 7488 15528 7497
rect 17868 7531 17920 7540
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 1492 7259 1544 7268
rect 1492 7225 1501 7259
rect 1501 7225 1535 7259
rect 1535 7225 1544 7259
rect 1492 7216 1544 7225
rect 2320 7284 2372 7336
rect 3148 7352 3200 7404
rect 2504 7191 2556 7200
rect 2504 7157 2513 7191
rect 2513 7157 2547 7191
rect 2547 7157 2556 7191
rect 2504 7148 2556 7157
rect 2964 7216 3016 7268
rect 3056 7148 3108 7200
rect 3792 7216 3844 7268
rect 4252 7352 4304 7404
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 7288 7352 7340 7404
rect 4344 7284 4396 7336
rect 4252 7216 4304 7268
rect 5908 7284 5960 7336
rect 8116 7420 8168 7472
rect 9404 7463 9456 7472
rect 8852 7352 8904 7404
rect 9404 7429 9438 7463
rect 9438 7429 9456 7463
rect 9404 7420 9456 7429
rect 11612 7420 11664 7472
rect 8944 7284 8996 7336
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 5264 7148 5316 7200
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 5908 7191 5960 7200
rect 5908 7157 5917 7191
rect 5917 7157 5951 7191
rect 5951 7157 5960 7191
rect 5908 7148 5960 7157
rect 10968 7352 11020 7404
rect 13820 7352 13872 7404
rect 11336 7327 11388 7336
rect 11336 7293 11345 7327
rect 11345 7293 11379 7327
rect 11379 7293 11388 7327
rect 11336 7284 11388 7293
rect 15752 7420 15804 7472
rect 17592 7420 17644 7472
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 16856 7352 16908 7404
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 17868 7488 17920 7497
rect 19340 7352 19392 7404
rect 15844 7284 15896 7336
rect 16212 7284 16264 7336
rect 17592 7284 17644 7336
rect 17868 7284 17920 7336
rect 18328 7327 18380 7336
rect 18328 7293 18337 7327
rect 18337 7293 18371 7327
rect 18371 7293 18380 7327
rect 18328 7284 18380 7293
rect 9496 7148 9548 7200
rect 10968 7191 11020 7200
rect 10968 7157 10977 7191
rect 10977 7157 11011 7191
rect 11011 7157 11020 7191
rect 10968 7148 11020 7157
rect 12808 7148 12860 7200
rect 15752 7191 15804 7200
rect 15752 7157 15761 7191
rect 15761 7157 15795 7191
rect 15795 7157 15804 7191
rect 15752 7148 15804 7157
rect 16304 7148 16356 7200
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 3430 7046 3482 7098
rect 7622 7046 7674 7098
rect 7686 7046 7738 7098
rect 7750 7046 7802 7098
rect 7814 7046 7866 7098
rect 7878 7046 7930 7098
rect 12070 7046 12122 7098
rect 12134 7046 12186 7098
rect 12198 7046 12250 7098
rect 12262 7046 12314 7098
rect 12326 7046 12378 7098
rect 16518 7046 16570 7098
rect 16582 7046 16634 7098
rect 16646 7046 16698 7098
rect 16710 7046 16762 7098
rect 16774 7046 16826 7098
rect 1676 6987 1728 6996
rect 1676 6953 1685 6987
rect 1685 6953 1719 6987
rect 1719 6953 1728 6987
rect 1676 6944 1728 6953
rect 2320 6944 2372 6996
rect 2596 6987 2648 6996
rect 2596 6953 2605 6987
rect 2605 6953 2639 6987
rect 2639 6953 2648 6987
rect 2596 6944 2648 6953
rect 2872 6944 2924 6996
rect 3056 6944 3108 6996
rect 3884 6987 3936 6996
rect 3884 6953 3893 6987
rect 3893 6953 3927 6987
rect 3927 6953 3936 6987
rect 3884 6944 3936 6953
rect 4068 6944 4120 6996
rect 7196 6944 7248 6996
rect 7472 6944 7524 6996
rect 9772 6944 9824 6996
rect 11428 6987 11480 6996
rect 11428 6953 11437 6987
rect 11437 6953 11471 6987
rect 11471 6953 11480 6987
rect 11428 6944 11480 6953
rect 13452 6944 13504 6996
rect 18052 6987 18104 6996
rect 2504 6876 2556 6928
rect 2136 6851 2188 6860
rect 2136 6817 2145 6851
rect 2145 6817 2179 6851
rect 2179 6817 2188 6851
rect 2136 6808 2188 6817
rect 2320 6740 2372 6792
rect 4344 6876 4396 6928
rect 5632 6876 5684 6928
rect 7380 6919 7432 6928
rect 7380 6885 7389 6919
rect 7389 6885 7423 6919
rect 7423 6885 7432 6919
rect 7380 6876 7432 6885
rect 3056 6808 3108 6860
rect 12900 6808 12952 6860
rect 13544 6876 13596 6928
rect 18052 6953 18061 6987
rect 18061 6953 18095 6987
rect 18095 6953 18104 6987
rect 18052 6944 18104 6953
rect 17040 6876 17092 6928
rect 17224 6876 17276 6928
rect 3608 6740 3660 6792
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 4344 6740 4396 6792
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 6000 6740 6052 6792
rect 7104 6740 7156 6792
rect 1492 6604 1544 6656
rect 2688 6604 2740 6656
rect 3056 6604 3108 6656
rect 3608 6647 3660 6656
rect 3608 6613 3617 6647
rect 3617 6613 3651 6647
rect 3651 6613 3660 6647
rect 3608 6604 3660 6613
rect 4804 6672 4856 6724
rect 5080 6672 5132 6724
rect 5724 6604 5776 6656
rect 7380 6672 7432 6724
rect 8668 6672 8720 6724
rect 8852 6604 8904 6656
rect 11060 6783 11112 6792
rect 11060 6749 11078 6783
rect 11078 6749 11112 6783
rect 11060 6740 11112 6749
rect 10968 6672 11020 6724
rect 12072 6740 12124 6792
rect 11704 6672 11756 6724
rect 11980 6672 12032 6724
rect 17592 6851 17644 6860
rect 17592 6817 17601 6851
rect 17601 6817 17635 6851
rect 17635 6817 17644 6851
rect 17592 6808 17644 6817
rect 18420 6808 18472 6860
rect 13636 6740 13688 6792
rect 16396 6740 16448 6792
rect 17224 6740 17276 6792
rect 16580 6672 16632 6724
rect 16856 6672 16908 6724
rect 17316 6672 17368 6724
rect 19156 6740 19208 6792
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 12992 6647 13044 6656
rect 12992 6613 13001 6647
rect 13001 6613 13035 6647
rect 13035 6613 13044 6647
rect 12992 6604 13044 6613
rect 13728 6604 13780 6656
rect 15384 6604 15436 6656
rect 15568 6647 15620 6656
rect 15568 6613 15577 6647
rect 15577 6613 15611 6647
rect 15611 6613 15620 6647
rect 15568 6604 15620 6613
rect 16120 6604 16172 6656
rect 17224 6604 17276 6656
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 5398 6502 5450 6554
rect 5462 6502 5514 6554
rect 5526 6502 5578 6554
rect 5590 6502 5642 6554
rect 5654 6502 5706 6554
rect 9846 6502 9898 6554
rect 9910 6502 9962 6554
rect 9974 6502 10026 6554
rect 10038 6502 10090 6554
rect 10102 6502 10154 6554
rect 14294 6502 14346 6554
rect 14358 6502 14410 6554
rect 14422 6502 14474 6554
rect 14486 6502 14538 6554
rect 14550 6502 14602 6554
rect 1124 6400 1176 6452
rect 3608 6400 3660 6452
rect 4620 6400 4672 6452
rect 9588 6400 9640 6452
rect 10968 6443 11020 6452
rect 1492 6264 1544 6316
rect 2412 6307 2464 6316
rect 1308 6196 1360 6248
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 3608 6307 3660 6316
rect 2136 6196 2188 6248
rect 2320 6196 2372 6248
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 5724 6332 5776 6384
rect 8392 6332 8444 6384
rect 9312 6332 9364 6384
rect 10968 6409 10977 6443
rect 10977 6409 11011 6443
rect 11011 6409 11020 6443
rect 10968 6400 11020 6409
rect 13452 6400 13504 6452
rect 10692 6332 10744 6384
rect 13544 6332 13596 6384
rect 15108 6400 15160 6452
rect 15936 6400 15988 6452
rect 17224 6443 17276 6452
rect 17224 6409 17233 6443
rect 17233 6409 17267 6443
rect 17267 6409 17276 6443
rect 17224 6400 17276 6409
rect 18328 6400 18380 6452
rect 18420 6400 18472 6452
rect 15568 6332 15620 6384
rect 3424 6239 3476 6248
rect 2964 6128 3016 6180
rect 3056 6128 3108 6180
rect 3424 6205 3433 6239
rect 3433 6205 3467 6239
rect 3467 6205 3476 6239
rect 3424 6196 3476 6205
rect 3884 6196 3936 6248
rect 4068 6196 4120 6248
rect 4436 6264 4488 6316
rect 6092 6264 6144 6316
rect 4620 6239 4672 6248
rect 4620 6205 4629 6239
rect 4629 6205 4663 6239
rect 4663 6205 4672 6239
rect 4620 6196 4672 6205
rect 4804 6239 4856 6248
rect 4804 6205 4813 6239
rect 4813 6205 4847 6239
rect 4847 6205 4856 6239
rect 4804 6196 4856 6205
rect 4528 6128 4580 6180
rect 6000 6128 6052 6180
rect 9128 6264 9180 6316
rect 1400 6060 1452 6112
rect 1676 6060 1728 6112
rect 8944 6196 8996 6248
rect 12900 6264 12952 6316
rect 12992 6264 13044 6316
rect 14096 6264 14148 6316
rect 14832 6307 14884 6316
rect 14832 6273 14841 6307
rect 14841 6273 14875 6307
rect 14875 6273 14884 6307
rect 14832 6264 14884 6273
rect 16028 6307 16080 6316
rect 18052 6332 18104 6384
rect 16028 6273 16046 6307
rect 16046 6273 16080 6307
rect 16028 6264 16080 6273
rect 16396 6264 16448 6316
rect 17500 6264 17552 6316
rect 18236 6264 18288 6316
rect 14924 6196 14976 6248
rect 16764 6239 16816 6248
rect 16764 6205 16773 6239
rect 16773 6205 16807 6239
rect 16807 6205 16816 6239
rect 17868 6239 17920 6248
rect 16764 6196 16816 6205
rect 8116 6128 8168 6180
rect 3884 6060 3936 6112
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 8300 6060 8352 6112
rect 9220 6128 9272 6180
rect 10232 6128 10284 6180
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12440 6060 12492 6069
rect 12900 6060 12952 6112
rect 13820 6128 13872 6180
rect 16580 6128 16632 6180
rect 17868 6205 17877 6239
rect 17877 6205 17911 6239
rect 17911 6205 17920 6239
rect 17868 6196 17920 6205
rect 13176 6103 13228 6112
rect 13176 6069 13185 6103
rect 13185 6069 13219 6103
rect 13219 6069 13228 6103
rect 13176 6060 13228 6069
rect 18420 6128 18472 6180
rect 17132 6060 17184 6112
rect 17316 6103 17368 6112
rect 17316 6069 17325 6103
rect 17325 6069 17359 6103
rect 17359 6069 17368 6103
rect 17316 6060 17368 6069
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 3430 5958 3482 6010
rect 7622 5958 7674 6010
rect 7686 5958 7738 6010
rect 7750 5958 7802 6010
rect 7814 5958 7866 6010
rect 7878 5958 7930 6010
rect 12070 5958 12122 6010
rect 12134 5958 12186 6010
rect 12198 5958 12250 6010
rect 12262 5958 12314 6010
rect 12326 5958 12378 6010
rect 16518 5958 16570 6010
rect 16582 5958 16634 6010
rect 16646 5958 16698 6010
rect 16710 5958 16762 6010
rect 16774 5958 16826 6010
rect 1492 5899 1544 5908
rect 1492 5865 1501 5899
rect 1501 5865 1535 5899
rect 1535 5865 1544 5899
rect 1492 5856 1544 5865
rect 2412 5856 2464 5908
rect 2872 5856 2924 5908
rect 3608 5899 3660 5908
rect 3608 5865 3617 5899
rect 3617 5865 3651 5899
rect 3651 5865 3660 5899
rect 3608 5856 3660 5865
rect 4620 5856 4672 5908
rect 1952 5720 2004 5772
rect 1860 5652 1912 5704
rect 2780 5720 2832 5772
rect 4160 5720 4212 5772
rect 3608 5652 3660 5704
rect 4436 5584 4488 5636
rect 5816 5788 5868 5840
rect 6092 5831 6144 5840
rect 6092 5797 6101 5831
rect 6101 5797 6135 5831
rect 6135 5797 6144 5831
rect 6092 5788 6144 5797
rect 4712 5652 4764 5704
rect 6368 5652 6420 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 1308 5516 1360 5568
rect 1768 5516 1820 5568
rect 4528 5559 4580 5568
rect 4528 5525 4537 5559
rect 4537 5525 4571 5559
rect 4571 5525 4580 5559
rect 4528 5516 4580 5525
rect 5908 5584 5960 5636
rect 7196 5627 7248 5636
rect 7196 5593 7214 5627
rect 7214 5593 7248 5627
rect 7196 5584 7248 5593
rect 8024 5584 8076 5636
rect 9680 5584 9732 5636
rect 10692 5652 10744 5704
rect 10968 5584 11020 5636
rect 12072 5899 12124 5908
rect 12072 5865 12081 5899
rect 12081 5865 12115 5899
rect 12115 5865 12124 5899
rect 12072 5856 12124 5865
rect 13452 5856 13504 5908
rect 15568 5899 15620 5908
rect 15568 5865 15577 5899
rect 15577 5865 15611 5899
rect 15611 5865 15620 5899
rect 15568 5856 15620 5865
rect 15660 5856 15712 5908
rect 15844 5856 15896 5908
rect 17224 5856 17276 5908
rect 16304 5720 16356 5772
rect 16856 5720 16908 5772
rect 17500 5763 17552 5772
rect 17500 5729 17509 5763
rect 17509 5729 17543 5763
rect 17543 5729 17552 5763
rect 17500 5720 17552 5729
rect 12072 5652 12124 5704
rect 13452 5695 13504 5704
rect 13452 5661 13461 5695
rect 13461 5661 13495 5695
rect 13495 5661 13504 5695
rect 13452 5652 13504 5661
rect 14832 5652 14884 5704
rect 17316 5652 17368 5704
rect 13820 5584 13872 5636
rect 15108 5584 15160 5636
rect 16764 5584 16816 5636
rect 17592 5584 17644 5636
rect 6000 5516 6052 5568
rect 6092 5516 6144 5568
rect 10232 5516 10284 5568
rect 11888 5516 11940 5568
rect 12072 5516 12124 5568
rect 15660 5516 15712 5568
rect 16120 5559 16172 5568
rect 16120 5525 16129 5559
rect 16129 5525 16163 5559
rect 16163 5525 16172 5559
rect 16120 5516 16172 5525
rect 16212 5516 16264 5568
rect 17316 5559 17368 5568
rect 17316 5525 17325 5559
rect 17325 5525 17359 5559
rect 17359 5525 17368 5559
rect 17316 5516 17368 5525
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18144 5516 18196 5525
rect 18236 5559 18288 5568
rect 18236 5525 18245 5559
rect 18245 5525 18279 5559
rect 18279 5525 18288 5559
rect 18236 5516 18288 5525
rect 5398 5414 5450 5466
rect 5462 5414 5514 5466
rect 5526 5414 5578 5466
rect 5590 5414 5642 5466
rect 5654 5414 5706 5466
rect 9846 5414 9898 5466
rect 9910 5414 9962 5466
rect 9974 5414 10026 5466
rect 10038 5414 10090 5466
rect 10102 5414 10154 5466
rect 14294 5414 14346 5466
rect 14358 5414 14410 5466
rect 14422 5414 14474 5466
rect 14486 5414 14538 5466
rect 14550 5414 14602 5466
rect 2780 5312 2832 5364
rect 3976 5355 4028 5364
rect 3976 5321 3985 5355
rect 3985 5321 4019 5355
rect 4019 5321 4028 5355
rect 3976 5312 4028 5321
rect 4804 5312 4856 5364
rect 6368 5355 6420 5364
rect 6368 5321 6377 5355
rect 6377 5321 6411 5355
rect 6411 5321 6420 5355
rect 6368 5312 6420 5321
rect 6460 5312 6512 5364
rect 13912 5312 13964 5364
rect 4160 5244 4212 5296
rect 4712 5244 4764 5296
rect 2228 5176 2280 5228
rect 2504 5176 2556 5228
rect 3056 5176 3108 5228
rect 4344 5176 4396 5228
rect 4528 5176 4580 5228
rect 5632 5219 5684 5228
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5176 5684 5185
rect 6644 5219 6696 5228
rect 2688 5108 2740 5160
rect 2872 5108 2924 5160
rect 4436 5108 4488 5160
rect 4528 5040 4580 5092
rect 4988 5151 5040 5160
rect 4988 5117 4997 5151
rect 4997 5117 5031 5151
rect 5031 5117 5040 5151
rect 5724 5151 5776 5160
rect 4988 5108 5040 5117
rect 5724 5117 5733 5151
rect 5733 5117 5767 5151
rect 5767 5117 5776 5151
rect 5724 5108 5776 5117
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 6920 5219 6972 5228
rect 6920 5185 6954 5219
rect 6954 5185 6972 5219
rect 6920 5176 6972 5185
rect 9680 5244 9732 5296
rect 8668 5176 8720 5228
rect 10968 5244 11020 5296
rect 11796 5287 11848 5296
rect 11796 5253 11830 5287
rect 11830 5253 11848 5287
rect 11796 5244 11848 5253
rect 13820 5244 13872 5296
rect 9956 5219 10008 5228
rect 9956 5185 9965 5219
rect 9965 5185 9999 5219
rect 9999 5185 10008 5219
rect 9956 5176 10008 5185
rect 11612 5176 11664 5228
rect 13176 5176 13228 5228
rect 14832 5244 14884 5296
rect 15568 5312 15620 5364
rect 16396 5355 16448 5364
rect 16396 5321 16405 5355
rect 16405 5321 16439 5355
rect 16439 5321 16448 5355
rect 16396 5312 16448 5321
rect 17316 5312 17368 5364
rect 18236 5355 18288 5364
rect 18236 5321 18245 5355
rect 18245 5321 18279 5355
rect 18279 5321 18288 5355
rect 18236 5312 18288 5321
rect 18328 5355 18380 5364
rect 18328 5321 18337 5355
rect 18337 5321 18371 5355
rect 18371 5321 18380 5355
rect 18328 5312 18380 5321
rect 15476 5176 15528 5228
rect 16948 5244 17000 5296
rect 17500 5244 17552 5296
rect 16304 5176 16356 5228
rect 17408 5176 17460 5228
rect 16764 5151 16816 5160
rect 8024 5083 8076 5092
rect 8024 5049 8033 5083
rect 8033 5049 8067 5083
rect 8067 5049 8076 5083
rect 8024 5040 8076 5049
rect 9404 5040 9456 5092
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 2780 5015 2832 5024
rect 2780 4981 2789 5015
rect 2789 4981 2823 5015
rect 2823 4981 2832 5015
rect 2780 4972 2832 4981
rect 3792 4972 3844 5024
rect 4344 4972 4396 5024
rect 5632 4972 5684 5024
rect 13084 5040 13136 5092
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 16764 5117 16773 5151
rect 16773 5117 16807 5151
rect 16807 5117 16816 5151
rect 16764 5108 16816 5117
rect 16948 5151 17000 5160
rect 16948 5117 16957 5151
rect 16957 5117 16991 5151
rect 16991 5117 17000 5151
rect 16948 5108 17000 5117
rect 17316 5108 17368 5160
rect 16028 5040 16080 5092
rect 16672 5040 16724 5092
rect 17224 5040 17276 5092
rect 18328 5176 18380 5228
rect 12992 4972 13044 4981
rect 19156 4972 19208 5024
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 3430 4870 3482 4922
rect 7622 4870 7674 4922
rect 7686 4870 7738 4922
rect 7750 4870 7802 4922
rect 7814 4870 7866 4922
rect 7878 4870 7930 4922
rect 12070 4870 12122 4922
rect 12134 4870 12186 4922
rect 12198 4870 12250 4922
rect 12262 4870 12314 4922
rect 12326 4870 12378 4922
rect 16518 4870 16570 4922
rect 16582 4870 16634 4922
rect 16646 4870 16698 4922
rect 16710 4870 16762 4922
rect 16774 4870 16826 4922
rect 1952 4768 2004 4820
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 5080 4768 5132 4820
rect 8024 4768 8076 4820
rect 8852 4768 8904 4820
rect 9956 4811 10008 4820
rect 9956 4777 9965 4811
rect 9965 4777 9999 4811
rect 9999 4777 10008 4811
rect 9956 4768 10008 4777
rect 10232 4768 10284 4820
rect 10416 4768 10468 4820
rect 12992 4768 13044 4820
rect 13452 4811 13504 4820
rect 13452 4777 13461 4811
rect 13461 4777 13495 4811
rect 13495 4777 13504 4811
rect 13452 4768 13504 4777
rect 3056 4700 3108 4752
rect 2136 4675 2188 4684
rect 2136 4641 2145 4675
rect 2145 4641 2179 4675
rect 2179 4641 2188 4675
rect 2136 4632 2188 4641
rect 2780 4632 2832 4684
rect 3424 4700 3476 4752
rect 4068 4700 4120 4752
rect 5908 4743 5960 4752
rect 5908 4709 5917 4743
rect 5917 4709 5951 4743
rect 5951 4709 5960 4743
rect 5908 4700 5960 4709
rect 9680 4700 9732 4752
rect 4252 4564 4304 4616
rect 2964 4496 3016 4548
rect 3240 4539 3292 4548
rect 3240 4505 3249 4539
rect 3249 4505 3283 4539
rect 3283 4505 3292 4539
rect 3240 4496 3292 4505
rect 3056 4428 3108 4480
rect 4068 4428 4120 4480
rect 9312 4632 9364 4684
rect 13544 4700 13596 4752
rect 15568 4632 15620 4684
rect 17040 4768 17092 4820
rect 17592 4768 17644 4820
rect 18144 4768 18196 4820
rect 18420 4811 18472 4820
rect 18420 4777 18429 4811
rect 18429 4777 18463 4811
rect 18463 4777 18472 4811
rect 18420 4768 18472 4777
rect 6644 4564 6696 4616
rect 7472 4564 7524 4616
rect 8484 4564 8536 4616
rect 9404 4607 9456 4616
rect 9404 4573 9413 4607
rect 9413 4573 9447 4607
rect 9447 4573 9456 4607
rect 9404 4564 9456 4573
rect 9772 4564 9824 4616
rect 4712 4539 4764 4548
rect 4712 4505 4746 4539
rect 4746 4505 4764 4539
rect 4712 4496 4764 4505
rect 4804 4496 4856 4548
rect 6920 4496 6972 4548
rect 7012 4539 7064 4548
rect 7012 4505 7030 4539
rect 7030 4505 7064 4539
rect 7012 4496 7064 4505
rect 9496 4496 9548 4548
rect 6000 4428 6052 4480
rect 10416 4496 10468 4548
rect 12900 4564 12952 4616
rect 15752 4564 15804 4616
rect 16672 4632 16724 4684
rect 16856 4632 16908 4684
rect 17040 4632 17092 4684
rect 17316 4675 17368 4684
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 17592 4607 17644 4616
rect 14096 4496 14148 4548
rect 15200 4539 15252 4548
rect 15200 4505 15218 4539
rect 15218 4505 15252 4539
rect 15200 4496 15252 4505
rect 11612 4471 11664 4480
rect 11612 4437 11621 4471
rect 11621 4437 11655 4471
rect 11655 4437 11664 4471
rect 11612 4428 11664 4437
rect 16672 4496 16724 4548
rect 17224 4496 17276 4548
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 18512 4564 18564 4616
rect 19248 4564 19300 4616
rect 17776 4496 17828 4548
rect 15936 4428 15988 4480
rect 16212 4428 16264 4480
rect 16396 4471 16448 4480
rect 16396 4437 16405 4471
rect 16405 4437 16439 4471
rect 16439 4437 16448 4471
rect 16396 4428 16448 4437
rect 16856 4471 16908 4480
rect 16856 4437 16865 4471
rect 16865 4437 16899 4471
rect 16899 4437 16908 4471
rect 16856 4428 16908 4437
rect 17132 4428 17184 4480
rect 18236 4471 18288 4480
rect 18236 4437 18245 4471
rect 18245 4437 18279 4471
rect 18279 4437 18288 4471
rect 18236 4428 18288 4437
rect 5398 4326 5450 4378
rect 5462 4326 5514 4378
rect 5526 4326 5578 4378
rect 5590 4326 5642 4378
rect 5654 4326 5706 4378
rect 9846 4326 9898 4378
rect 9910 4326 9962 4378
rect 9974 4326 10026 4378
rect 10038 4326 10090 4378
rect 10102 4326 10154 4378
rect 14294 4326 14346 4378
rect 14358 4326 14410 4378
rect 14422 4326 14474 4378
rect 14486 4326 14538 4378
rect 14550 4326 14602 4378
rect 3240 4224 3292 4276
rect 1584 4156 1636 4208
rect 3424 4199 3476 4208
rect 3424 4165 3433 4199
rect 3433 4165 3467 4199
rect 3467 4165 3476 4199
rect 3424 4156 3476 4165
rect 4252 4224 4304 4276
rect 6736 4224 6788 4276
rect 9312 4224 9364 4276
rect 11612 4267 11664 4276
rect 11612 4233 11621 4267
rect 11621 4233 11655 4267
rect 11655 4233 11664 4267
rect 11612 4224 11664 4233
rect 13452 4224 13504 4276
rect 4160 4156 4212 4208
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 2596 4088 2648 4140
rect 9588 4156 9640 4208
rect 4436 4088 4488 4140
rect 4160 4063 4212 4072
rect 4160 4029 4169 4063
rect 4169 4029 4203 4063
rect 4203 4029 4212 4063
rect 4160 4020 4212 4029
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 4620 3952 4672 4004
rect 6184 4088 6236 4140
rect 8024 4131 8076 4140
rect 8024 4097 8042 4131
rect 8042 4097 8076 4131
rect 9772 4131 9824 4140
rect 8024 4088 8076 4097
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 9956 4088 10008 4140
rect 12808 4088 12860 4140
rect 16396 4224 16448 4276
rect 16948 4224 17000 4276
rect 17776 4224 17828 4276
rect 18144 4267 18196 4276
rect 18144 4233 18153 4267
rect 18153 4233 18187 4267
rect 18187 4233 18196 4267
rect 18144 4224 18196 4233
rect 16120 4156 16172 4208
rect 1676 3884 1728 3936
rect 1952 3884 2004 3936
rect 4252 3884 4304 3936
rect 5724 3884 5776 3936
rect 7012 3884 7064 3936
rect 8392 4020 8444 4072
rect 14188 4088 14240 4140
rect 16304 4088 16356 4140
rect 17500 4088 17552 4140
rect 17960 4131 18012 4140
rect 17960 4097 17969 4131
rect 17969 4097 18003 4131
rect 18003 4097 18012 4131
rect 17960 4088 18012 4097
rect 19340 4088 19392 4140
rect 15476 4020 15528 4072
rect 11244 3995 11296 4004
rect 11244 3961 11253 3995
rect 11253 3961 11287 3995
rect 11287 3961 11296 3995
rect 11244 3952 11296 3961
rect 12532 3952 12584 4004
rect 17316 4020 17368 4072
rect 17408 4020 17460 4072
rect 10232 3884 10284 3936
rect 10784 3884 10836 3936
rect 15108 3884 15160 3936
rect 16304 3952 16356 4004
rect 17776 4020 17828 4072
rect 19064 4020 19116 4072
rect 15752 3884 15804 3936
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 3430 3782 3482 3834
rect 7622 3782 7674 3834
rect 7686 3782 7738 3834
rect 7750 3782 7802 3834
rect 7814 3782 7866 3834
rect 7878 3782 7930 3834
rect 12070 3782 12122 3834
rect 12134 3782 12186 3834
rect 12198 3782 12250 3834
rect 12262 3782 12314 3834
rect 12326 3782 12378 3834
rect 16518 3782 16570 3834
rect 16582 3782 16634 3834
rect 16646 3782 16698 3834
rect 16710 3782 16762 3834
rect 16774 3782 16826 3834
rect 1584 3680 1636 3732
rect 2320 3680 2372 3732
rect 4804 3723 4856 3732
rect 4804 3689 4813 3723
rect 4813 3689 4847 3723
rect 4847 3689 4856 3723
rect 4804 3680 4856 3689
rect 1216 3612 1268 3664
rect 2504 3612 2556 3664
rect 2596 3612 2648 3664
rect 2964 3612 3016 3664
rect 4712 3612 4764 3664
rect 2412 3544 2464 3596
rect 2044 3408 2096 3460
rect 2780 3519 2832 3528
rect 2780 3485 2789 3519
rect 2789 3485 2823 3519
rect 2823 3485 2832 3519
rect 2780 3476 2832 3485
rect 3056 3544 3108 3596
rect 3516 3476 3568 3528
rect 4528 3544 4580 3596
rect 6368 3680 6420 3732
rect 11152 3680 11204 3732
rect 11428 3680 11480 3732
rect 13452 3723 13504 3732
rect 13452 3689 13461 3723
rect 13461 3689 13495 3723
rect 13495 3689 13504 3723
rect 13452 3680 13504 3689
rect 15200 3680 15252 3732
rect 15476 3680 15528 3732
rect 17224 3680 17276 3732
rect 18052 3680 18104 3732
rect 8024 3612 8076 3664
rect 6644 3476 6696 3528
rect 8392 3544 8444 3596
rect 8484 3476 8536 3528
rect 3056 3408 3108 3460
rect 4436 3451 4488 3460
rect 4436 3417 4445 3451
rect 4445 3417 4479 3451
rect 4479 3417 4488 3451
rect 4436 3408 4488 3417
rect 4620 3408 4672 3460
rect 4712 3340 4764 3392
rect 6460 3408 6512 3460
rect 8208 3408 8260 3460
rect 8668 3408 8720 3460
rect 8852 3612 8904 3664
rect 15568 3544 15620 3596
rect 17868 3544 17920 3596
rect 9956 3408 10008 3460
rect 10140 3451 10192 3460
rect 10140 3417 10158 3451
rect 10158 3417 10192 3451
rect 10140 3408 10192 3417
rect 11612 3476 11664 3528
rect 11704 3476 11756 3528
rect 10876 3408 10928 3460
rect 8760 3340 8812 3392
rect 9680 3340 9732 3392
rect 10508 3340 10560 3392
rect 13544 3476 13596 3528
rect 15844 3476 15896 3528
rect 17224 3476 17276 3528
rect 17684 3476 17736 3528
rect 15660 3408 15712 3460
rect 17040 3408 17092 3460
rect 17960 3476 18012 3528
rect 16580 3340 16632 3392
rect 17408 3340 17460 3392
rect 17592 3340 17644 3392
rect 5398 3238 5450 3290
rect 5462 3238 5514 3290
rect 5526 3238 5578 3290
rect 5590 3238 5642 3290
rect 5654 3238 5706 3290
rect 9846 3238 9898 3290
rect 9910 3238 9962 3290
rect 9974 3238 10026 3290
rect 10038 3238 10090 3290
rect 10102 3238 10154 3290
rect 14294 3238 14346 3290
rect 14358 3238 14410 3290
rect 14422 3238 14474 3290
rect 14486 3238 14538 3290
rect 14550 3238 14602 3290
rect 2412 3068 2464 3120
rect 2596 3068 2648 3120
rect 3700 3136 3752 3188
rect 4252 3179 4304 3188
rect 4252 3145 4261 3179
rect 4261 3145 4295 3179
rect 4295 3145 4304 3179
rect 4252 3136 4304 3145
rect 4344 3179 4396 3188
rect 4344 3145 4353 3179
rect 4353 3145 4387 3179
rect 4387 3145 4396 3179
rect 4344 3136 4396 3145
rect 5632 3136 5684 3188
rect 5264 3068 5316 3120
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 3608 3000 3660 3052
rect 6644 3068 6696 3120
rect 8116 3136 8168 3188
rect 2872 2864 2924 2916
rect 4160 2975 4212 2984
rect 4160 2941 4169 2975
rect 4169 2941 4203 2975
rect 4203 2941 4212 2975
rect 4160 2932 4212 2941
rect 4528 2864 4580 2916
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 4896 2864 4948 2916
rect 6092 3000 6144 3052
rect 6920 3000 6972 3052
rect 8576 3068 8628 3120
rect 8760 3111 8812 3120
rect 8760 3077 8794 3111
rect 8794 3077 8812 3111
rect 8760 3068 8812 3077
rect 9220 3136 9272 3188
rect 10324 3136 10376 3188
rect 6184 2975 6236 2984
rect 6184 2941 6193 2975
rect 6193 2941 6227 2975
rect 6227 2941 6236 2975
rect 6184 2932 6236 2941
rect 6644 2932 6696 2984
rect 9036 3000 9088 3052
rect 9588 3068 9640 3120
rect 14464 3179 14516 3188
rect 10508 3068 10560 3120
rect 10784 3000 10836 3052
rect 11060 3043 11112 3052
rect 11060 3009 11078 3043
rect 11078 3009 11112 3043
rect 11060 3000 11112 3009
rect 8116 2932 8168 2984
rect 8484 2975 8536 2984
rect 6736 2864 6788 2916
rect 6368 2839 6420 2848
rect 6368 2805 6377 2839
rect 6377 2805 6411 2839
rect 6411 2805 6420 2839
rect 6368 2796 6420 2805
rect 8024 2796 8076 2848
rect 8484 2941 8493 2975
rect 8493 2941 8527 2975
rect 8527 2941 8536 2975
rect 8484 2932 8536 2941
rect 11612 3068 11664 3120
rect 13452 3068 13504 3120
rect 13084 3000 13136 3052
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 15568 3111 15620 3120
rect 15568 3077 15586 3111
rect 15586 3077 15620 3111
rect 16856 3136 16908 3188
rect 18328 3136 18380 3188
rect 15568 3068 15620 3077
rect 15844 3043 15896 3052
rect 15844 3009 15853 3043
rect 15853 3009 15887 3043
rect 15887 3009 15896 3043
rect 15844 3000 15896 3009
rect 15936 3043 15988 3052
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 16580 3000 16632 3052
rect 17040 3000 17092 3052
rect 17132 3000 17184 3052
rect 16028 2932 16080 2984
rect 17868 2932 17920 2984
rect 10324 2796 10376 2848
rect 14096 2864 14148 2916
rect 14372 2907 14424 2916
rect 14372 2873 14381 2907
rect 14381 2873 14415 2907
rect 14415 2873 14424 2907
rect 14372 2864 14424 2873
rect 16856 2907 16908 2916
rect 16856 2873 16865 2907
rect 16865 2873 16899 2907
rect 16899 2873 16908 2907
rect 16856 2864 16908 2873
rect 17500 2864 17552 2916
rect 11152 2796 11204 2848
rect 12900 2796 12952 2848
rect 15476 2796 15528 2848
rect 17040 2796 17092 2848
rect 17316 2796 17368 2848
rect 18144 2796 18196 2848
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 3430 2694 3482 2746
rect 7622 2694 7674 2746
rect 7686 2694 7738 2746
rect 7750 2694 7802 2746
rect 7814 2694 7866 2746
rect 7878 2694 7930 2746
rect 12070 2694 12122 2746
rect 12134 2694 12186 2746
rect 12198 2694 12250 2746
rect 12262 2694 12314 2746
rect 12326 2694 12378 2746
rect 16518 2694 16570 2746
rect 16582 2694 16634 2746
rect 16646 2694 16698 2746
rect 16710 2694 16762 2746
rect 16774 2694 16826 2746
rect 1308 2592 1360 2644
rect 2688 2635 2740 2644
rect 2688 2601 2697 2635
rect 2697 2601 2731 2635
rect 2731 2601 2740 2635
rect 2688 2592 2740 2601
rect 3056 2635 3108 2644
rect 3056 2601 3065 2635
rect 3065 2601 3099 2635
rect 3099 2601 3108 2635
rect 3056 2592 3108 2601
rect 1216 2524 1268 2576
rect 2780 2456 2832 2508
rect 2504 2431 2556 2440
rect 2504 2397 2513 2431
rect 2513 2397 2547 2431
rect 2547 2397 2556 2431
rect 2504 2388 2556 2397
rect 3884 2456 3936 2508
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 6000 2592 6052 2644
rect 6184 2635 6236 2644
rect 6184 2601 6193 2635
rect 6193 2601 6227 2635
rect 6227 2601 6236 2635
rect 6184 2592 6236 2601
rect 7472 2592 7524 2644
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 9404 2592 9456 2644
rect 11612 2635 11664 2644
rect 11612 2601 11621 2635
rect 11621 2601 11655 2635
rect 11655 2601 11664 2635
rect 11612 2592 11664 2601
rect 15844 2635 15896 2644
rect 4160 2456 4212 2508
rect 4804 2456 4856 2508
rect 4344 2388 4396 2440
rect 4436 2388 4488 2440
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 5632 2456 5684 2508
rect 9680 2456 9732 2508
rect 15844 2601 15853 2635
rect 15853 2601 15887 2635
rect 15887 2601 15896 2635
rect 15844 2592 15896 2601
rect 16672 2524 16724 2576
rect 16856 2524 16908 2576
rect 17132 2592 17184 2644
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 17224 2524 17276 2576
rect 4712 2388 4764 2397
rect 6460 2431 6512 2440
rect 6460 2397 6469 2431
rect 6469 2397 6503 2431
rect 6503 2397 6512 2431
rect 6460 2388 6512 2397
rect 3700 2320 3752 2372
rect 8300 2388 8352 2440
rect 12348 2431 12400 2440
rect 7840 2320 7892 2372
rect 7932 2320 7984 2372
rect 9220 2320 9272 2372
rect 9680 2363 9732 2372
rect 9680 2329 9689 2363
rect 9689 2329 9723 2363
rect 9723 2329 9732 2363
rect 9680 2320 9732 2329
rect 11980 2320 12032 2372
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 12532 2388 12584 2440
rect 14004 2388 14056 2440
rect 11060 2252 11112 2304
rect 13820 2320 13872 2372
rect 18604 2456 18656 2508
rect 15476 2431 15528 2440
rect 15476 2397 15485 2431
rect 15485 2397 15519 2431
rect 15519 2397 15528 2431
rect 15476 2388 15528 2397
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 17868 2431 17920 2440
rect 14924 2320 14976 2372
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 18144 2388 18196 2440
rect 17040 2252 17092 2304
rect 17316 2295 17368 2304
rect 17316 2261 17325 2295
rect 17325 2261 17359 2295
rect 17359 2261 17368 2295
rect 17316 2252 17368 2261
rect 17684 2295 17736 2304
rect 17684 2261 17693 2295
rect 17693 2261 17727 2295
rect 17727 2261 17736 2295
rect 17684 2252 17736 2261
rect 18420 2295 18472 2304
rect 18420 2261 18429 2295
rect 18429 2261 18463 2295
rect 18463 2261 18472 2295
rect 18420 2252 18472 2261
rect 5398 2150 5450 2202
rect 5462 2150 5514 2202
rect 5526 2150 5578 2202
rect 5590 2150 5642 2202
rect 5654 2150 5706 2202
rect 9846 2150 9898 2202
rect 9910 2150 9962 2202
rect 9974 2150 10026 2202
rect 10038 2150 10090 2202
rect 10102 2150 10154 2202
rect 14294 2150 14346 2202
rect 14358 2150 14410 2202
rect 14422 2150 14474 2202
rect 14486 2150 14538 2202
rect 14550 2150 14602 2202
rect 4712 1980 4764 2032
rect 12440 1980 12492 2032
rect 17868 2048 17920 2100
rect 16672 1980 16724 2032
rect 18512 1980 18564 2032
rect 14464 1504 14516 1556
rect 16028 1504 16080 1556
<< metal2 >>
rect 1122 16400 1178 17200
rect 3330 16538 3386 17200
rect 4434 16688 4490 16697
rect 4434 16623 4490 16632
rect 3330 16510 3648 16538
rect 3330 16400 3386 16510
rect 1136 14482 1164 16400
rect 3422 15464 3478 15473
rect 3422 15399 3478 15408
rect 3436 15298 3464 15399
rect 3424 15292 3476 15298
rect 3424 15234 3476 15240
rect 3056 15224 3108 15230
rect 3056 15166 3108 15172
rect 2778 14648 2834 14657
rect 2778 14583 2834 14592
rect 1124 14476 1176 14482
rect 1124 14418 1176 14424
rect 2792 13734 2820 14583
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2792 13530 2820 13670
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2792 13326 2820 13466
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2412 13252 2464 13258
rect 2412 13194 2464 13200
rect 1308 13184 1360 13190
rect 1308 13126 1360 13132
rect 940 12096 992 12102
rect 940 12038 992 12044
rect 952 5273 980 12038
rect 1124 11824 1176 11830
rect 1124 11766 1176 11772
rect 1136 11014 1164 11766
rect 1214 11384 1270 11393
rect 1214 11319 1270 11328
rect 1124 11008 1176 11014
rect 1124 10950 1176 10956
rect 1136 10169 1164 10950
rect 1122 10160 1178 10169
rect 1122 10095 1178 10104
rect 1124 8424 1176 8430
rect 1124 8366 1176 8372
rect 1136 6458 1164 8366
rect 1124 6452 1176 6458
rect 1124 6394 1176 6400
rect 938 5264 994 5273
rect 938 5199 994 5208
rect 1228 3670 1256 11319
rect 1320 6254 1348 13126
rect 1858 13016 1914 13025
rect 1858 12951 1914 12960
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1688 11762 1716 12786
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1400 11280 1452 11286
rect 1400 11222 1452 11228
rect 1308 6248 1360 6254
rect 1412 6225 1440 11222
rect 1504 7721 1532 11494
rect 1688 11354 1716 11698
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1766 10568 1822 10577
rect 1766 10503 1822 10512
rect 1780 10033 1808 10503
rect 1766 10024 1822 10033
rect 1766 9959 1822 9968
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 8537 1716 8774
rect 1674 8528 1730 8537
rect 1674 8463 1730 8472
rect 1674 7848 1730 7857
rect 1674 7783 1730 7792
rect 1584 7744 1636 7750
rect 1490 7712 1546 7721
rect 1584 7686 1636 7692
rect 1490 7647 1546 7656
rect 1490 7304 1546 7313
rect 1490 7239 1492 7248
rect 1544 7239 1546 7248
rect 1492 7210 1544 7216
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 1504 6662 1532 6831
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1596 6497 1624 7686
rect 1688 7410 1716 7783
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1688 7002 1716 7346
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1582 6488 1638 6497
rect 1582 6423 1638 6432
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1308 6190 1360 6196
rect 1398 6216 1454 6225
rect 1320 5574 1348 6190
rect 1398 6151 1454 6160
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1308 5568 1360 5574
rect 1308 5510 1360 5516
rect 1216 3664 1268 3670
rect 1268 3624 1348 3652
rect 1216 3606 1268 3612
rect 1320 2650 1348 3624
rect 1308 2644 1360 2650
rect 1308 2586 1360 2592
rect 1216 2576 1268 2582
rect 1216 2518 1268 2524
rect 1228 800 1256 2518
rect 1412 1193 1440 6054
rect 1504 5914 1532 6258
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1504 3233 1532 4966
rect 1584 4208 1636 4214
rect 1584 4150 1636 4156
rect 1596 3738 1624 4150
rect 1688 4049 1716 6054
rect 1780 5681 1808 9862
rect 1872 8378 1900 12951
rect 2136 12912 2188 12918
rect 2136 12854 2188 12860
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 2056 11744 2084 12650
rect 2148 12238 2176 12854
rect 2226 12744 2282 12753
rect 2226 12679 2282 12688
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2136 11756 2188 11762
rect 2056 11716 2136 11744
rect 2136 11698 2188 11704
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 9178 1992 10542
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2056 8634 2084 9454
rect 2148 9364 2176 11698
rect 2240 10266 2268 12679
rect 2318 12336 2374 12345
rect 2318 12271 2374 12280
rect 2332 11150 2360 12271
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2424 10810 2452 13194
rect 2964 12640 3016 12646
rect 2778 12608 2834 12617
rect 2964 12582 3016 12588
rect 2778 12543 2834 12552
rect 2792 12442 2820 12543
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2596 12164 2648 12170
rect 2596 12106 2648 12112
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2516 11898 2544 12038
rect 2608 11898 2636 12106
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2504 11756 2556 11762
rect 2556 11716 2636 11744
rect 2504 11698 2556 11704
rect 2502 11656 2558 11665
rect 2502 11591 2558 11600
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2424 10674 2452 10746
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2240 10062 2268 10202
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2318 10024 2374 10033
rect 2318 9959 2374 9968
rect 2228 9376 2280 9382
rect 2148 9336 2228 9364
rect 2228 9318 2280 9324
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 1952 8560 2004 8566
rect 1950 8528 1952 8537
rect 2004 8528 2006 8537
rect 2006 8486 2084 8514
rect 1950 8463 2006 8472
rect 1872 8350 1992 8378
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1872 5710 1900 8230
rect 1964 5778 1992 8350
rect 2056 6712 2084 8486
rect 2148 7886 2176 8570
rect 2240 8362 2268 9318
rect 2332 9042 2360 9959
rect 2424 9722 2452 10406
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2332 8498 2360 8978
rect 2516 8514 2544 11591
rect 2608 11014 2636 11716
rect 2700 11218 2728 12242
rect 2792 11354 2820 12378
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2884 11121 2912 12038
rect 2976 11898 3004 12582
rect 3068 12434 3096 15166
rect 3174 14716 3482 14725
rect 3174 14714 3180 14716
rect 3236 14714 3260 14716
rect 3316 14714 3340 14716
rect 3396 14714 3420 14716
rect 3476 14714 3482 14716
rect 3236 14662 3238 14714
rect 3418 14662 3420 14714
rect 3174 14660 3180 14662
rect 3236 14660 3260 14662
rect 3316 14660 3340 14662
rect 3396 14660 3420 14662
rect 3476 14660 3482 14662
rect 3174 14651 3482 14660
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3436 13841 3464 14350
rect 3620 14346 3648 16510
rect 3974 16280 4030 16289
rect 3974 16215 4030 16224
rect 3988 15230 4016 16215
rect 4066 15872 4122 15881
rect 4066 15807 4122 15816
rect 3976 15224 4028 15230
rect 4080 15212 4108 15807
rect 4080 15184 4200 15212
rect 3976 15166 4028 15172
rect 4172 14618 4200 15184
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3514 14240 3570 14249
rect 3514 14175 3570 14184
rect 3528 14006 3556 14175
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3422 13832 3478 13841
rect 3422 13767 3478 13776
rect 3174 13628 3482 13637
rect 3174 13626 3180 13628
rect 3236 13626 3260 13628
rect 3316 13626 3340 13628
rect 3396 13626 3420 13628
rect 3476 13626 3482 13628
rect 3236 13574 3238 13626
rect 3418 13574 3420 13626
rect 3174 13572 3180 13574
rect 3236 13572 3260 13574
rect 3316 13572 3340 13574
rect 3396 13572 3420 13574
rect 3476 13572 3482 13574
rect 3174 13563 3482 13572
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3174 12540 3482 12549
rect 3174 12538 3180 12540
rect 3236 12538 3260 12540
rect 3316 12538 3340 12540
rect 3396 12538 3420 12540
rect 3476 12538 3482 12540
rect 3236 12486 3238 12538
rect 3418 12486 3420 12538
rect 3174 12484 3180 12486
rect 3236 12484 3260 12486
rect 3316 12484 3340 12486
rect 3396 12484 3420 12486
rect 3476 12484 3482 12486
rect 3174 12475 3482 12484
rect 3068 12406 3188 12434
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3160 11778 3188 12406
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3238 12200 3294 12209
rect 3238 12135 3294 12144
rect 2976 11750 3188 11778
rect 2870 11112 2926 11121
rect 2688 11076 2740 11082
rect 2870 11047 2926 11056
rect 2688 11018 2740 11024
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2700 10810 2728 11018
rect 2872 11008 2924 11014
rect 2778 10976 2834 10985
rect 2872 10950 2924 10956
rect 2778 10911 2834 10920
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2424 8486 2544 8514
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2226 8120 2282 8129
rect 2226 8055 2228 8064
rect 2280 8055 2282 8064
rect 2228 8026 2280 8032
rect 2424 7936 2452 8486
rect 2332 7908 2452 7936
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 7721 2268 7822
rect 2226 7712 2282 7721
rect 2226 7647 2282 7656
rect 2226 7440 2282 7449
rect 2136 7404 2188 7410
rect 2332 7426 2360 7908
rect 2608 7585 2636 8978
rect 2700 8430 2728 10610
rect 2792 10266 2820 10911
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2778 9752 2834 9761
rect 2778 9687 2834 9696
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2700 8022 2728 8366
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2594 7576 2650 7585
rect 2594 7511 2650 7520
rect 2700 7460 2728 7686
rect 2608 7432 2728 7460
rect 2332 7398 2452 7426
rect 2226 7375 2282 7384
rect 2136 7346 2188 7352
rect 2148 6866 2176 7346
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2056 6684 2176 6712
rect 2042 6624 2098 6633
rect 2042 6559 2098 6568
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1860 5704 1912 5710
rect 1766 5672 1822 5681
rect 1912 5652 1992 5658
rect 1860 5646 1992 5652
rect 1872 5630 1992 5646
rect 1766 5607 1822 5616
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1674 4040 1730 4049
rect 1674 3975 1730 3984
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1490 3224 1546 3233
rect 1490 3159 1546 3168
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1504 1601 1532 2790
rect 1688 2417 1716 3878
rect 1674 2408 1730 2417
rect 1674 2343 1730 2352
rect 1780 2009 1808 5510
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1872 3641 1900 4966
rect 1964 4826 1992 5630
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2056 4146 2084 6559
rect 2148 6254 2176 6684
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2240 5234 2268 7375
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2332 7002 2360 7278
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2332 6798 2360 6938
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2424 6610 2452 7398
rect 2504 7200 2556 7206
rect 2608 7177 2636 7432
rect 2792 7392 2820 9687
rect 2884 9586 2912 10950
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2884 9450 2912 9522
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2884 9353 2912 9386
rect 2870 9344 2926 9353
rect 2870 9279 2926 9288
rect 2700 7364 2820 7392
rect 2504 7142 2556 7148
rect 2594 7168 2650 7177
rect 2516 6934 2544 7142
rect 2594 7103 2650 7112
rect 2594 7032 2650 7041
rect 2594 6967 2596 6976
rect 2648 6967 2650 6976
rect 2596 6938 2648 6944
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2594 6760 2650 6769
rect 2594 6695 2650 6704
rect 2424 6582 2544 6610
rect 2410 6488 2466 6497
rect 2410 6423 2466 6432
rect 2424 6322 2452 6423
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2228 5228 2280 5234
rect 2332 5216 2360 6190
rect 2424 5914 2452 6258
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2516 5234 2544 6582
rect 2504 5228 2556 5234
rect 2332 5188 2452 5216
rect 2228 5170 2280 5176
rect 2240 5114 2268 5170
rect 2240 5086 2360 5114
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2134 4720 2190 4729
rect 2134 4655 2136 4664
rect 2188 4655 2190 4664
rect 2136 4626 2188 4632
rect 2240 4457 2268 4966
rect 2226 4448 2282 4457
rect 2226 4383 2282 4392
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1858 3632 1914 3641
rect 1858 3567 1914 3576
rect 1964 2825 1992 3878
rect 2332 3738 2360 5086
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2424 3602 2452 5188
rect 2504 5170 2556 5176
rect 2516 3670 2544 5170
rect 2608 4146 2636 6695
rect 2700 6662 2728 7364
rect 2884 7324 2912 9279
rect 2976 9178 3004 11750
rect 3252 11642 3280 12135
rect 3344 11830 3372 12242
rect 3528 12238 3556 12582
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3332 11824 3384 11830
rect 3332 11766 3384 11772
rect 3068 11614 3280 11642
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3068 11257 3096 11614
rect 3174 11452 3482 11461
rect 3174 11450 3180 11452
rect 3236 11450 3260 11452
rect 3316 11450 3340 11452
rect 3396 11450 3420 11452
rect 3476 11450 3482 11452
rect 3236 11398 3238 11450
rect 3418 11398 3420 11450
rect 3174 11396 3180 11398
rect 3236 11396 3260 11398
rect 3316 11396 3340 11398
rect 3396 11396 3420 11398
rect 3476 11396 3482 11398
rect 3174 11387 3482 11396
rect 3054 11248 3110 11257
rect 3054 11183 3110 11192
rect 3068 10810 3096 11183
rect 3422 10976 3478 10985
rect 3422 10911 3478 10920
rect 3436 10810 3464 10911
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3436 10674 3464 10746
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3528 10606 3556 11630
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3174 10364 3482 10373
rect 3174 10362 3180 10364
rect 3236 10362 3260 10364
rect 3316 10362 3340 10364
rect 3396 10362 3420 10364
rect 3476 10362 3482 10364
rect 3236 10310 3238 10362
rect 3418 10310 3420 10362
rect 3174 10308 3180 10310
rect 3236 10308 3260 10310
rect 3316 10308 3340 10310
rect 3396 10308 3420 10310
rect 3476 10308 3482 10310
rect 3174 10299 3482 10308
rect 3054 10160 3110 10169
rect 3054 10095 3056 10104
rect 3108 10095 3110 10104
rect 3056 10066 3108 10072
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2964 8832 3016 8838
rect 2962 8800 2964 8809
rect 3016 8800 3018 8809
rect 2962 8735 3018 8744
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2792 7296 2912 7324
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2686 6352 2742 6361
rect 2686 6287 2742 6296
rect 2700 5166 2728 6287
rect 2792 5778 2820 7296
rect 2976 7274 3004 8434
rect 3068 7546 3096 10066
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3160 9489 3188 9590
rect 3146 9480 3202 9489
rect 3528 9466 3556 10542
rect 3620 9654 3648 14010
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4158 13424 4214 13433
rect 4158 13359 4214 13368
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3712 11558 3740 12174
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4080 11898 4108 12038
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4066 11792 4122 11801
rect 4172 11762 4200 13359
rect 4264 13258 4292 13874
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4252 13252 4304 13258
rect 4252 13194 4304 13200
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4066 11727 4122 11736
rect 4160 11756 4212 11762
rect 3700 11552 3752 11558
rect 3884 11552 3936 11558
rect 3700 11494 3752 11500
rect 3882 11520 3884 11529
rect 3976 11552 4028 11558
rect 3936 11520 3938 11529
rect 3976 11494 4028 11500
rect 3882 11455 3938 11464
rect 3884 10532 3936 10538
rect 3884 10474 3936 10480
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3712 9761 3740 10134
rect 3698 9752 3754 9761
rect 3698 9687 3754 9696
rect 3608 9648 3660 9654
rect 3608 9590 3660 9596
rect 3528 9438 3648 9466
rect 3146 9415 3202 9424
rect 3174 9276 3482 9285
rect 3174 9274 3180 9276
rect 3236 9274 3260 9276
rect 3316 9274 3340 9276
rect 3396 9274 3420 9276
rect 3476 9274 3482 9276
rect 3236 9222 3238 9274
rect 3418 9222 3420 9274
rect 3174 9220 3180 9222
rect 3236 9220 3260 9222
rect 3316 9220 3340 9222
rect 3396 9220 3420 9222
rect 3476 9220 3482 9222
rect 3174 9211 3482 9220
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3160 8634 3188 8910
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3424 8424 3476 8430
rect 3422 8392 3424 8401
rect 3476 8392 3478 8401
rect 3422 8327 3478 8336
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 3174 8188 3482 8197
rect 3174 8186 3180 8188
rect 3236 8186 3260 8188
rect 3316 8186 3340 8188
rect 3396 8186 3420 8188
rect 3476 8186 3482 8188
rect 3236 8134 3238 8186
rect 3418 8134 3420 8186
rect 3174 8132 3180 8134
rect 3236 8132 3260 8134
rect 3316 8132 3340 8134
rect 3396 8132 3420 8134
rect 3476 8132 3482 8134
rect 3174 8123 3482 8132
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3332 8016 3384 8022
rect 3436 7993 3464 8026
rect 3332 7958 3384 7964
rect 3422 7984 3478 7993
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3160 7410 3188 7890
rect 3344 7886 3372 7958
rect 3422 7919 3478 7928
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3436 7818 3464 7919
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3344 7313 3372 7686
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3436 7449 3464 7482
rect 3422 7440 3478 7449
rect 3422 7375 3478 7384
rect 3330 7304 3386 7313
rect 2964 7268 3016 7274
rect 3330 7239 3386 7248
rect 2964 7210 3016 7216
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 2962 7032 3018 7041
rect 2872 6996 2924 7002
rect 3068 7002 3096 7142
rect 3174 7100 3482 7109
rect 3174 7098 3180 7100
rect 3236 7098 3260 7100
rect 3316 7098 3340 7100
rect 3396 7098 3420 7100
rect 3476 7098 3482 7100
rect 3236 7046 3238 7098
rect 3418 7046 3420 7098
rect 3174 7044 3180 7046
rect 3236 7044 3260 7046
rect 3316 7044 3340 7046
rect 3396 7044 3420 7046
rect 3476 7044 3482 7046
rect 3174 7035 3482 7044
rect 2962 6967 3018 6976
rect 3056 6996 3108 7002
rect 2872 6938 2924 6944
rect 2884 5914 2912 6938
rect 2976 6848 3004 6967
rect 3056 6938 3108 6944
rect 3056 6860 3108 6866
rect 2976 6820 3056 6848
rect 3056 6802 3108 6808
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 6186 3096 6598
rect 3424 6248 3476 6254
rect 3422 6216 3424 6225
rect 3476 6216 3478 6225
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 3056 6180 3108 6186
rect 3422 6151 3478 6160
rect 3056 6122 3108 6128
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2792 5370 2820 5714
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2504 3664 2556 3670
rect 2504 3606 2556 3612
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2044 3460 2096 3466
rect 2044 3402 2096 3408
rect 1950 2816 2006 2825
rect 1950 2751 2006 2760
rect 1766 2000 1822 2009
rect 1766 1935 1822 1944
rect 1490 1592 1546 1601
rect 1490 1527 1546 1536
rect 1398 1184 1454 1193
rect 1398 1119 1454 1128
rect 2056 800 2084 3402
rect 2424 3126 2452 3538
rect 2608 3126 2636 3606
rect 2412 3120 2464 3126
rect 2412 3062 2464 3068
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2700 2650 2728 5102
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4690 2820 4966
rect 2884 4826 2912 5102
rect 2976 4865 3004 6122
rect 3068 5234 3096 6122
rect 3174 6012 3482 6021
rect 3174 6010 3180 6012
rect 3236 6010 3260 6012
rect 3316 6010 3340 6012
rect 3396 6010 3420 6012
rect 3476 6010 3482 6012
rect 3236 5958 3238 6010
rect 3418 5958 3420 6010
rect 3174 5956 3180 5958
rect 3236 5956 3260 5958
rect 3316 5956 3340 5958
rect 3396 5956 3420 5958
rect 3476 5956 3482 5958
rect 3174 5947 3482 5956
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2962 4856 3018 4865
rect 2872 4820 2924 4826
rect 2962 4791 3018 4800
rect 2872 4762 2924 4768
rect 3068 4758 3096 5170
rect 3174 4924 3482 4933
rect 3174 4922 3180 4924
rect 3236 4922 3260 4924
rect 3316 4922 3340 4924
rect 3396 4922 3420 4924
rect 3476 4922 3482 4924
rect 3236 4870 3238 4922
rect 3418 4870 3420 4922
rect 3174 4868 3180 4870
rect 3236 4868 3260 4870
rect 3316 4868 3340 4870
rect 3396 4868 3420 4870
rect 3476 4868 3482 4870
rect 3174 4859 3482 4868
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 3240 4548 3292 4554
rect 3240 4490 3292 4496
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 2792 3534 2820 4111
rect 2976 3670 3004 4490
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 3068 3602 3096 4422
rect 3252 4282 3280 4490
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3436 4214 3464 4694
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3174 3836 3482 3845
rect 3174 3834 3180 3836
rect 3236 3834 3260 3836
rect 3316 3834 3340 3836
rect 3396 3834 3420 3836
rect 3476 3834 3482 3836
rect 3236 3782 3238 3834
rect 3418 3782 3420 3834
rect 3174 3780 3180 3782
rect 3236 3780 3260 3782
rect 3316 3780 3340 3782
rect 3396 3780 3420 3782
rect 3476 3780 3482 3782
rect 3174 3771 3482 3780
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3528 3534 3556 8298
rect 3620 8265 3648 9438
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3606 8256 3662 8265
rect 3606 8191 3662 8200
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3620 6798 3648 7414
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 6458 3648 6598
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3620 5914 3648 6258
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3620 5710 3648 5850
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3606 3496 3662 3505
rect 3056 3460 3108 3466
rect 3606 3431 3662 3440
rect 3056 3402 3108 3408
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2502 2544 2558 2553
rect 2502 2479 2558 2488
rect 2780 2508 2832 2514
rect 2516 2446 2544 2479
rect 2780 2450 2832 2456
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 1214 0 1270 800
rect 2042 0 2098 800
rect 2792 377 2820 2450
rect 2884 800 2912 2858
rect 3068 2650 3096 3402
rect 3330 3088 3386 3097
rect 3620 3058 3648 3431
rect 3712 3194 3740 9318
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3804 8634 3832 8774
rect 3896 8634 3924 10474
rect 3988 9110 4016 11494
rect 4080 10985 4108 11727
rect 4160 11698 4212 11704
rect 4264 11354 4292 12038
rect 4356 11778 4384 13738
rect 4448 12102 4476 16623
rect 5538 16400 5594 17200
rect 7746 16538 7802 17200
rect 9954 16538 10010 17200
rect 12162 16538 12218 17200
rect 7746 16510 8064 16538
rect 7746 16400 7802 16510
rect 5552 14278 5580 16400
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5000 13870 5028 14214
rect 5398 14172 5706 14181
rect 5398 14170 5404 14172
rect 5460 14170 5484 14172
rect 5540 14170 5564 14172
rect 5620 14170 5644 14172
rect 5700 14170 5706 14172
rect 5460 14118 5462 14170
rect 5642 14118 5644 14170
rect 5398 14116 5404 14118
rect 5460 14116 5484 14118
rect 5540 14116 5564 14118
rect 5620 14116 5644 14118
rect 5700 14116 5706 14118
rect 5398 14107 5706 14116
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4632 13530 4660 13806
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 5092 13274 5120 14010
rect 5736 13802 5764 14554
rect 5908 14000 5960 14006
rect 6092 14000 6144 14006
rect 5960 13948 6092 13954
rect 5908 13942 6144 13948
rect 5920 13926 6132 13942
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 4632 13246 5120 13274
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4540 12986 4568 13126
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4540 11898 4568 12106
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4356 11750 4476 11778
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4066 10976 4122 10985
rect 4066 10911 4122 10920
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 4080 9761 4108 10678
rect 4066 9752 4122 9761
rect 4066 9687 4122 9696
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3974 8936 4030 8945
rect 3974 8871 4030 8880
rect 3988 8838 4016 8871
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3988 8480 4016 8774
rect 3896 8452 4016 8480
rect 3790 7576 3846 7585
rect 3896 7546 3924 8452
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3790 7511 3846 7520
rect 3884 7540 3936 7546
rect 3804 7274 3832 7511
rect 3884 7482 3936 7488
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3804 6225 3832 7210
rect 3896 7002 3924 7482
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3896 6254 3924 6938
rect 3884 6248 3936 6254
rect 3790 6216 3846 6225
rect 3884 6190 3936 6196
rect 3790 6151 3846 6160
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3330 3023 3332 3032
rect 3384 3023 3386 3032
rect 3608 3052 3660 3058
rect 3332 2994 3384 3000
rect 3608 2994 3660 3000
rect 3174 2748 3482 2757
rect 3174 2746 3180 2748
rect 3236 2746 3260 2748
rect 3316 2746 3340 2748
rect 3396 2746 3420 2748
rect 3476 2746 3482 2748
rect 3236 2694 3238 2746
rect 3418 2694 3420 2746
rect 3174 2692 3180 2694
rect 3236 2692 3260 2694
rect 3316 2692 3340 2694
rect 3396 2692 3420 2694
rect 3476 2692 3482 2694
rect 3174 2683 3482 2692
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3804 2446 3832 4966
rect 3896 2514 3924 6054
rect 3988 5370 4016 8298
rect 4080 7002 4108 9454
rect 4172 9450 4200 11086
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10266 4292 10950
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4356 9722 4384 11562
rect 4448 11014 4476 11750
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4540 10810 4568 11630
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4448 10130 4476 10542
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4344 9716 4396 9722
rect 4264 9664 4344 9674
rect 4264 9658 4396 9664
rect 4264 9646 4384 9658
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4264 8566 4292 9646
rect 4448 9602 4476 10066
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4540 9654 4568 9930
rect 4356 9574 4476 9602
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4356 9518 4384 9574
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4356 8514 4384 9454
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8634 4476 8774
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4356 8486 4476 8514
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4066 6896 4122 6905
rect 4066 6831 4122 6840
rect 4080 6798 4108 6831
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 4080 4758 4108 6190
rect 4172 5778 4200 7890
rect 4264 7886 4292 8366
rect 4448 8362 4476 8486
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4356 8090 4384 8298
rect 4434 8256 4490 8265
rect 4434 8191 4490 8200
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4252 7744 4304 7750
rect 4250 7712 4252 7721
rect 4304 7712 4306 7721
rect 4250 7647 4306 7656
rect 4264 7410 4292 7647
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4172 5302 4200 5714
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4068 4752 4120 4758
rect 4120 4712 4200 4740
rect 4068 4694 4120 4700
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 3712 800 3740 2314
rect 2778 368 2834 377
rect 2778 303 2834 312
rect 2870 0 2926 800
rect 3698 0 3754 800
rect 4080 785 4108 4422
rect 4172 4214 4200 4712
rect 4264 4622 4292 7210
rect 4356 6934 4384 7278
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 4344 6792 4396 6798
rect 4342 6760 4344 6769
rect 4396 6760 4398 6769
rect 4342 6695 4398 6704
rect 4448 6322 4476 8191
rect 4540 7954 4568 8978
rect 4632 8974 4660 13246
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4724 12306 4752 12718
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4724 10810 4752 12242
rect 4908 12238 4936 12854
rect 5000 12850 5028 13126
rect 5092 12986 5120 13126
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4896 12232 4948 12238
rect 4802 12200 4858 12209
rect 4896 12174 4948 12180
rect 4986 12200 5042 12209
rect 4802 12135 4804 12144
rect 4856 12135 4858 12144
rect 4986 12135 5042 12144
rect 4804 12106 4856 12112
rect 5000 12102 5028 12135
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 11898 5028 12038
rect 4804 11892 4856 11898
rect 4988 11892 5040 11898
rect 4856 11852 4936 11880
rect 4804 11834 4856 11840
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4816 11082 4844 11630
rect 4908 11218 4936 11852
rect 4988 11834 5040 11840
rect 5184 11694 5212 13330
rect 5736 13326 5764 13738
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5398 13084 5706 13093
rect 5398 13082 5404 13084
rect 5460 13082 5484 13084
rect 5540 13082 5564 13084
rect 5620 13082 5644 13084
rect 5700 13082 5706 13084
rect 5460 13030 5462 13082
rect 5642 13030 5644 13082
rect 5398 13028 5404 13030
rect 5460 13028 5484 13030
rect 5540 13028 5564 13030
rect 5620 13028 5644 13030
rect 5700 13028 5706 13030
rect 5398 13019 5706 13028
rect 5828 12986 5856 13466
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5828 12481 5856 12922
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5814 12472 5870 12481
rect 5814 12407 5870 12416
rect 5920 12238 5948 12582
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5276 11898 5304 12038
rect 5398 11996 5706 12005
rect 5398 11994 5404 11996
rect 5460 11994 5484 11996
rect 5540 11994 5564 11996
rect 5620 11994 5644 11996
rect 5700 11994 5706 11996
rect 5460 11942 5462 11994
rect 5642 11942 5644 11994
rect 5398 11940 5404 11942
rect 5460 11940 5484 11942
rect 5540 11940 5564 11942
rect 5620 11940 5644 11942
rect 5700 11940 5706 11942
rect 5398 11931 5706 11940
rect 5736 11898 5764 12038
rect 5828 11898 5856 12038
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5080 11620 5132 11626
rect 5080 11562 5132 11568
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4710 10704 4766 10713
rect 4710 10639 4712 10648
rect 4764 10639 4766 10648
rect 4712 10610 4764 10616
rect 4710 10432 4766 10441
rect 4710 10367 4766 10376
rect 4724 9110 4752 10367
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4526 7576 4582 7585
rect 4526 7511 4582 7520
rect 4540 7478 4568 7511
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4632 7324 4660 8502
rect 4540 7296 4660 7324
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4540 6186 4568 7296
rect 4618 6896 4674 6905
rect 4618 6831 4674 6840
rect 4632 6458 4660 6831
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 4632 5914 4660 6190
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4724 5794 4752 9046
rect 4816 8378 4844 11018
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4908 10169 4936 10746
rect 4894 10160 4950 10169
rect 4894 10095 4950 10104
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4908 9450 4936 9998
rect 5000 9489 5028 10950
rect 5092 10810 5120 11562
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5184 10062 5212 11222
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5276 10130 5304 10950
rect 5398 10908 5706 10917
rect 5398 10906 5404 10908
rect 5460 10906 5484 10908
rect 5540 10906 5564 10908
rect 5620 10906 5644 10908
rect 5700 10906 5706 10908
rect 5460 10854 5462 10906
rect 5642 10854 5644 10906
rect 5398 10852 5404 10854
rect 5460 10852 5484 10854
rect 5540 10852 5564 10854
rect 5620 10852 5644 10854
rect 5700 10852 5706 10854
rect 5398 10843 5706 10852
rect 5736 10810 5764 11698
rect 5920 11642 5948 12174
rect 5828 11626 5948 11642
rect 5816 11620 5948 11626
rect 5868 11614 5948 11620
rect 5816 11562 5868 11568
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5356 10600 5408 10606
rect 5354 10568 5356 10577
rect 5408 10568 5410 10577
rect 5354 10503 5410 10512
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 10305 5580 10406
rect 5538 10296 5594 10305
rect 5538 10231 5594 10240
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5172 10056 5224 10062
rect 5460 10033 5488 10066
rect 5172 9998 5224 10004
rect 5446 10024 5502 10033
rect 5552 9994 5580 10231
rect 5644 10062 5672 10746
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5446 9959 5502 9968
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5092 9586 5120 9862
rect 5398 9820 5706 9829
rect 5398 9818 5404 9820
rect 5460 9818 5484 9820
rect 5540 9818 5564 9820
rect 5620 9818 5644 9820
rect 5700 9818 5706 9820
rect 5460 9766 5462 9818
rect 5642 9766 5644 9818
rect 5398 9764 5404 9766
rect 5460 9764 5484 9766
rect 5540 9764 5564 9766
rect 5620 9764 5644 9766
rect 5700 9764 5706 9766
rect 5398 9755 5706 9764
rect 5736 9722 5764 9862
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5828 9654 5856 10202
rect 5920 9654 5948 11494
rect 6012 10674 6040 13670
rect 6288 13530 6316 15302
rect 7012 15224 7064 15230
rect 7012 15166 7064 15172
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6472 13274 6500 14010
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6276 13252 6328 13258
rect 6276 13194 6328 13200
rect 6380 13246 6500 13274
rect 6644 13320 6696 13326
rect 6748 13308 6776 13670
rect 6840 13326 6868 13738
rect 6696 13280 6776 13308
rect 6644 13262 6696 13268
rect 6288 12986 6316 13194
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6288 12073 6316 12106
rect 6274 12064 6330 12073
rect 6274 11999 6330 12008
rect 6380 11830 6408 13246
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6656 12986 6684 13126
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6748 12918 6776 13280
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 7024 12850 7052 15166
rect 7622 14716 7930 14725
rect 7622 14714 7628 14716
rect 7684 14714 7708 14716
rect 7764 14714 7788 14716
rect 7844 14714 7868 14716
rect 7924 14714 7930 14716
rect 7684 14662 7686 14714
rect 7866 14662 7868 14714
rect 7622 14660 7628 14662
rect 7684 14660 7708 14662
rect 7764 14660 7788 14662
rect 7844 14660 7868 14662
rect 7924 14660 7930 14662
rect 7622 14651 7930 14660
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7024 12646 7052 12786
rect 6828 12640 6880 12646
rect 7012 12640 7064 12646
rect 6880 12588 6960 12594
rect 6828 12582 6960 12588
rect 7012 12582 7064 12588
rect 6840 12566 6960 12582
rect 6932 12374 6960 12566
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6092 11824 6144 11830
rect 6368 11824 6420 11830
rect 6092 11766 6144 11772
rect 6366 11792 6368 11801
rect 6420 11792 6422 11801
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6012 9722 6040 9998
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4986 9480 5042 9489
rect 4896 9444 4948 9450
rect 4986 9415 5042 9424
rect 5448 9444 5500 9450
rect 4896 9386 4948 9392
rect 5448 9386 5500 9392
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5000 8838 5028 9114
rect 4988 8832 5040 8838
rect 5080 8832 5132 8838
rect 4988 8774 5040 8780
rect 5078 8800 5080 8809
rect 5132 8800 5134 8809
rect 5000 8673 5028 8774
rect 5078 8735 5134 8744
rect 4986 8664 5042 8673
rect 4986 8599 5042 8608
rect 4896 8492 4948 8498
rect 4948 8452 5028 8480
rect 4896 8434 4948 8440
rect 4816 8350 4936 8378
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4816 6905 4844 7482
rect 4802 6896 4858 6905
rect 4802 6831 4858 6840
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4816 6254 4844 6666
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4632 5766 4752 5794
rect 4434 5672 4490 5681
rect 4434 5607 4436 5616
rect 4488 5607 4490 5616
rect 4436 5578 4488 5584
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4540 5234 4568 5510
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4356 5030 4384 5170
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4356 4826 4384 4966
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4282 4292 4558
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 4160 4072 4212 4078
rect 4158 4040 4160 4049
rect 4212 4040 4214 4049
rect 4158 3975 4214 3984
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4264 3194 4292 3878
rect 4356 3194 4384 4762
rect 4448 4146 4476 5102
rect 4528 5092 4580 5098
rect 4632 5080 4660 5766
rect 4712 5704 4764 5710
rect 4816 5658 4844 6190
rect 4764 5652 4844 5658
rect 4712 5646 4844 5652
rect 4724 5630 4844 5646
rect 4816 5370 4844 5630
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4580 5052 4660 5080
rect 4528 5034 4580 5040
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4540 3602 4568 5034
rect 4724 4554 4752 5238
rect 4816 4554 4844 5306
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4632 3466 4660 3946
rect 4724 3670 4752 4490
rect 4816 4078 4844 4490
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4816 3738 4844 4014
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4172 2514 4200 2926
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4356 2446 4384 3130
rect 4448 2446 4476 3402
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4528 2916 4580 2922
rect 4528 2858 4580 2864
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 4540 800 4568 2858
rect 4724 2446 4752 3334
rect 4908 2922 4936 8350
rect 5000 5166 5028 8452
rect 5184 7954 5212 9318
rect 5460 8974 5488 9386
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5448 8968 5500 8974
rect 5552 8945 5580 8978
rect 5448 8910 5500 8916
rect 5538 8936 5594 8945
rect 5644 8906 5672 9386
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5998 9072 6054 9081
rect 5814 8936 5870 8945
rect 5538 8871 5594 8880
rect 5632 8900 5684 8906
rect 5814 8871 5816 8880
rect 5632 8842 5684 8848
rect 5868 8871 5870 8880
rect 5816 8842 5868 8848
rect 5724 8832 5776 8838
rect 5920 8809 5948 9046
rect 5998 9007 6054 9016
rect 5724 8774 5776 8780
rect 5906 8800 5962 8809
rect 5398 8732 5706 8741
rect 5398 8730 5404 8732
rect 5460 8730 5484 8732
rect 5540 8730 5564 8732
rect 5620 8730 5644 8732
rect 5700 8730 5706 8732
rect 5460 8678 5462 8730
rect 5642 8678 5644 8730
rect 5398 8676 5404 8678
rect 5460 8676 5484 8678
rect 5540 8676 5564 8678
rect 5620 8676 5644 8678
rect 5700 8676 5706 8678
rect 5398 8667 5706 8676
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5276 7818 5304 8570
rect 5736 8090 5764 8774
rect 5906 8735 5962 8744
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5632 8016 5684 8022
rect 5630 7984 5632 7993
rect 5684 7984 5686 7993
rect 5686 7942 5764 7970
rect 5630 7919 5686 7928
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5092 6730 5120 7754
rect 5398 7644 5706 7653
rect 5398 7642 5404 7644
rect 5460 7642 5484 7644
rect 5540 7642 5564 7644
rect 5620 7642 5644 7644
rect 5700 7642 5706 7644
rect 5460 7590 5462 7642
rect 5642 7590 5644 7642
rect 5398 7588 5404 7590
rect 5460 7588 5484 7590
rect 5540 7588 5564 7590
rect 5620 7588 5644 7590
rect 5700 7588 5706 7590
rect 5398 7579 5706 7588
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5184 7449 5212 7482
rect 5170 7440 5226 7449
rect 5170 7375 5226 7384
rect 5276 7206 5304 7482
rect 5630 7440 5686 7449
rect 5630 7375 5632 7384
rect 5684 7375 5686 7384
rect 5632 7346 5684 7352
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5630 7168 5686 7177
rect 5552 7041 5580 7142
rect 5630 7103 5686 7112
rect 5538 7032 5594 7041
rect 5538 6967 5594 6976
rect 5644 6934 5672 7103
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 5736 6662 5764 7942
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5398 6556 5706 6565
rect 5398 6554 5404 6556
rect 5460 6554 5484 6556
rect 5540 6554 5564 6556
rect 5620 6554 5644 6556
rect 5700 6554 5706 6556
rect 5460 6502 5462 6554
rect 5642 6502 5644 6554
rect 5398 6500 5404 6502
rect 5460 6500 5484 6502
rect 5540 6500 5564 6502
rect 5620 6500 5644 6502
rect 5700 6500 5706 6502
rect 5398 6491 5706 6500
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 5398 5468 5706 5477
rect 5398 5466 5404 5468
rect 5460 5466 5484 5468
rect 5540 5466 5564 5468
rect 5620 5466 5644 5468
rect 5700 5466 5706 5468
rect 5460 5414 5462 5466
rect 5642 5414 5644 5466
rect 5398 5412 5404 5414
rect 5460 5412 5484 5414
rect 5540 5412 5564 5414
rect 5620 5412 5644 5414
rect 5700 5412 5706 5414
rect 5398 5403 5706 5412
rect 5736 5250 5764 6326
rect 5828 5846 5856 8434
rect 5920 7750 5948 8502
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5920 7342 5948 7686
rect 6012 7478 6040 9007
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5920 7206 5948 7278
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5920 6798 5948 7142
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6012 6610 6040 6734
rect 5920 6582 6040 6610
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 5920 5642 5948 6582
rect 6104 6474 6132 11766
rect 6366 11727 6422 11736
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6196 11218 6224 11290
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6196 9110 6224 11154
rect 6380 10198 6408 11630
rect 6472 11121 6500 12038
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6458 11112 6514 11121
rect 6458 11047 6514 11056
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6288 9761 6316 10066
rect 6274 9752 6330 9761
rect 6274 9687 6330 9696
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6012 6446 6132 6474
rect 6012 6186 6040 6446
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 6104 5846 6132 6258
rect 6092 5840 6144 5846
rect 6092 5782 6144 5788
rect 6090 5672 6146 5681
rect 5908 5636 5960 5642
rect 6090 5607 6146 5616
rect 5908 5578 5960 5584
rect 5644 5234 5764 5250
rect 5632 5228 5764 5234
rect 5684 5222 5764 5228
rect 5632 5170 5684 5176
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5000 4842 5028 5102
rect 5644 5030 5672 5170
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5000 4826 5120 4842
rect 5000 4820 5132 4826
rect 5000 4814 5080 4820
rect 5080 4762 5132 4768
rect 5398 4380 5706 4389
rect 5398 4378 5404 4380
rect 5460 4378 5484 4380
rect 5540 4378 5564 4380
rect 5620 4378 5644 4380
rect 5700 4378 5706 4380
rect 5460 4326 5462 4378
rect 5642 4326 5644 4378
rect 5398 4324 5404 4326
rect 5460 4324 5484 4326
rect 5540 4324 5564 4326
rect 5620 4324 5644 4326
rect 5700 4324 5706 4326
rect 5398 4315 5706 4324
rect 5736 3942 5764 5102
rect 5920 4758 5948 5578
rect 6104 5574 6132 5607
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 6012 4486 6040 5510
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 6196 4146 6224 8774
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 6288 3505 6316 9318
rect 6380 8498 6408 10134
rect 6472 10130 6500 10950
rect 6564 10742 6592 11222
rect 6656 11218 6684 11766
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6748 11150 6776 11630
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6552 10736 6604 10742
rect 6552 10678 6604 10684
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 9722 6500 9862
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6748 9625 6776 10610
rect 6734 9616 6790 9625
rect 6734 9551 6790 9560
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6472 8430 6500 9454
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6564 8974 6592 9318
rect 6656 8974 6684 9454
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6564 8566 6592 8910
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6656 8362 6684 8910
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6748 8634 6776 8774
rect 6840 8673 6868 12310
rect 7116 12238 7144 13126
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7208 12782 7236 12922
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7392 12646 7420 14350
rect 7622 13628 7930 13637
rect 7622 13626 7628 13628
rect 7684 13626 7708 13628
rect 7764 13626 7788 13628
rect 7844 13626 7868 13628
rect 7924 13626 7930 13628
rect 7684 13574 7686 13626
rect 7866 13574 7868 13626
rect 7622 13572 7628 13574
rect 7684 13572 7708 13574
rect 7764 13572 7788 13574
rect 7844 13572 7868 13574
rect 7924 13572 7930 13574
rect 7622 13563 7930 13572
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 6932 11898 6960 12038
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6932 11218 6960 11698
rect 7116 11218 7144 12038
rect 7194 11520 7250 11529
rect 7194 11455 7250 11464
rect 7208 11354 7236 11455
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6932 9926 6960 10406
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6826 8664 6882 8673
rect 6736 8628 6788 8634
rect 6826 8599 6882 8608
rect 6736 8570 6788 8576
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5710 6408 6054
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6380 5370 6408 5646
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6472 4049 6500 5306
rect 6458 4040 6514 4049
rect 6458 3975 6514 3984
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6274 3496 6330 3505
rect 6274 3431 6330 3440
rect 5398 3292 5706 3301
rect 5398 3290 5404 3292
rect 5460 3290 5484 3292
rect 5540 3290 5564 3292
rect 5620 3290 5644 3292
rect 5700 3290 5706 3292
rect 5460 3238 5462 3290
rect 5642 3238 5644 3290
rect 5398 3236 5404 3238
rect 5460 3236 5484 3238
rect 5540 3236 5564 3238
rect 5620 3236 5644 3238
rect 5700 3236 5706 3238
rect 5398 3227 5706 3236
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4712 2440 4764 2446
rect 4816 2417 4844 2450
rect 4712 2382 4764 2388
rect 4802 2408 4858 2417
rect 4724 2038 4752 2382
rect 4802 2343 4858 2352
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 5276 1442 5304 3062
rect 5644 2514 5672 3130
rect 6090 3088 6146 3097
rect 6090 3023 6092 3032
rect 6144 3023 6146 3032
rect 6092 2994 6144 3000
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 6196 2650 6224 2926
rect 6380 2854 6408 3674
rect 6472 3466 6500 3975
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6564 3097 6592 8230
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6656 4622 6684 5170
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6656 3534 6684 4558
rect 6748 4282 6776 8298
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 7546 6868 8230
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6932 7426 6960 9590
rect 6840 7398 6960 7426
rect 6840 6361 6868 7398
rect 6918 7168 6974 7177
rect 6918 7103 6974 7112
rect 6826 6352 6882 6361
rect 6826 6287 6882 6296
rect 6932 5234 6960 7103
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 7024 4554 7052 10474
rect 7116 6798 7144 11154
rect 7300 11082 7328 12038
rect 7484 11694 7512 13330
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7576 12753 7604 12786
rect 7562 12744 7618 12753
rect 7562 12679 7618 12688
rect 7622 12540 7930 12549
rect 7622 12538 7628 12540
rect 7684 12538 7708 12540
rect 7764 12538 7788 12540
rect 7844 12538 7868 12540
rect 7924 12538 7930 12540
rect 7684 12486 7686 12538
rect 7866 12486 7868 12538
rect 7622 12484 7628 12486
rect 7684 12484 7708 12486
rect 7764 12484 7788 12486
rect 7844 12484 7868 12486
rect 7924 12484 7930 12486
rect 7622 12475 7930 12484
rect 8036 12481 8064 16510
rect 9954 16510 10272 16538
rect 9954 16400 10010 16510
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9784 14074 9812 14486
rect 9846 14172 10154 14181
rect 9846 14170 9852 14172
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 10148 14170 10154 14172
rect 9908 14118 9910 14170
rect 10090 14118 10092 14170
rect 9846 14116 9852 14118
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 10148 14116 10154 14118
rect 9846 14107 10154 14116
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 8114 13288 8170 13297
rect 8114 13223 8170 13232
rect 8128 12850 8156 13223
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 8022 12472 8078 12481
rect 8022 12407 8078 12416
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7656 12096 7708 12102
rect 7654 12064 7656 12073
rect 7748 12096 7800 12102
rect 7708 12064 7710 12073
rect 7748 12038 7800 12044
rect 7654 11999 7710 12008
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7472 11688 7524 11694
rect 7760 11665 7788 12038
rect 7852 11762 7880 12242
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7472 11630 7524 11636
rect 7746 11656 7802 11665
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7208 10441 7236 10542
rect 7194 10432 7250 10441
rect 7194 10367 7250 10376
rect 7194 10296 7250 10305
rect 7194 10231 7250 10240
rect 7208 9994 7236 10231
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7300 8838 7328 10678
rect 7392 10266 7420 11630
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7286 8664 7342 8673
rect 7286 8599 7342 8608
rect 7300 8566 7328 8599
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7300 8090 7328 8502
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7208 7002 7236 7958
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7300 7410 7328 7686
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7392 7324 7420 10066
rect 7484 7886 7512 11630
rect 7944 11626 7972 12038
rect 8036 11676 8064 12174
rect 8128 11880 8156 12582
rect 8220 12238 8248 12718
rect 9404 12368 9456 12374
rect 9456 12328 9536 12356
rect 9404 12310 9456 12316
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 9508 12102 9536 12328
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 8956 11898 8984 12038
rect 9324 11898 9352 12038
rect 9508 11898 9536 12038
rect 8208 11892 8260 11898
rect 8128 11852 8208 11880
rect 8208 11834 8260 11840
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 8116 11688 8168 11694
rect 8036 11648 8116 11676
rect 8116 11630 8168 11636
rect 7746 11591 7802 11600
rect 7932 11620 7984 11626
rect 7984 11580 8064 11608
rect 7932 11562 7984 11568
rect 7622 11452 7930 11461
rect 7622 11450 7628 11452
rect 7684 11450 7708 11452
rect 7764 11450 7788 11452
rect 7844 11450 7868 11452
rect 7924 11450 7930 11452
rect 7684 11398 7686 11450
rect 7866 11398 7868 11450
rect 7622 11396 7628 11398
rect 7684 11396 7708 11398
rect 7764 11396 7788 11398
rect 7844 11396 7868 11398
rect 7924 11396 7930 11398
rect 7622 11387 7930 11396
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7576 10810 7604 10950
rect 7668 10810 7696 11018
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10470 7604 10610
rect 7760 10606 7788 11154
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7852 10554 7880 11290
rect 8036 11268 8064 11580
rect 7944 11240 8064 11268
rect 7944 11082 7972 11240
rect 8024 11144 8076 11150
rect 8022 11112 8024 11121
rect 8076 11112 8078 11121
rect 7932 11076 7984 11082
rect 8022 11047 8078 11056
rect 7932 11018 7984 11024
rect 7852 10526 8064 10554
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7622 10364 7930 10373
rect 7622 10362 7628 10364
rect 7684 10362 7708 10364
rect 7764 10362 7788 10364
rect 7844 10362 7868 10364
rect 7924 10362 7930 10364
rect 7684 10310 7686 10362
rect 7866 10310 7868 10362
rect 7622 10308 7628 10310
rect 7684 10308 7708 10310
rect 7764 10308 7788 10310
rect 7844 10308 7868 10310
rect 7924 10308 7930 10310
rect 7622 10299 7930 10308
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7760 9926 7788 10202
rect 8036 10010 8064 10526
rect 8128 10130 8156 11630
rect 8220 10742 8248 11834
rect 9692 11762 9720 13942
rect 10244 13870 10272 16510
rect 11992 16510 12218 16538
rect 11244 15292 11296 15298
rect 11244 15234 11296 15240
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10336 14074 10364 14418
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10416 13932 10468 13938
rect 10612 13920 10640 14350
rect 10468 13892 10640 13920
rect 10416 13874 10468 13880
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 9846 13084 10154 13093
rect 9846 13082 9852 13084
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 10148 13082 10154 13084
rect 9908 13030 9910 13082
rect 10090 13030 10092 13082
rect 9846 13028 9852 13030
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 10148 13028 10154 13030
rect 9846 13019 10154 13028
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10230 12336 10286 12345
rect 10230 12271 10232 12280
rect 10284 12271 10286 12280
rect 10232 12242 10284 12248
rect 10520 12209 10548 12582
rect 10506 12200 10562 12209
rect 10506 12135 10562 12144
rect 10520 12102 10548 12135
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 9784 11830 9812 12038
rect 9846 11996 10154 12005
rect 9846 11994 9852 11996
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 10148 11994 10154 11996
rect 9908 11942 9910 11994
rect 10090 11942 10092 11994
rect 9846 11940 9852 11942
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 10148 11940 10154 11942
rect 9846 11931 10154 11940
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8312 11014 8340 11494
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8496 11014 8524 11290
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10810 8524 10950
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 10266 8248 10406
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8312 10198 8340 10610
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8404 10130 8432 10542
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8036 9982 8156 10010
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 8022 9888 8078 9897
rect 7576 9654 7604 9862
rect 7852 9722 7880 9862
rect 8022 9823 8078 9832
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7654 9616 7710 9625
rect 7576 9382 7604 9590
rect 7654 9551 7656 9560
rect 7708 9551 7710 9560
rect 7656 9522 7708 9528
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7622 9276 7930 9285
rect 7622 9274 7628 9276
rect 7684 9274 7708 9276
rect 7764 9274 7788 9276
rect 7844 9274 7868 9276
rect 7924 9274 7930 9276
rect 7684 9222 7686 9274
rect 7866 9222 7868 9274
rect 7622 9220 7628 9222
rect 7684 9220 7708 9222
rect 7764 9220 7788 9222
rect 7844 9220 7868 9222
rect 7924 9220 7930 9222
rect 7622 9211 7930 9220
rect 7562 8664 7618 8673
rect 7562 8599 7618 8608
rect 7576 8401 7604 8599
rect 7562 8392 7618 8401
rect 7562 8327 7618 8336
rect 7622 8188 7930 8197
rect 7622 8186 7628 8188
rect 7684 8186 7708 8188
rect 7764 8186 7788 8188
rect 7844 8186 7868 8188
rect 7924 8186 7930 8188
rect 7684 8134 7686 8186
rect 7866 8134 7868 8186
rect 7622 8132 7628 8134
rect 7684 8132 7708 8134
rect 7764 8132 7788 8134
rect 7844 8132 7868 8134
rect 7924 8132 7930 8134
rect 7622 8123 7930 8132
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7484 7546 7512 7822
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7372 7296 7420 7324
rect 7372 7256 7400 7296
rect 7372 7228 7420 7256
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7208 5642 7236 6938
rect 7392 6934 7420 7228
rect 7668 7188 7696 7482
rect 7484 7160 7696 7188
rect 7484 7002 7512 7160
rect 7622 7100 7930 7109
rect 7622 7098 7628 7100
rect 7684 7098 7708 7100
rect 7764 7098 7788 7100
rect 7844 7098 7868 7100
rect 7924 7098 7930 7100
rect 7684 7046 7686 7098
rect 7866 7046 7868 7098
rect 7622 7044 7628 7046
rect 7684 7044 7708 7046
rect 7764 7044 7788 7046
rect 7844 7044 7868 7046
rect 7924 7044 7930 7046
rect 7622 7035 7930 7044
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7392 6730 7420 6870
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 8036 6168 8064 9823
rect 8128 7478 8156 9982
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8312 9466 8340 9862
rect 8220 9438 8340 9466
rect 8220 8498 8248 9438
rect 8300 9376 8352 9382
rect 8298 9344 8300 9353
rect 8352 9344 8354 9353
rect 8298 9279 8354 9288
rect 8404 9178 8432 9930
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8496 8974 8524 10406
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8300 7540 8352 7546
rect 8220 7500 8300 7528
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8116 6180 8168 6186
rect 8036 6140 8116 6168
rect 8116 6122 8168 6128
rect 7622 6012 7930 6021
rect 7622 6010 7628 6012
rect 7684 6010 7708 6012
rect 7764 6010 7788 6012
rect 7844 6010 7868 6012
rect 7924 6010 7930 6012
rect 7684 5958 7686 6010
rect 7866 5958 7868 6010
rect 7622 5956 7628 5958
rect 7684 5956 7708 5958
rect 7764 5956 7788 5958
rect 7844 5956 7868 5958
rect 7924 5956 7930 5958
rect 7622 5947 7930 5956
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 8036 5098 8064 5578
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 7622 4924 7930 4933
rect 7622 4922 7628 4924
rect 7684 4922 7708 4924
rect 7764 4922 7788 4924
rect 7844 4922 7868 4924
rect 7924 4922 7930 4924
rect 7684 4870 7686 4922
rect 7866 4870 7868 4922
rect 7622 4868 7628 4870
rect 7684 4868 7708 4870
rect 7764 4868 7788 4870
rect 7844 4868 7868 4870
rect 7924 4868 7930 4870
rect 7622 4859 7930 4868
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6656 3126 6684 3470
rect 6644 3120 6696 3126
rect 6550 3088 6606 3097
rect 6644 3062 6696 3068
rect 6550 3023 6606 3032
rect 6656 2990 6684 3062
rect 6932 3058 6960 4490
rect 7024 3942 7052 4490
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 6748 2922 7052 2938
rect 6736 2916 7052 2922
rect 6788 2910 7052 2916
rect 6736 2858 6788 2864
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6458 2680 6514 2689
rect 6000 2644 6052 2650
rect 6184 2644 6236 2650
rect 6052 2604 6132 2632
rect 6000 2586 6052 2592
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5398 2204 5706 2213
rect 5398 2202 5404 2204
rect 5460 2202 5484 2204
rect 5540 2202 5564 2204
rect 5620 2202 5644 2204
rect 5700 2202 5706 2204
rect 5460 2150 5462 2202
rect 5642 2150 5644 2202
rect 5398 2148 5404 2150
rect 5460 2148 5484 2150
rect 5540 2148 5564 2150
rect 5620 2148 5644 2150
rect 5700 2148 5706 2150
rect 5398 2139 5706 2148
rect 5276 1414 5396 1442
rect 5368 800 5396 1414
rect 6104 1170 6132 2604
rect 6458 2615 6514 2624
rect 6184 2586 6236 2592
rect 6472 2446 6500 2615
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6104 1142 6224 1170
rect 6196 800 6224 1142
rect 7024 800 7052 2910
rect 7484 2650 7512 4558
rect 8036 4146 8064 4762
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7622 3836 7930 3845
rect 7622 3834 7628 3836
rect 7684 3834 7708 3836
rect 7764 3834 7788 3836
rect 7844 3834 7868 3836
rect 7924 3834 7930 3836
rect 7684 3782 7686 3834
rect 7866 3782 7868 3834
rect 7622 3780 7628 3782
rect 7684 3780 7708 3782
rect 7764 3780 7788 3782
rect 7844 3780 7868 3782
rect 7924 3780 7930 3782
rect 7622 3771 7930 3780
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 8036 2854 8064 3606
rect 8220 3466 8248 7500
rect 8300 7482 8352 7488
rect 8404 6390 8432 8502
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8128 2990 8156 3130
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 7622 2748 7930 2757
rect 7622 2746 7628 2748
rect 7684 2746 7708 2748
rect 7764 2746 7788 2748
rect 7844 2746 7868 2748
rect 7924 2746 7930 2748
rect 7684 2694 7686 2746
rect 7866 2694 7868 2746
rect 7622 2692 7628 2694
rect 7684 2692 7708 2694
rect 7764 2692 7788 2694
rect 7844 2692 7868 2694
rect 7924 2692 7930 2694
rect 7622 2683 7930 2692
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 8312 2446 8340 6054
rect 8496 4622 8524 8774
rect 8588 7546 8616 11154
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8680 10985 8708 11018
rect 8666 10976 8722 10985
rect 8666 10911 8722 10920
rect 8666 10840 8722 10849
rect 8956 10810 8984 11698
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9140 11354 9168 11630
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8666 10775 8722 10784
rect 8944 10804 8996 10810
rect 8680 10062 8708 10775
rect 8944 10746 8996 10752
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8680 9926 8708 9998
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8680 9110 8708 9454
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8680 6730 8708 9046
rect 8772 9042 8800 9318
rect 8956 9217 8984 9862
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 8942 9208 8998 9217
rect 8942 9143 8998 9152
rect 9048 9081 9076 9658
rect 9034 9072 9090 9081
rect 8760 9036 8812 9042
rect 9034 9007 9090 9016
rect 8760 8978 8812 8984
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8772 8537 8800 8774
rect 8864 8673 8892 8774
rect 8850 8664 8906 8673
rect 8850 8599 8906 8608
rect 8956 8566 8984 8842
rect 8944 8560 8996 8566
rect 8758 8528 8814 8537
rect 8944 8502 8996 8508
rect 8758 8463 8814 8472
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8864 7886 8892 8230
rect 9048 7970 9076 9007
rect 8956 7942 9076 7970
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8864 7410 8892 7822
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8956 7342 8984 7942
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8942 6760 8998 6769
rect 8668 6724 8720 6730
rect 8942 6695 8998 6704
rect 8668 6666 8720 6672
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8668 5228 8720 5234
rect 8588 5188 8668 5216
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8404 3602 8432 4014
rect 8482 3632 8538 3641
rect 8392 3596 8444 3602
rect 8482 3567 8538 3576
rect 8392 3538 8444 3544
rect 8404 2972 8432 3538
rect 8496 3534 8524 3567
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8588 3126 8616 5188
rect 8668 5170 8720 5176
rect 8864 4826 8892 6598
rect 8956 6254 8984 6695
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8864 3670 8892 4762
rect 8852 3664 8904 3670
rect 8852 3606 8904 3612
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8484 2984 8536 2990
rect 8404 2944 8484 2972
rect 8484 2926 8536 2932
rect 8496 2650 8524 2926
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8300 2440 8352 2446
rect 7930 2408 7986 2417
rect 7840 2372 7892 2378
rect 8300 2382 8352 2388
rect 7930 2343 7932 2352
rect 7840 2314 7892 2320
rect 7984 2343 7986 2352
rect 7932 2314 7984 2320
rect 7852 800 7880 2314
rect 8680 800 8708 3402
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8772 3126 8800 3334
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 9048 3058 9076 7822
rect 9140 7750 9168 11290
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 10810 9444 11018
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9416 10538 9444 10746
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9402 10160 9458 10169
rect 9312 10124 9364 10130
rect 9402 10095 9458 10104
rect 9312 10066 9364 10072
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9232 9926 9260 9998
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9220 9648 9272 9654
rect 9218 9616 9220 9625
rect 9272 9616 9274 9625
rect 9218 9551 9274 9560
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9232 9217 9260 9454
rect 9218 9208 9274 9217
rect 9218 9143 9274 9152
rect 9218 8800 9274 8809
rect 9218 8735 9274 8744
rect 9232 8566 9260 8735
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 6662 9168 7278
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9140 6322 9168 6598
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 5710 9168 6258
rect 9232 6186 9260 8502
rect 9324 7954 9352 10066
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9324 6390 9352 7890
rect 9416 7478 9444 10095
rect 9508 9382 9536 10542
rect 9586 10160 9642 10169
rect 9586 10095 9642 10104
rect 9600 9926 9628 10095
rect 9692 10062 9720 11562
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10336 11150 10364 11494
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 9846 10908 10154 10917
rect 9846 10906 9852 10908
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 10148 10906 10154 10908
rect 9908 10854 9910 10906
rect 10090 10854 10092 10906
rect 9846 10852 9852 10854
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 10148 10852 10154 10854
rect 9846 10843 10154 10852
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9876 10266 9904 10610
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9968 10130 9996 10610
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9586 9752 9642 9761
rect 9586 9687 9642 9696
rect 9496 9376 9548 9382
rect 9600 9353 9628 9687
rect 9496 9318 9548 9324
rect 9586 9344 9642 9353
rect 9508 9042 9536 9318
rect 9586 9279 9642 9288
rect 9692 9178 9720 9998
rect 9846 9820 10154 9829
rect 9846 9818 9852 9820
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 10148 9818 10154 9820
rect 9908 9766 9910 9818
rect 10090 9766 10092 9818
rect 9846 9764 9852 9766
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 10148 9764 10154 9766
rect 9846 9755 10154 9764
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9784 9353 9812 9454
rect 9770 9344 9826 9353
rect 9770 9279 9826 9288
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9600 8673 9628 8774
rect 9586 8664 9642 8673
rect 9586 8599 9642 8608
rect 9494 8528 9550 8537
rect 9494 8463 9550 8472
rect 9508 7886 9536 8463
rect 9784 8294 9812 9279
rect 9876 8974 9904 9658
rect 10336 9654 10364 10542
rect 10428 10198 10456 11494
rect 10520 11121 10548 12038
rect 10506 11112 10562 11121
rect 10506 11047 10562 11056
rect 10612 10810 10640 13892
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10704 11665 10732 11698
rect 10796 11694 10824 12242
rect 10784 11688 10836 11694
rect 10690 11656 10746 11665
rect 10784 11630 10836 11636
rect 10690 11591 10746 11600
rect 10796 11218 10824 11630
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10506 10024 10562 10033
rect 10506 9959 10562 9968
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9968 9178 9996 9522
rect 10230 9480 10286 9489
rect 10230 9415 10286 9424
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9968 8838 9996 9114
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9846 8732 10154 8741
rect 9846 8730 9852 8732
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 10148 8730 10154 8732
rect 9908 8678 9910 8730
rect 10090 8678 10092 8730
rect 9846 8676 9852 8678
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 10148 8676 10154 8678
rect 9846 8667 10154 8676
rect 9692 8266 9812 8294
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9220 6180 9272 6186
rect 9220 6122 9272 6128
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9324 4690 9352 6326
rect 9416 5098 9444 7414
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9508 6440 9536 7142
rect 9588 6452 9640 6458
rect 9508 6412 9588 6440
rect 9588 6394 9640 6400
rect 9692 5642 9720 8266
rect 10244 7886 10272 9415
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9784 7002 9812 7754
rect 9846 7644 10154 7653
rect 9846 7642 9852 7644
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 10148 7642 10154 7644
rect 9908 7590 9910 7642
rect 10090 7590 10092 7642
rect 9846 7588 9852 7590
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 10148 7588 10154 7590
rect 9846 7579 10154 7588
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9846 6556 10154 6565
rect 9846 6554 9852 6556
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 10148 6554 10154 6556
rect 9908 6502 9910 6554
rect 10090 6502 10092 6554
rect 9846 6500 9852 6502
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 10148 6500 10154 6502
rect 9846 6491 10154 6500
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 10244 5574 10272 6122
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 9846 5468 10154 5477
rect 9846 5466 9852 5468
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 10148 5466 10154 5468
rect 9908 5414 9910 5466
rect 10090 5414 10092 5466
rect 9846 5412 9852 5414
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 10148 5412 10154 5414
rect 9678 5400 9734 5409
rect 9846 5403 10154 5412
rect 9678 5335 9734 5344
rect 9692 5302 9720 5335
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9968 4826 9996 5170
rect 9956 4820 10008 4826
rect 9784 4780 9956 4808
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9324 4049 9352 4218
rect 9310 4040 9366 4049
rect 9310 3975 9366 3984
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9232 2378 9260 3130
rect 9416 2650 9444 4558
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 9508 800 9536 4490
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9600 3233 9628 4150
rect 9692 3398 9720 4694
rect 9784 4622 9812 4780
rect 9956 4762 10008 4768
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9784 4146 9812 4558
rect 9846 4380 10154 4389
rect 9846 4378 9852 4380
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 10148 4378 10154 4380
rect 9908 4326 9910 4378
rect 10090 4326 10092 4378
rect 9846 4324 9852 4326
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 10148 4324 10154 4326
rect 9846 4315 10154 4324
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9968 3466 9996 4082
rect 10244 4026 10272 4762
rect 10152 3998 10272 4026
rect 10152 3466 10180 3998
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9586 3224 9642 3233
rect 9586 3159 9642 3168
rect 9600 3126 9628 3159
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9692 2514 9720 3334
rect 9846 3292 10154 3301
rect 9846 3290 9852 3292
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 10148 3290 10154 3292
rect 9908 3238 9910 3290
rect 10090 3238 10092 3290
rect 9846 3236 9852 3238
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 10148 3236 10154 3238
rect 9846 3227 10154 3236
rect 10244 2774 10272 3878
rect 10336 3194 10364 9590
rect 10414 9208 10470 9217
rect 10414 9143 10470 9152
rect 10428 8838 10456 9143
rect 10416 8832 10468 8838
rect 10414 8800 10416 8809
rect 10468 8800 10470 8809
rect 10414 8735 10470 8744
rect 10520 8634 10548 9959
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10520 7750 10548 8570
rect 10704 8537 10732 8774
rect 10690 8528 10746 8537
rect 10690 8463 10746 8472
rect 10796 7818 10824 11154
rect 10784 7812 10836 7818
rect 10784 7754 10836 7760
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10414 6216 10470 6225
rect 10414 6151 10470 6160
rect 10428 4826 10456 6151
rect 10704 5710 10732 6326
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10416 4548 10468 4554
rect 10416 4490 10468 4496
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10428 3074 10456 4490
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10520 3126 10548 3334
rect 10336 3046 10456 3074
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10796 3058 10824 3878
rect 10888 3466 10916 13874
rect 10968 13456 11020 13462
rect 10968 13398 11020 13404
rect 10980 12209 11008 13398
rect 10966 12200 11022 12209
rect 10966 12135 11022 12144
rect 10980 10266 11008 12135
rect 11152 11552 11204 11558
rect 11150 11520 11152 11529
rect 11204 11520 11206 11529
rect 11150 11455 11206 11464
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11072 10810 11100 11018
rect 11256 10810 11284 15234
rect 11992 14006 12020 16510
rect 12162 16400 12218 16510
rect 14370 16400 14426 17200
rect 16578 16538 16634 17200
rect 17958 16552 18014 16561
rect 16578 16510 16896 16538
rect 16578 16400 16634 16510
rect 13544 15224 13596 15230
rect 13544 15166 13596 15172
rect 12070 14716 12378 14725
rect 12070 14714 12076 14716
rect 12132 14714 12156 14716
rect 12212 14714 12236 14716
rect 12292 14714 12316 14716
rect 12372 14714 12378 14716
rect 12132 14662 12134 14714
rect 12314 14662 12316 14714
rect 12070 14660 12076 14662
rect 12132 14660 12156 14662
rect 12212 14660 12236 14662
rect 12292 14660 12316 14662
rect 12372 14660 12378 14662
rect 12070 14651 12378 14660
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12070 13628 12378 13637
rect 12070 13626 12076 13628
rect 12132 13626 12156 13628
rect 12212 13626 12236 13628
rect 12292 13626 12316 13628
rect 12372 13626 12378 13628
rect 12132 13574 12134 13626
rect 12314 13574 12316 13626
rect 12070 13572 12076 13574
rect 12132 13572 12156 13574
rect 12212 13572 12236 13574
rect 12292 13572 12316 13574
rect 12372 13572 12378 13574
rect 12070 13563 12378 13572
rect 12452 13326 12480 13806
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12070 12540 12378 12549
rect 12070 12538 12076 12540
rect 12132 12538 12156 12540
rect 12212 12538 12236 12540
rect 12292 12538 12316 12540
rect 12372 12538 12378 12540
rect 12132 12486 12134 12538
rect 12314 12486 12316 12538
rect 12070 12484 12076 12486
rect 12132 12484 12156 12486
rect 12212 12484 12236 12486
rect 12292 12484 12316 12486
rect 12372 12484 12378 12486
rect 12070 12475 12378 12484
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11808 12238 11836 12378
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11992 11898 12020 12038
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11348 11150 11376 11494
rect 11440 11218 11468 11562
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11440 10996 11468 11154
rect 11348 10968 11468 10996
rect 11060 10804 11112 10810
rect 11244 10804 11296 10810
rect 11112 10764 11192 10792
rect 11060 10746 11112 10752
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 10266 11100 10474
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11164 10010 11192 10764
rect 11244 10746 11296 10752
rect 11164 9994 11284 10010
rect 11164 9988 11296 9994
rect 11164 9982 11244 9988
rect 11244 9930 11296 9936
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11072 8974 11100 9862
rect 11164 9042 11192 9862
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11348 8498 11376 10968
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11532 10130 11560 10406
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11624 10010 11652 11698
rect 12084 11694 12112 12242
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11898 12388 12038
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 11808 11529 11836 11630
rect 11794 11520 11850 11529
rect 11794 11455 11850 11464
rect 12070 11452 12378 11461
rect 12070 11450 12076 11452
rect 12132 11450 12156 11452
rect 12212 11450 12236 11452
rect 12292 11450 12316 11452
rect 12372 11450 12378 11452
rect 12132 11398 12134 11450
rect 12314 11398 12316 11450
rect 12070 11396 12076 11398
rect 12132 11396 12156 11398
rect 12212 11396 12236 11398
rect 12292 11396 12316 11398
rect 12372 11396 12378 11398
rect 12070 11387 12378 11396
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11532 9982 11652 10010
rect 11532 9110 11560 9982
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11624 9722 11652 9862
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 7886 11008 8230
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10980 7410 11008 7822
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10980 7206 11008 7346
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 6730 11008 7142
rect 11072 6798 11100 8434
rect 11440 7886 11468 8978
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 11256 7324 11284 7754
rect 11336 7336 11388 7342
rect 11256 7296 11336 7324
rect 11336 7278 11388 7284
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10980 6458 11008 6666
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10980 5642 11008 6394
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10980 5302 11008 5578
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 11242 4720 11298 4729
rect 11242 4655 11298 4664
rect 11256 4010 11284 4655
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11152 3732 11204 3738
rect 11072 3692 11152 3720
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 11072 3058 11100 3692
rect 11348 3720 11376 7278
rect 11440 7002 11468 7822
rect 11612 7472 11664 7478
rect 11610 7440 11612 7449
rect 11664 7440 11666 7449
rect 11610 7375 11666 7384
rect 11624 7324 11652 7375
rect 11532 7296 11652 7324
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11532 4049 11560 7296
rect 11716 6730 11744 10066
rect 11808 8634 11836 10134
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11624 4486 11652 5170
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11624 4282 11652 4422
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11518 4040 11574 4049
rect 11518 3975 11574 3984
rect 11428 3732 11480 3738
rect 11348 3692 11428 3720
rect 11152 3674 11204 3680
rect 11428 3674 11480 3680
rect 11624 3534 11652 4218
rect 11716 3534 11744 6054
rect 11808 5302 11836 8570
rect 11900 5574 11928 9318
rect 11992 8956 12020 11018
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12636 10470 12664 10678
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12070 10364 12378 10373
rect 12070 10362 12076 10364
rect 12132 10362 12156 10364
rect 12212 10362 12236 10364
rect 12292 10362 12316 10364
rect 12372 10362 12378 10364
rect 12132 10310 12134 10362
rect 12314 10310 12316 10362
rect 12070 10308 12076 10310
rect 12132 10308 12156 10310
rect 12212 10308 12236 10310
rect 12292 10308 12316 10310
rect 12372 10308 12378 10310
rect 12070 10299 12378 10308
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12360 9722 12388 9998
rect 12636 9994 12664 10406
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9722 12572 9862
rect 12728 9738 12756 11018
rect 12820 10810 12848 13874
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13004 12238 13032 12582
rect 13372 12306 13400 12786
rect 13556 12434 13584 15166
rect 14384 14482 14412 16400
rect 15014 15736 15070 15745
rect 15014 15671 15070 15680
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14294 14172 14602 14181
rect 14294 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14516 14170 14540 14172
rect 14596 14170 14602 14172
rect 14356 14118 14358 14170
rect 14538 14118 14540 14170
rect 14294 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14516 14116 14540 14118
rect 14596 14116 14602 14118
rect 14294 14107 14602 14116
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 13728 13864 13780 13870
rect 13726 13832 13728 13841
rect 13780 13832 13782 13841
rect 13726 13767 13782 13776
rect 14292 13530 14320 13942
rect 14752 13870 14780 14214
rect 14922 14104 14978 14113
rect 14922 14039 14978 14048
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13924 12850 13952 13194
rect 14294 13084 14602 13093
rect 14294 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14516 13082 14540 13084
rect 14596 13082 14602 13084
rect 14356 13030 14358 13082
rect 14538 13030 14540 13082
rect 14294 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14516 13028 14540 13030
rect 14596 13028 14602 13030
rect 14294 13019 14602 13028
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 13464 12406 13584 12434
rect 13084 12300 13136 12306
rect 13360 12300 13412 12306
rect 13136 12260 13216 12288
rect 13084 12242 13136 12248
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13096 11150 13124 11494
rect 13188 11150 13216 12260
rect 13360 12242 13412 12248
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13280 11558 13308 11630
rect 13464 11558 13492 12406
rect 14476 12102 14504 12786
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14844 12306 14872 12718
rect 14936 12374 14964 14039
rect 15028 12986 15056 15671
rect 15198 15464 15254 15473
rect 15198 15399 15254 15408
rect 15212 15366 15240 15399
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15290 15328 15346 15337
rect 15290 15263 15346 15272
rect 15304 15230 15332 15263
rect 15292 15224 15344 15230
rect 15292 15166 15344 15172
rect 15290 14920 15346 14929
rect 15290 14855 15346 14864
rect 15304 14550 15332 14855
rect 16518 14716 16826 14725
rect 16518 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16740 14714 16764 14716
rect 16820 14714 16826 14716
rect 16580 14662 16582 14714
rect 16762 14662 16764 14714
rect 16518 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16740 14660 16764 14662
rect 16820 14660 16826 14662
rect 16518 14651 16826 14660
rect 15292 14544 15344 14550
rect 15198 14512 15254 14521
rect 15108 14476 15160 14482
rect 15292 14486 15344 14492
rect 15198 14447 15254 14456
rect 15108 14418 15160 14424
rect 15120 14090 15148 14418
rect 15212 14414 15240 14447
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15304 14226 15332 14486
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 15304 14198 15424 14226
rect 15120 14062 15332 14090
rect 15120 13326 15148 14062
rect 15304 14006 15332 14062
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15212 13190 15240 13942
rect 15290 13288 15346 13297
rect 15290 13223 15346 13232
rect 15200 13184 15252 13190
rect 15198 13152 15200 13161
rect 15252 13152 15254 13161
rect 15198 13087 15254 13096
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 14924 12368 14976 12374
rect 14922 12336 14924 12345
rect 15016 12368 15068 12374
rect 14976 12336 14978 12345
rect 14832 12300 14884 12306
rect 15016 12310 15068 12316
rect 15106 12336 15162 12345
rect 14922 12271 14978 12280
rect 14832 12242 14884 12248
rect 14936 12245 14964 12271
rect 14844 12186 14872 12242
rect 14844 12158 14964 12186
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13004 10130 13032 10542
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9761 12940 9862
rect 12898 9752 12954 9761
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12532 9716 12584 9722
rect 12728 9710 12848 9738
rect 12532 9658 12584 9664
rect 12176 9602 12204 9658
rect 12176 9574 12480 9602
rect 12072 9512 12124 9518
rect 12070 9480 12072 9489
rect 12124 9480 12126 9489
rect 12070 9415 12126 9424
rect 12070 9276 12378 9285
rect 12070 9274 12076 9276
rect 12132 9274 12156 9276
rect 12212 9274 12236 9276
rect 12292 9274 12316 9276
rect 12372 9274 12378 9276
rect 12132 9222 12134 9274
rect 12314 9222 12316 9274
rect 12070 9220 12076 9222
rect 12132 9220 12156 9222
rect 12212 9220 12236 9222
rect 12292 9220 12316 9222
rect 12372 9220 12378 9222
rect 12070 9211 12378 9220
rect 12452 9110 12480 9574
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12440 9104 12492 9110
rect 12438 9072 12440 9081
rect 12492 9072 12494 9081
rect 12438 9007 12494 9016
rect 12072 8968 12124 8974
rect 11992 8928 12072 8956
rect 12072 8910 12124 8916
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 11992 6882 12020 8774
rect 12070 8188 12378 8197
rect 12070 8186 12076 8188
rect 12132 8186 12156 8188
rect 12212 8186 12236 8188
rect 12292 8186 12316 8188
rect 12372 8186 12378 8188
rect 12132 8134 12134 8186
rect 12314 8134 12316 8186
rect 12070 8132 12076 8134
rect 12132 8132 12156 8134
rect 12212 8132 12236 8134
rect 12292 8132 12316 8134
rect 12372 8132 12378 8134
rect 12070 8123 12378 8132
rect 12070 7100 12378 7109
rect 12070 7098 12076 7100
rect 12132 7098 12156 7100
rect 12212 7098 12236 7100
rect 12292 7098 12316 7100
rect 12372 7098 12378 7100
rect 12132 7046 12134 7098
rect 12314 7046 12316 7098
rect 12070 7044 12076 7046
rect 12132 7044 12156 7046
rect 12212 7044 12236 7046
rect 12292 7044 12316 7046
rect 12372 7044 12378 7046
rect 12070 7035 12378 7044
rect 11992 6854 12112 6882
rect 12084 6798 12112 6854
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 11992 5896 12020 6666
rect 12452 6118 12480 8774
rect 12636 7290 12664 9386
rect 12728 9042 12756 9522
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12820 8974 12848 9710
rect 12898 9687 12954 9696
rect 13004 9636 13032 10066
rect 12912 9608 13032 9636
rect 12912 9518 12940 9608
rect 13280 9586 13308 11494
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13464 10810 13492 10950
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13556 10062 13584 12038
rect 14294 11996 14602 12005
rect 14294 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14516 11994 14540 11996
rect 14596 11994 14602 11996
rect 14356 11942 14358 11994
rect 14538 11942 14540 11994
rect 14294 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14516 11940 14540 11942
rect 14596 11940 14602 11942
rect 14294 11931 14602 11940
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13648 11218 13676 11630
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12912 9382 12940 9454
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 13004 8838 13032 9454
rect 13280 8838 13308 9522
rect 13452 9172 13504 9178
rect 13372 9110 13400 9141
rect 13452 9114 13504 9120
rect 13360 9104 13412 9110
rect 13358 9072 13360 9081
rect 13412 9072 13414 9081
rect 13358 9007 13414 9016
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 12898 7848 12954 7857
rect 12898 7783 12954 7792
rect 12912 7546 12940 7783
rect 13280 7721 13308 8774
rect 13266 7712 13322 7721
rect 13266 7647 13322 7656
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12636 7262 12940 7290
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12070 6012 12378 6021
rect 12070 6010 12076 6012
rect 12132 6010 12156 6012
rect 12212 6010 12236 6012
rect 12292 6010 12316 6012
rect 12372 6010 12378 6012
rect 12132 5958 12134 6010
rect 12314 5958 12316 6010
rect 12070 5956 12076 5958
rect 12132 5956 12156 5958
rect 12212 5956 12236 5958
rect 12292 5956 12316 5958
rect 12372 5956 12378 5958
rect 12070 5947 12378 5956
rect 12072 5908 12124 5914
rect 11992 5868 12072 5896
rect 12072 5850 12124 5856
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12084 5574 12112 5646
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 12070 4924 12378 4933
rect 12070 4922 12076 4924
rect 12132 4922 12156 4924
rect 12212 4922 12236 4924
rect 12292 4922 12316 4924
rect 12372 4922 12378 4924
rect 12132 4870 12134 4922
rect 12314 4870 12316 4922
rect 12070 4868 12076 4870
rect 12132 4868 12156 4870
rect 12212 4868 12236 4870
rect 12292 4868 12316 4870
rect 12372 4868 12378 4870
rect 12070 4859 12378 4868
rect 12070 3836 12378 3845
rect 12070 3834 12076 3836
rect 12132 3834 12156 3836
rect 12212 3834 12236 3836
rect 12292 3834 12316 3836
rect 12372 3834 12378 3836
rect 12132 3782 12134 3834
rect 12314 3782 12316 3834
rect 12070 3780 12076 3782
rect 12132 3780 12156 3782
rect 12212 3780 12236 3782
rect 12292 3780 12316 3782
rect 12372 3780 12378 3782
rect 12070 3771 12378 3780
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11624 3126 11652 3470
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 10784 3052 10836 3058
rect 10336 2854 10364 3046
rect 10784 2994 10836 3000
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10152 2746 10272 2774
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9678 2408 9734 2417
rect 10152 2394 10180 2746
rect 10152 2366 10364 2394
rect 9678 2343 9680 2352
rect 9732 2343 9734 2352
rect 9680 2314 9732 2320
rect 9846 2204 10154 2213
rect 9846 2202 9852 2204
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 10148 2202 10154 2204
rect 9908 2150 9910 2202
rect 10090 2150 10092 2202
rect 9846 2148 9852 2150
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 10148 2148 10154 2150
rect 9846 2139 10154 2148
rect 10336 800 10364 2366
rect 11072 2310 11100 2994
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11164 800 11192 2790
rect 11624 2650 11652 3062
rect 12070 2748 12378 2757
rect 12070 2746 12076 2748
rect 12132 2746 12156 2748
rect 12212 2746 12236 2748
rect 12292 2746 12316 2748
rect 12372 2746 12378 2748
rect 12132 2694 12134 2746
rect 12314 2694 12316 2746
rect 12070 2692 12076 2694
rect 12132 2692 12156 2694
rect 12212 2692 12236 2694
rect 12292 2692 12316 2694
rect 12372 2692 12378 2694
rect 12070 2683 12378 2692
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 12346 2544 12402 2553
rect 12346 2479 12402 2488
rect 12360 2446 12388 2479
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 11980 2372 12032 2378
rect 11980 2314 12032 2320
rect 11992 800 12020 2314
rect 12452 2038 12480 6054
rect 12820 4146 12848 7142
rect 12912 6866 12940 7262
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 13280 6769 13308 7647
rect 13372 7546 13400 9007
rect 13464 8514 13492 9114
rect 13556 8809 13584 9658
rect 13648 9382 13676 11018
rect 13740 10810 13768 11698
rect 14752 11558 14780 11698
rect 14830 11656 14886 11665
rect 14830 11591 14886 11600
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14462 11384 14518 11393
rect 14752 11354 14780 11494
rect 14844 11354 14872 11591
rect 14462 11319 14518 11328
rect 14740 11348 14792 11354
rect 14200 11286 14228 11317
rect 14188 11280 14240 11286
rect 14186 11248 14188 11257
rect 14240 11248 14242 11257
rect 14186 11183 14242 11192
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13832 10742 13860 11086
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13542 8800 13598 8809
rect 13542 8735 13598 8744
rect 13464 8486 13584 8514
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13464 7886 13492 8366
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13464 7546 13492 7822
rect 13556 7750 13584 8486
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13266 6760 13322 6769
rect 13266 6695 13322 6704
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 13004 6322 13032 6598
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12912 6118 12940 6258
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 12912 4622 12940 6054
rect 13188 5234 13216 6054
rect 13372 5896 13400 7482
rect 13464 7002 13492 7482
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13464 6458 13492 6938
rect 13556 6934 13584 7686
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13556 6390 13584 6870
rect 13648 6798 13676 9318
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13740 6662 13768 10542
rect 13832 7546 13860 10542
rect 13924 10130 13952 10950
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13924 8566 13952 10066
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 13924 8022 13952 8502
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13832 6186 13860 7346
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13452 5908 13504 5914
rect 13372 5868 13452 5896
rect 13452 5850 13504 5856
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 4826 13032 4966
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12544 2446 12572 3946
rect 13096 3058 13124 5034
rect 13464 4826 13492 5646
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13832 5302 13860 5578
rect 13924 5370 13952 7686
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13464 4282 13492 4762
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13464 3738 13492 4218
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13464 3126 13492 3674
rect 13556 3534 13584 4694
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 12900 2848 12952 2854
rect 12820 2796 12900 2802
rect 12820 2790 12952 2796
rect 12820 2774 12940 2790
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12440 2032 12492 2038
rect 12440 1974 12492 1980
rect 12820 800 12848 2774
rect 14016 2446 14044 10406
rect 14200 9518 14228 11183
rect 14476 11150 14504 11319
rect 14740 11290 14792 11296
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14738 11248 14794 11257
rect 14738 11183 14794 11192
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14294 10908 14602 10917
rect 14294 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14516 10906 14540 10908
rect 14596 10906 14602 10908
rect 14356 10854 14358 10906
rect 14538 10854 14540 10906
rect 14294 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14516 10852 14540 10854
rect 14596 10852 14602 10854
rect 14294 10843 14602 10852
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14476 10062 14504 10406
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14294 9820 14602 9829
rect 14294 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14516 9818 14540 9820
rect 14596 9818 14602 9820
rect 14356 9766 14358 9818
rect 14538 9766 14540 9818
rect 14294 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14516 9764 14540 9766
rect 14596 9764 14602 9766
rect 14294 9755 14602 9764
rect 14648 9716 14700 9722
rect 14752 9704 14780 11183
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14844 9722 14872 10610
rect 14936 10606 14964 12158
rect 15028 12102 15056 12310
rect 15106 12271 15162 12280
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15120 11898 15148 12271
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 15028 11540 15056 11766
rect 15108 11688 15160 11694
rect 15160 11648 15240 11676
rect 15108 11630 15160 11636
rect 15028 11512 15148 11540
rect 15120 11354 15148 11512
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15028 10742 15056 11290
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 10810 15148 10950
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14936 10130 14964 10542
rect 15108 10464 15160 10470
rect 15212 10452 15240 11648
rect 15304 10538 15332 13223
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15160 10424 15240 10452
rect 15108 10406 15160 10412
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14700 9676 14780 9704
rect 14648 9658 14700 9664
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14108 9042 14136 9454
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14108 8498 14136 8978
rect 14200 8838 14228 9454
rect 14384 9110 14412 9590
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14108 8090 14136 8434
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14200 7970 14228 8774
rect 14294 8732 14602 8741
rect 14294 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14516 8730 14540 8732
rect 14596 8730 14602 8732
rect 14356 8678 14358 8730
rect 14538 8678 14540 8730
rect 14294 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14516 8676 14540 8678
rect 14596 8676 14602 8678
rect 14294 8667 14602 8676
rect 14660 8634 14688 9318
rect 14752 9178 14780 9676
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14844 9178 14872 9454
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14832 8832 14884 8838
rect 14830 8800 14832 8809
rect 14884 8800 14886 8809
rect 14830 8735 14886 8744
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14936 8401 14964 10066
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 15028 9450 15056 9862
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 14922 8392 14978 8401
rect 14922 8327 14924 8336
rect 14976 8327 14978 8336
rect 14924 8298 14976 8304
rect 14108 7942 14228 7970
rect 14108 6322 14136 7942
rect 14294 7644 14602 7653
rect 14294 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14516 7642 14540 7644
rect 14596 7642 14602 7644
rect 14356 7590 14358 7642
rect 14538 7590 14540 7642
rect 14294 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14516 7588 14540 7590
rect 14596 7588 14602 7590
rect 14294 7579 14602 7588
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 14108 2922 14136 4490
rect 14200 4146 14228 7482
rect 14294 6556 14602 6565
rect 14294 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14516 6554 14540 6556
rect 14596 6554 14602 6556
rect 14356 6502 14358 6554
rect 14538 6502 14540 6554
rect 14294 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14516 6500 14540 6502
rect 14596 6500 14602 6502
rect 14294 6491 14602 6500
rect 15120 6458 15148 10406
rect 15396 10112 15424 14198
rect 16684 13938 16712 14350
rect 16868 14074 16896 16510
rect 17958 16487 18014 16496
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16304 13864 16356 13870
rect 16302 13832 16304 13841
rect 16356 13832 16358 13841
rect 16302 13767 16358 13776
rect 16518 13628 16826 13637
rect 16518 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16740 13626 16764 13628
rect 16820 13626 16826 13628
rect 16580 13574 16582 13626
rect 16762 13574 16764 13626
rect 16518 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16740 13572 16764 13574
rect 16820 13572 16826 13574
rect 16518 13563 16826 13572
rect 17866 13152 17922 13161
rect 17866 13087 17922 13096
rect 17880 12986 17908 13087
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 16026 12880 16082 12889
rect 16026 12815 16082 12824
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 11014 15516 11494
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15580 10130 15608 11154
rect 15672 10674 15700 11630
rect 15936 11552 15988 11558
rect 15856 11500 15936 11506
rect 15856 11494 15988 11500
rect 15856 11478 15976 11494
rect 15856 11218 15884 11478
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15568 10124 15620 10130
rect 15396 10084 15516 10112
rect 15290 10024 15346 10033
rect 15290 9959 15346 9968
rect 15304 9654 15332 9959
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15396 8838 15424 9862
rect 15488 9654 15516 10084
rect 15568 10066 15620 10072
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15304 7546 15332 8230
rect 15488 7993 15516 9386
rect 15580 8974 15608 10066
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15764 9722 15792 9862
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15580 8566 15608 8910
rect 15672 8566 15700 9454
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15474 7984 15530 7993
rect 15474 7919 15530 7928
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15488 7546 15516 7822
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15580 6662 15608 8502
rect 15672 7449 15700 8502
rect 15764 8090 15792 8774
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15750 7984 15806 7993
rect 15750 7919 15806 7928
rect 15764 7478 15792 7919
rect 15752 7472 15804 7478
rect 15658 7440 15714 7449
rect 15752 7414 15804 7420
rect 15658 7375 15714 7384
rect 15764 7290 15792 7414
rect 15856 7342 15884 11154
rect 16040 11150 16068 12815
rect 16518 12540 16826 12549
rect 16518 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16740 12538 16764 12540
rect 16820 12538 16826 12540
rect 16580 12486 16582 12538
rect 16762 12486 16764 12538
rect 16518 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16740 12484 16764 12486
rect 16820 12484 16826 12486
rect 16518 12475 16826 12484
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17500 12232 17552 12238
rect 17052 12158 17356 12186
rect 17500 12174 17552 12180
rect 16948 12096 17000 12102
rect 17052 12084 17080 12158
rect 17328 12102 17356 12158
rect 17000 12056 17080 12084
rect 17132 12096 17184 12102
rect 16948 12038 17000 12044
rect 17132 12038 17184 12044
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 16854 11656 16910 11665
rect 16396 11620 16448 11626
rect 16854 11591 16910 11600
rect 16396 11562 16448 11568
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 15936 9648 15988 9654
rect 15936 9590 15988 9596
rect 15948 8673 15976 9590
rect 16040 9450 16068 11086
rect 16132 10674 16160 11086
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 15934 8664 15990 8673
rect 15934 8599 15990 8608
rect 15934 8256 15990 8265
rect 15934 8191 15990 8200
rect 15948 7993 15976 8191
rect 15934 7984 15990 7993
rect 15934 7919 15990 7928
rect 15672 7262 15792 7290
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15672 7041 15700 7262
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15658 7032 15714 7041
rect 15658 6967 15714 6976
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14844 5710 14872 6258
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14294 5468 14602 5477
rect 14294 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14516 5466 14540 5468
rect 14596 5466 14602 5468
rect 14356 5414 14358 5466
rect 14538 5414 14540 5466
rect 14294 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14516 5412 14540 5414
rect 14596 5412 14602 5414
rect 14294 5403 14602 5412
rect 14844 5302 14872 5646
rect 14832 5296 14884 5302
rect 14832 5238 14884 5244
rect 14294 4380 14602 4389
rect 14294 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14516 4378 14540 4380
rect 14596 4378 14602 4380
rect 14356 4326 14358 4378
rect 14538 4326 14540 4378
rect 14294 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14516 4324 14540 4326
rect 14596 4324 14602 4326
rect 14294 4315 14602 4324
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14294 3292 14602 3301
rect 14294 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14516 3290 14540 3292
rect 14596 3290 14602 3292
rect 14356 3238 14358 3290
rect 14538 3238 14540 3290
rect 14294 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14516 3236 14540 3238
rect 14596 3236 14602 3238
rect 14294 3227 14602 3236
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14476 3097 14504 3130
rect 14462 3088 14518 3097
rect 14462 3023 14518 3032
rect 14370 2952 14426 2961
rect 14096 2916 14148 2922
rect 14370 2887 14372 2896
rect 14096 2858 14148 2864
rect 14424 2887 14426 2896
rect 14372 2858 14424 2864
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 14936 2378 14964 6190
rect 15198 5672 15254 5681
rect 15108 5636 15160 5642
rect 15198 5607 15254 5616
rect 15108 5578 15160 5584
rect 15120 3942 15148 5578
rect 15212 4554 15240 5607
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15212 3738 15240 4490
rect 15290 4040 15346 4049
rect 15290 3975 15346 3984
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 14924 2372 14976 2378
rect 14924 2314 14976 2320
rect 13832 1442 13860 2314
rect 14294 2204 14602 2213
rect 14294 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14516 2202 14540 2204
rect 14596 2202 14602 2204
rect 14356 2150 14358 2202
rect 14538 2150 14540 2202
rect 14294 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14516 2148 14540 2150
rect 14596 2148 14602 2150
rect 14294 2139 14602 2148
rect 14464 1556 14516 1562
rect 14464 1498 14516 1504
rect 13648 1414 13860 1442
rect 13648 800 13676 1414
rect 14476 800 14504 1498
rect 15304 800 15332 3975
rect 15396 3108 15424 6598
rect 15568 6384 15620 6390
rect 15568 6326 15620 6332
rect 15580 5914 15608 6326
rect 15672 5914 15700 6967
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15580 5370 15608 5850
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15488 4078 15516 5170
rect 15580 4690 15608 5306
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15488 3738 15516 4014
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15580 3602 15608 4626
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15672 3466 15700 5510
rect 15764 4622 15792 7142
rect 15948 6458 15976 7919
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15948 6066 15976 6394
rect 16040 6322 16068 8842
rect 16132 8378 16160 10610
rect 16224 10606 16252 10950
rect 16212 10600 16264 10606
rect 16210 10568 16212 10577
rect 16304 10600 16356 10606
rect 16264 10568 16266 10577
rect 16304 10542 16356 10548
rect 16210 10503 16266 10512
rect 16224 10169 16252 10503
rect 16210 10160 16266 10169
rect 16210 10095 16266 10104
rect 16210 8936 16266 8945
rect 16210 8871 16266 8880
rect 16224 8838 16252 8871
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16316 8650 16344 10542
rect 16408 10033 16436 11562
rect 16518 11452 16826 11461
rect 16518 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16740 11450 16764 11452
rect 16820 11450 16826 11452
rect 16580 11398 16582 11450
rect 16762 11398 16764 11450
rect 16518 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16740 11396 16764 11398
rect 16820 11396 16826 11398
rect 16518 11387 16826 11396
rect 16764 11280 16816 11286
rect 16764 11222 16816 11228
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16592 10810 16620 11018
rect 16776 10810 16804 11222
rect 16868 11150 16896 11591
rect 16856 11144 16908 11150
rect 16960 11121 16988 12038
rect 17144 11898 17172 12038
rect 17512 11898 17540 12174
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17130 11792 17186 11801
rect 17040 11756 17092 11762
rect 17130 11727 17186 11736
rect 17040 11698 17092 11704
rect 17052 11354 17080 11698
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16856 11086 16908 11092
rect 16946 11112 17002 11121
rect 16946 11047 17002 11056
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16518 10364 16826 10373
rect 16518 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16740 10362 16764 10364
rect 16820 10362 16826 10364
rect 16580 10310 16582 10362
rect 16762 10310 16764 10362
rect 16518 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16740 10308 16764 10310
rect 16820 10308 16826 10310
rect 16518 10299 16826 10308
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16394 10024 16450 10033
rect 16394 9959 16450 9968
rect 16592 9654 16620 10066
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16684 9722 16712 9930
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16776 9518 16804 10066
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16408 8974 16436 9318
rect 16518 9276 16826 9285
rect 16518 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16740 9274 16764 9276
rect 16820 9274 16826 9276
rect 16580 9222 16582 9274
rect 16762 9222 16764 9274
rect 16518 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16740 9220 16764 9222
rect 16820 9220 16826 9222
rect 16518 9211 16826 9220
rect 16868 9058 16896 10950
rect 16776 9030 16896 9058
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16224 8622 16344 8650
rect 16592 8634 16620 8774
rect 16580 8628 16632 8634
rect 16224 8498 16252 8622
rect 16580 8570 16632 8576
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16316 8486 16528 8514
rect 16776 8498 16804 9030
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16316 8378 16344 8486
rect 16500 8430 16528 8486
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16132 8350 16344 8378
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16132 6662 16160 7346
rect 16212 7336 16264 7342
rect 16316 7313 16344 8350
rect 16408 7886 16436 8366
rect 16518 8188 16826 8197
rect 16518 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16740 8186 16764 8188
rect 16820 8186 16826 8188
rect 16580 8134 16582 8186
rect 16762 8134 16764 8186
rect 16518 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16740 8132 16764 8134
rect 16820 8132 16826 8134
rect 16518 8123 16826 8132
rect 16396 7880 16448 7886
rect 16868 7857 16896 8910
rect 16960 8634 16988 11047
rect 17144 11014 17172 11727
rect 17604 11218 17632 12242
rect 17880 12238 17908 12922
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17420 10810 17448 10950
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17604 10606 17632 11154
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17038 10432 17094 10441
rect 17038 10367 17094 10376
rect 17052 9654 17080 10367
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 17052 9353 17080 9454
rect 17038 9344 17094 9353
rect 17038 9279 17094 9288
rect 17144 9178 17172 10542
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17316 9512 17368 9518
rect 17222 9480 17278 9489
rect 17316 9454 17368 9460
rect 17222 9415 17278 9424
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17052 8974 17080 9114
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16960 8362 16988 8570
rect 17052 8498 17080 8774
rect 17144 8673 17172 8842
rect 17130 8664 17186 8673
rect 17130 8599 17186 8608
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 17038 8392 17094 8401
rect 16948 8356 17000 8362
rect 17038 8327 17094 8336
rect 16948 8298 17000 8304
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 16396 7822 16448 7828
rect 16854 7848 16910 7857
rect 16212 7278 16264 7284
rect 16302 7304 16358 7313
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15856 6038 15976 6066
rect 15856 5914 15884 6038
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 16040 5098 16068 6258
rect 16224 5681 16252 7278
rect 16302 7239 16358 7248
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16316 5778 16344 7142
rect 16408 6798 16436 7822
rect 16854 7783 16910 7792
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16518 7100 16826 7109
rect 16518 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16740 7098 16764 7100
rect 16820 7098 16826 7100
rect 16580 7046 16582 7098
rect 16762 7046 16764 7098
rect 16518 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16740 7044 16764 7046
rect 16820 7044 16826 7046
rect 16518 7035 16826 7044
rect 16868 6914 16896 7346
rect 16776 6886 16896 6914
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16486 6760 16542 6769
rect 16408 6322 16436 6734
rect 16486 6695 16542 6704
rect 16580 6724 16632 6730
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16500 6202 16528 6695
rect 16580 6666 16632 6672
rect 16408 6174 16528 6202
rect 16592 6186 16620 6666
rect 16776 6254 16804 6886
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16580 6180 16632 6186
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 16210 5672 16266 5681
rect 16210 5607 16266 5616
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15660 3460 15712 3466
rect 15660 3402 15712 3408
rect 15568 3120 15620 3126
rect 15396 3080 15568 3108
rect 15568 3062 15620 3068
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15488 2446 15516 2790
rect 15764 2446 15792 3878
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15856 3058 15884 3470
rect 15948 3058 15976 4422
rect 16132 4214 16160 5510
rect 16224 4486 16252 5510
rect 16408 5370 16436 6174
rect 16580 6122 16632 6128
rect 16518 6012 16826 6021
rect 16518 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16740 6010 16764 6012
rect 16820 6010 16826 6012
rect 16580 5958 16582 6010
rect 16762 5958 16764 6010
rect 16518 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16740 5956 16764 5958
rect 16820 5956 16826 5958
rect 16518 5947 16826 5956
rect 16868 5896 16896 6666
rect 16684 5868 16896 5896
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16120 4208 16172 4214
rect 16120 4150 16172 4156
rect 16316 4146 16344 5170
rect 16684 5098 16712 5868
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 16776 5166 16804 5578
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16672 5092 16724 5098
rect 16672 5034 16724 5040
rect 16518 4924 16826 4933
rect 16518 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16740 4922 16764 4924
rect 16820 4922 16826 4924
rect 16580 4870 16582 4922
rect 16762 4870 16764 4922
rect 16518 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16740 4868 16764 4870
rect 16820 4868 16826 4870
rect 16518 4859 16826 4868
rect 16868 4690 16896 5714
rect 16960 5302 16988 7958
rect 17052 7818 17080 8327
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17144 8022 17172 8230
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 17236 7886 17264 9415
rect 17328 7954 17356 9454
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17040 7812 17092 7818
rect 17040 7754 17092 7760
rect 17132 7812 17184 7818
rect 17132 7754 17184 7760
rect 17040 6928 17092 6934
rect 17040 6870 17092 6876
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16684 4554 16712 4626
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16396 4480 16448 4486
rect 16396 4422 16448 4428
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16408 4282 16436 4422
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16118 3904 16174 3913
rect 16118 3839 16174 3848
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 15856 2650 15884 2994
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 16040 1562 16068 2926
rect 16028 1556 16080 1562
rect 16028 1498 16080 1504
rect 16132 800 16160 3839
rect 4066 776 4122 785
rect 4066 711 4122 720
rect 4526 0 4582 800
rect 5354 0 5410 800
rect 6182 0 6238 800
rect 7010 0 7066 800
rect 7838 0 7894 800
rect 8666 0 8722 800
rect 9494 0 9550 800
rect 10322 0 10378 800
rect 11150 0 11206 800
rect 11978 0 12034 800
rect 12806 0 12862 800
rect 13634 0 13690 800
rect 14462 0 14518 800
rect 15290 0 15346 800
rect 16118 0 16174 800
rect 16316 649 16344 3946
rect 16518 3836 16826 3845
rect 16518 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16740 3834 16764 3836
rect 16820 3834 16826 3836
rect 16580 3782 16582 3834
rect 16762 3782 16764 3834
rect 16518 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16740 3780 16764 3782
rect 16820 3780 16826 3782
rect 16518 3771 16826 3780
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16592 3058 16620 3334
rect 16868 3194 16896 4422
rect 16960 4282 16988 5102
rect 17052 4826 17080 6870
rect 17144 6118 17172 7754
rect 17236 6934 17264 7822
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17224 6792 17276 6798
rect 17222 6760 17224 6769
rect 17276 6760 17278 6769
rect 17328 6730 17356 7890
rect 17222 6695 17278 6704
rect 17316 6724 17368 6730
rect 17316 6666 17368 6672
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6458 17264 6598
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 16946 3632 17002 3641
rect 16946 3567 17002 3576
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 16518 2748 16826 2757
rect 16518 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16740 2746 16764 2748
rect 16820 2746 16826 2748
rect 16580 2694 16582 2746
rect 16762 2694 16764 2746
rect 16518 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16740 2692 16764 2694
rect 16820 2692 16826 2694
rect 16518 2683 16826 2692
rect 16868 2582 16896 2858
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 16684 2038 16712 2518
rect 16672 2032 16724 2038
rect 16672 1974 16724 1980
rect 16960 800 16988 3567
rect 17052 3466 17080 4626
rect 17144 4486 17172 6054
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17236 5098 17264 5850
rect 17328 5710 17356 6054
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17316 5568 17368 5574
rect 17316 5510 17368 5516
rect 17328 5370 17356 5510
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17420 5234 17448 9862
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17512 9110 17540 9318
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17512 8090 17540 8774
rect 17604 8566 17632 9590
rect 17696 9217 17724 12038
rect 17972 11898 18000 16487
rect 18786 16400 18842 17200
rect 18800 14006 18828 16400
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18892 12434 18920 13806
rect 18892 12406 19104 12434
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17788 11150 17816 11834
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17880 11098 17908 11494
rect 17972 11286 18000 11834
rect 17960 11280 18012 11286
rect 17960 11222 18012 11228
rect 17880 11070 18000 11098
rect 17866 10976 17922 10985
rect 17866 10911 17922 10920
rect 17880 10674 17908 10911
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17972 10554 18000 11070
rect 18156 10962 18184 12310
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18248 11150 18276 11766
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18696 11280 18748 11286
rect 18696 11222 18748 11228
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18156 10934 18276 10962
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 17880 10526 18000 10554
rect 17880 9722 17908 10526
rect 18156 10062 18184 10678
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17682 9208 17738 9217
rect 17682 9143 17738 9152
rect 17696 8974 17724 9143
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17684 8832 17736 8838
rect 17682 8800 17684 8809
rect 17736 8800 17738 8809
rect 17682 8735 17738 8744
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17590 8392 17646 8401
rect 17590 8327 17646 8336
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17604 7478 17632 8327
rect 17696 7818 17724 8735
rect 17788 8650 17816 9522
rect 17880 9081 17908 9658
rect 17866 9072 17922 9081
rect 17866 9007 17922 9016
rect 17880 8809 17908 9007
rect 17866 8800 17922 8809
rect 17866 8735 17922 8744
rect 17788 8622 17908 8650
rect 17776 8560 17828 8566
rect 17776 8502 17828 8508
rect 17684 7812 17736 7818
rect 17684 7754 17736 7760
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17592 7336 17644 7342
rect 17498 7304 17554 7313
rect 17592 7278 17644 7284
rect 17498 7239 17554 7248
rect 17512 6322 17540 7239
rect 17604 6866 17632 7278
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17512 5681 17540 5714
rect 17498 5672 17554 5681
rect 17604 5642 17632 6802
rect 17498 5607 17554 5616
rect 17592 5636 17644 5642
rect 17592 5578 17644 5584
rect 17500 5296 17552 5302
rect 17500 5238 17552 5244
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17224 5092 17276 5098
rect 17224 5034 17276 5040
rect 17328 4690 17356 5102
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 17144 3058 17172 4422
rect 17236 3738 17264 4490
rect 17328 4078 17356 4626
rect 17512 4146 17540 5238
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17604 4622 17632 4762
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17316 4072 17368 4078
rect 17408 4072 17460 4078
rect 17316 4014 17368 4020
rect 17406 4040 17408 4049
rect 17460 4040 17462 4049
rect 17406 3975 17462 3984
rect 17420 3890 17448 3975
rect 17328 3862 17448 3890
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17052 2854 17080 2994
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 2310 17080 2790
rect 17144 2650 17172 2994
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17144 2446 17172 2586
rect 17236 2582 17264 3470
rect 17328 2854 17356 3862
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17328 1465 17356 2246
rect 17314 1456 17370 1465
rect 17314 1391 17370 1400
rect 17420 1057 17448 3334
rect 17512 2922 17540 4082
rect 17604 3398 17632 4558
rect 17696 3534 17724 7754
rect 17788 4554 17816 8502
rect 17880 8362 17908 8622
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17866 7984 17922 7993
rect 17866 7919 17922 7928
rect 17880 7886 17908 7919
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17880 7546 17908 7822
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17880 6254 17908 7278
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17776 4548 17828 4554
rect 17776 4490 17828 4496
rect 17788 4282 17816 4490
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17696 1873 17724 2246
rect 17682 1864 17738 1873
rect 17682 1799 17738 1808
rect 17406 1048 17462 1057
rect 17406 983 17462 992
rect 17788 800 17816 4014
rect 17880 3602 17908 6190
rect 17972 5545 18000 9862
rect 18064 9722 18092 9998
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 18142 9616 18198 9625
rect 18142 9551 18198 9560
rect 18156 8498 18184 9551
rect 18248 8974 18276 10934
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18050 8392 18106 8401
rect 18050 8327 18052 8336
rect 18104 8327 18106 8336
rect 18052 8298 18104 8304
rect 18052 8016 18104 8022
rect 18050 7984 18052 7993
rect 18104 7984 18106 7993
rect 18050 7919 18106 7928
rect 18050 7168 18106 7177
rect 18050 7103 18106 7112
rect 18064 7002 18092 7103
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18050 6488 18106 6497
rect 18050 6423 18106 6432
rect 18064 6390 18092 6423
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17958 5536 18014 5545
rect 17958 5471 18014 5480
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17880 2990 17908 3538
rect 17972 3534 18000 4082
rect 18064 3738 18092 6326
rect 18156 6202 18184 8434
rect 18248 6322 18276 8910
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18340 7426 18368 8026
rect 18432 7585 18460 8774
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18418 7576 18474 7585
rect 18418 7511 18474 7520
rect 18340 7398 18460 7426
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18340 6458 18368 7278
rect 18432 6866 18460 7398
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18418 6760 18474 6769
rect 18418 6695 18474 6704
rect 18432 6662 18460 6695
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18156 6174 18368 6202
rect 18432 6186 18460 6394
rect 18524 6361 18552 8298
rect 18510 6352 18566 6361
rect 18510 6287 18566 6296
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18156 4826 18184 5510
rect 18248 5370 18276 5510
rect 18340 5370 18368 6174
rect 18420 6180 18472 6186
rect 18420 6122 18472 6128
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18142 4720 18198 4729
rect 18142 4655 18198 4664
rect 18156 4282 18184 4655
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17960 3528 18012 3534
rect 18248 3505 18276 4422
rect 17960 3470 18012 3476
rect 18234 3496 18290 3505
rect 18234 3431 18290 3440
rect 18340 3194 18368 5170
rect 18432 4826 18460 6122
rect 18616 5953 18644 9862
rect 18602 5944 18658 5953
rect 18602 5879 18658 5888
rect 18708 5137 18736 11222
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18694 5128 18750 5137
rect 18694 5063 18750 5072
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 18050 3088 18106 3097
rect 18050 3023 18106 3032
rect 17868 2984 17920 2990
rect 17866 2952 17868 2961
rect 17920 2952 17922 2961
rect 17866 2887 17922 2896
rect 18064 2650 18092 3023
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 18156 2446 18184 2790
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 17880 2106 17908 2382
rect 18420 2304 18472 2310
rect 18418 2272 18420 2281
rect 18472 2272 18474 2281
rect 18418 2207 18474 2216
rect 17868 2100 17920 2106
rect 17868 2042 17920 2048
rect 18524 2038 18552 4558
rect 18800 2689 18828 10474
rect 18892 4321 18920 11290
rect 18970 10568 19026 10577
rect 18970 10503 18972 10512
rect 19024 10503 19026 10512
rect 18972 10474 19024 10480
rect 18972 10192 19024 10198
rect 18972 10134 19024 10140
rect 18878 4312 18934 4321
rect 18878 4247 18934 4256
rect 18984 3913 19012 10134
rect 19076 4078 19104 12406
rect 19248 10532 19300 10538
rect 19248 10474 19300 10480
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19168 5030 19196 6734
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19260 4622 19288 10474
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19352 4146 19380 7346
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 18970 3904 19026 3913
rect 18970 3839 19026 3848
rect 18786 2680 18842 2689
rect 18786 2615 18842 2624
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 18512 2032 18564 2038
rect 18512 1974 18564 1980
rect 18616 800 18644 2450
rect 16302 640 16358 649
rect 16302 575 16358 584
rect 16946 0 17002 800
rect 17774 0 17830 800
rect 18602 0 18658 800
<< via2 >>
rect 4434 16632 4490 16688
rect 3422 15408 3478 15464
rect 2778 14592 2834 14648
rect 1214 11328 1270 11384
rect 1122 10104 1178 10160
rect 938 5208 994 5264
rect 1858 12960 1914 13016
rect 1766 10512 1822 10568
rect 1766 9968 1822 10024
rect 1674 8472 1730 8528
rect 1674 7792 1730 7848
rect 1490 7656 1546 7712
rect 1490 7268 1546 7304
rect 1490 7248 1492 7268
rect 1492 7248 1544 7268
rect 1544 7248 1546 7268
rect 1490 6840 1546 6896
rect 1582 6432 1638 6488
rect 1398 6160 1454 6216
rect 2226 12688 2282 12744
rect 2318 12280 2374 12336
rect 2778 12552 2834 12608
rect 2502 11600 2558 11656
rect 2318 9968 2374 10024
rect 1950 8508 1952 8528
rect 1952 8508 2004 8528
rect 2004 8508 2006 8528
rect 1950 8472 2006 8508
rect 3180 14714 3236 14716
rect 3260 14714 3316 14716
rect 3340 14714 3396 14716
rect 3420 14714 3476 14716
rect 3180 14662 3226 14714
rect 3226 14662 3236 14714
rect 3260 14662 3290 14714
rect 3290 14662 3302 14714
rect 3302 14662 3316 14714
rect 3340 14662 3354 14714
rect 3354 14662 3366 14714
rect 3366 14662 3396 14714
rect 3420 14662 3430 14714
rect 3430 14662 3476 14714
rect 3180 14660 3236 14662
rect 3260 14660 3316 14662
rect 3340 14660 3396 14662
rect 3420 14660 3476 14662
rect 3974 16224 4030 16280
rect 4066 15816 4122 15872
rect 3514 14184 3570 14240
rect 3422 13776 3478 13832
rect 3180 13626 3236 13628
rect 3260 13626 3316 13628
rect 3340 13626 3396 13628
rect 3420 13626 3476 13628
rect 3180 13574 3226 13626
rect 3226 13574 3236 13626
rect 3260 13574 3290 13626
rect 3290 13574 3302 13626
rect 3302 13574 3316 13626
rect 3340 13574 3354 13626
rect 3354 13574 3366 13626
rect 3366 13574 3396 13626
rect 3420 13574 3430 13626
rect 3430 13574 3476 13626
rect 3180 13572 3236 13574
rect 3260 13572 3316 13574
rect 3340 13572 3396 13574
rect 3420 13572 3476 13574
rect 3180 12538 3236 12540
rect 3260 12538 3316 12540
rect 3340 12538 3396 12540
rect 3420 12538 3476 12540
rect 3180 12486 3226 12538
rect 3226 12486 3236 12538
rect 3260 12486 3290 12538
rect 3290 12486 3302 12538
rect 3302 12486 3316 12538
rect 3340 12486 3354 12538
rect 3354 12486 3366 12538
rect 3366 12486 3396 12538
rect 3420 12486 3430 12538
rect 3430 12486 3476 12538
rect 3180 12484 3236 12486
rect 3260 12484 3316 12486
rect 3340 12484 3396 12486
rect 3420 12484 3476 12486
rect 3238 12144 3294 12200
rect 2870 11056 2926 11112
rect 2778 10920 2834 10976
rect 2226 8084 2282 8120
rect 2226 8064 2228 8084
rect 2228 8064 2280 8084
rect 2280 8064 2282 8084
rect 2226 7656 2282 7712
rect 2226 7384 2282 7440
rect 2778 9696 2834 9752
rect 2594 7520 2650 7576
rect 2042 6568 2098 6624
rect 1766 5616 1822 5672
rect 1674 3984 1730 4040
rect 1490 3168 1546 3224
rect 1674 2352 1730 2408
rect 2870 9288 2926 9344
rect 2594 7112 2650 7168
rect 2594 6996 2650 7032
rect 2594 6976 2596 6996
rect 2596 6976 2648 6996
rect 2648 6976 2650 6996
rect 2594 6704 2650 6760
rect 2410 6432 2466 6488
rect 2134 4684 2190 4720
rect 2134 4664 2136 4684
rect 2136 4664 2188 4684
rect 2188 4664 2190 4684
rect 2226 4392 2282 4448
rect 1858 3576 1914 3632
rect 3180 11450 3236 11452
rect 3260 11450 3316 11452
rect 3340 11450 3396 11452
rect 3420 11450 3476 11452
rect 3180 11398 3226 11450
rect 3226 11398 3236 11450
rect 3260 11398 3290 11450
rect 3290 11398 3302 11450
rect 3302 11398 3316 11450
rect 3340 11398 3354 11450
rect 3354 11398 3366 11450
rect 3366 11398 3396 11450
rect 3420 11398 3430 11450
rect 3430 11398 3476 11450
rect 3180 11396 3236 11398
rect 3260 11396 3316 11398
rect 3340 11396 3396 11398
rect 3420 11396 3476 11398
rect 3054 11192 3110 11248
rect 3422 10920 3478 10976
rect 3180 10362 3236 10364
rect 3260 10362 3316 10364
rect 3340 10362 3396 10364
rect 3420 10362 3476 10364
rect 3180 10310 3226 10362
rect 3226 10310 3236 10362
rect 3260 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3316 10362
rect 3340 10310 3354 10362
rect 3354 10310 3366 10362
rect 3366 10310 3396 10362
rect 3420 10310 3430 10362
rect 3430 10310 3476 10362
rect 3180 10308 3236 10310
rect 3260 10308 3316 10310
rect 3340 10308 3396 10310
rect 3420 10308 3476 10310
rect 3054 10124 3110 10160
rect 3054 10104 3056 10124
rect 3056 10104 3108 10124
rect 3108 10104 3110 10124
rect 2962 8780 2964 8800
rect 2964 8780 3016 8800
rect 3016 8780 3018 8800
rect 2962 8744 3018 8780
rect 2686 6296 2742 6352
rect 3146 9424 3202 9480
rect 4158 13368 4214 13424
rect 4066 11736 4122 11792
rect 3882 11500 3884 11520
rect 3884 11500 3936 11520
rect 3936 11500 3938 11520
rect 3882 11464 3938 11500
rect 3698 9696 3754 9752
rect 3180 9274 3236 9276
rect 3260 9274 3316 9276
rect 3340 9274 3396 9276
rect 3420 9274 3476 9276
rect 3180 9222 3226 9274
rect 3226 9222 3236 9274
rect 3260 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3316 9274
rect 3340 9222 3354 9274
rect 3354 9222 3366 9274
rect 3366 9222 3396 9274
rect 3420 9222 3430 9274
rect 3430 9222 3476 9274
rect 3180 9220 3236 9222
rect 3260 9220 3316 9222
rect 3340 9220 3396 9222
rect 3420 9220 3476 9222
rect 3422 8372 3424 8392
rect 3424 8372 3476 8392
rect 3476 8372 3478 8392
rect 3422 8336 3478 8372
rect 3180 8186 3236 8188
rect 3260 8186 3316 8188
rect 3340 8186 3396 8188
rect 3420 8186 3476 8188
rect 3180 8134 3226 8186
rect 3226 8134 3236 8186
rect 3260 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3316 8186
rect 3340 8134 3354 8186
rect 3354 8134 3366 8186
rect 3366 8134 3396 8186
rect 3420 8134 3430 8186
rect 3430 8134 3476 8186
rect 3180 8132 3236 8134
rect 3260 8132 3316 8134
rect 3340 8132 3396 8134
rect 3420 8132 3476 8134
rect 3422 7928 3478 7984
rect 3422 7384 3478 7440
rect 3330 7248 3386 7304
rect 2962 6976 3018 7032
rect 3180 7098 3236 7100
rect 3260 7098 3316 7100
rect 3340 7098 3396 7100
rect 3420 7098 3476 7100
rect 3180 7046 3226 7098
rect 3226 7046 3236 7098
rect 3260 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3316 7098
rect 3340 7046 3354 7098
rect 3354 7046 3366 7098
rect 3366 7046 3396 7098
rect 3420 7046 3430 7098
rect 3430 7046 3476 7098
rect 3180 7044 3236 7046
rect 3260 7044 3316 7046
rect 3340 7044 3396 7046
rect 3420 7044 3476 7046
rect 3422 6196 3424 6216
rect 3424 6196 3476 6216
rect 3476 6196 3478 6216
rect 3422 6160 3478 6196
rect 1950 2760 2006 2816
rect 1766 1944 1822 2000
rect 1490 1536 1546 1592
rect 1398 1128 1454 1184
rect 3180 6010 3236 6012
rect 3260 6010 3316 6012
rect 3340 6010 3396 6012
rect 3420 6010 3476 6012
rect 3180 5958 3226 6010
rect 3226 5958 3236 6010
rect 3260 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3316 6010
rect 3340 5958 3354 6010
rect 3354 5958 3366 6010
rect 3366 5958 3396 6010
rect 3420 5958 3430 6010
rect 3430 5958 3476 6010
rect 3180 5956 3236 5958
rect 3260 5956 3316 5958
rect 3340 5956 3396 5958
rect 3420 5956 3476 5958
rect 2962 4800 3018 4856
rect 3180 4922 3236 4924
rect 3260 4922 3316 4924
rect 3340 4922 3396 4924
rect 3420 4922 3476 4924
rect 3180 4870 3226 4922
rect 3226 4870 3236 4922
rect 3260 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3316 4922
rect 3340 4870 3354 4922
rect 3354 4870 3366 4922
rect 3366 4870 3396 4922
rect 3420 4870 3430 4922
rect 3430 4870 3476 4922
rect 3180 4868 3236 4870
rect 3260 4868 3316 4870
rect 3340 4868 3396 4870
rect 3420 4868 3476 4870
rect 2778 4120 2834 4176
rect 3180 3834 3236 3836
rect 3260 3834 3316 3836
rect 3340 3834 3396 3836
rect 3420 3834 3476 3836
rect 3180 3782 3226 3834
rect 3226 3782 3236 3834
rect 3260 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3316 3834
rect 3340 3782 3354 3834
rect 3354 3782 3366 3834
rect 3366 3782 3396 3834
rect 3420 3782 3430 3834
rect 3430 3782 3476 3834
rect 3180 3780 3236 3782
rect 3260 3780 3316 3782
rect 3340 3780 3396 3782
rect 3420 3780 3476 3782
rect 3606 8200 3662 8256
rect 3606 3440 3662 3496
rect 2502 2488 2558 2544
rect 3330 3052 3386 3088
rect 5404 14170 5460 14172
rect 5484 14170 5540 14172
rect 5564 14170 5620 14172
rect 5644 14170 5700 14172
rect 5404 14118 5450 14170
rect 5450 14118 5460 14170
rect 5484 14118 5514 14170
rect 5514 14118 5526 14170
rect 5526 14118 5540 14170
rect 5564 14118 5578 14170
rect 5578 14118 5590 14170
rect 5590 14118 5620 14170
rect 5644 14118 5654 14170
rect 5654 14118 5700 14170
rect 5404 14116 5460 14118
rect 5484 14116 5540 14118
rect 5564 14116 5620 14118
rect 5644 14116 5700 14118
rect 4066 10920 4122 10976
rect 4066 9696 4122 9752
rect 3974 8880 4030 8936
rect 3790 7520 3846 7576
rect 3790 6160 3846 6216
rect 3330 3032 3332 3052
rect 3332 3032 3384 3052
rect 3384 3032 3386 3052
rect 3180 2746 3236 2748
rect 3260 2746 3316 2748
rect 3340 2746 3396 2748
rect 3420 2746 3476 2748
rect 3180 2694 3226 2746
rect 3226 2694 3236 2746
rect 3260 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3316 2746
rect 3340 2694 3354 2746
rect 3354 2694 3366 2746
rect 3366 2694 3396 2746
rect 3420 2694 3430 2746
rect 3430 2694 3476 2746
rect 3180 2692 3236 2694
rect 3260 2692 3316 2694
rect 3340 2692 3396 2694
rect 3420 2692 3476 2694
rect 4066 6840 4122 6896
rect 4434 8200 4490 8256
rect 4250 7692 4252 7712
rect 4252 7692 4304 7712
rect 4304 7692 4306 7712
rect 4250 7656 4306 7692
rect 2778 312 2834 368
rect 4342 6740 4344 6760
rect 4344 6740 4396 6760
rect 4396 6740 4398 6760
rect 4342 6704 4398 6740
rect 4802 12164 4858 12200
rect 4802 12144 4804 12164
rect 4804 12144 4856 12164
rect 4856 12144 4858 12164
rect 4986 12144 5042 12200
rect 5404 13082 5460 13084
rect 5484 13082 5540 13084
rect 5564 13082 5620 13084
rect 5644 13082 5700 13084
rect 5404 13030 5450 13082
rect 5450 13030 5460 13082
rect 5484 13030 5514 13082
rect 5514 13030 5526 13082
rect 5526 13030 5540 13082
rect 5564 13030 5578 13082
rect 5578 13030 5590 13082
rect 5590 13030 5620 13082
rect 5644 13030 5654 13082
rect 5654 13030 5700 13082
rect 5404 13028 5460 13030
rect 5484 13028 5540 13030
rect 5564 13028 5620 13030
rect 5644 13028 5700 13030
rect 5814 12416 5870 12472
rect 5404 11994 5460 11996
rect 5484 11994 5540 11996
rect 5564 11994 5620 11996
rect 5644 11994 5700 11996
rect 5404 11942 5450 11994
rect 5450 11942 5460 11994
rect 5484 11942 5514 11994
rect 5514 11942 5526 11994
rect 5526 11942 5540 11994
rect 5564 11942 5578 11994
rect 5578 11942 5590 11994
rect 5590 11942 5620 11994
rect 5644 11942 5654 11994
rect 5654 11942 5700 11994
rect 5404 11940 5460 11942
rect 5484 11940 5540 11942
rect 5564 11940 5620 11942
rect 5644 11940 5700 11942
rect 4710 10668 4766 10704
rect 4710 10648 4712 10668
rect 4712 10648 4764 10668
rect 4764 10648 4766 10668
rect 4710 10376 4766 10432
rect 4526 7520 4582 7576
rect 4618 6840 4674 6896
rect 4894 10104 4950 10160
rect 5404 10906 5460 10908
rect 5484 10906 5540 10908
rect 5564 10906 5620 10908
rect 5644 10906 5700 10908
rect 5404 10854 5450 10906
rect 5450 10854 5460 10906
rect 5484 10854 5514 10906
rect 5514 10854 5526 10906
rect 5526 10854 5540 10906
rect 5564 10854 5578 10906
rect 5578 10854 5590 10906
rect 5590 10854 5620 10906
rect 5644 10854 5654 10906
rect 5654 10854 5700 10906
rect 5404 10852 5460 10854
rect 5484 10852 5540 10854
rect 5564 10852 5620 10854
rect 5644 10852 5700 10854
rect 5354 10548 5356 10568
rect 5356 10548 5408 10568
rect 5408 10548 5410 10568
rect 5354 10512 5410 10548
rect 5538 10240 5594 10296
rect 5446 9968 5502 10024
rect 5404 9818 5460 9820
rect 5484 9818 5540 9820
rect 5564 9818 5620 9820
rect 5644 9818 5700 9820
rect 5404 9766 5450 9818
rect 5450 9766 5460 9818
rect 5484 9766 5514 9818
rect 5514 9766 5526 9818
rect 5526 9766 5540 9818
rect 5564 9766 5578 9818
rect 5578 9766 5590 9818
rect 5590 9766 5620 9818
rect 5644 9766 5654 9818
rect 5654 9766 5700 9818
rect 5404 9764 5460 9766
rect 5484 9764 5540 9766
rect 5564 9764 5620 9766
rect 5644 9764 5700 9766
rect 6274 12008 6330 12064
rect 7628 14714 7684 14716
rect 7708 14714 7764 14716
rect 7788 14714 7844 14716
rect 7868 14714 7924 14716
rect 7628 14662 7674 14714
rect 7674 14662 7684 14714
rect 7708 14662 7738 14714
rect 7738 14662 7750 14714
rect 7750 14662 7764 14714
rect 7788 14662 7802 14714
rect 7802 14662 7814 14714
rect 7814 14662 7844 14714
rect 7868 14662 7878 14714
rect 7878 14662 7924 14714
rect 7628 14660 7684 14662
rect 7708 14660 7764 14662
rect 7788 14660 7844 14662
rect 7868 14660 7924 14662
rect 6366 11772 6368 11792
rect 6368 11772 6420 11792
rect 6420 11772 6422 11792
rect 4986 9424 5042 9480
rect 5078 8780 5080 8800
rect 5080 8780 5132 8800
rect 5132 8780 5134 8800
rect 5078 8744 5134 8780
rect 4986 8608 5042 8664
rect 4802 6840 4858 6896
rect 4434 5636 4490 5672
rect 4434 5616 4436 5636
rect 4436 5616 4488 5636
rect 4488 5616 4490 5636
rect 4158 4020 4160 4040
rect 4160 4020 4212 4040
rect 4212 4020 4214 4040
rect 4158 3984 4214 4020
rect 5538 8880 5594 8936
rect 5814 8900 5870 8936
rect 5814 8880 5816 8900
rect 5816 8880 5868 8900
rect 5868 8880 5870 8900
rect 5998 9016 6054 9072
rect 5404 8730 5460 8732
rect 5484 8730 5540 8732
rect 5564 8730 5620 8732
rect 5644 8730 5700 8732
rect 5404 8678 5450 8730
rect 5450 8678 5460 8730
rect 5484 8678 5514 8730
rect 5514 8678 5526 8730
rect 5526 8678 5540 8730
rect 5564 8678 5578 8730
rect 5578 8678 5590 8730
rect 5590 8678 5620 8730
rect 5644 8678 5654 8730
rect 5654 8678 5700 8730
rect 5404 8676 5460 8678
rect 5484 8676 5540 8678
rect 5564 8676 5620 8678
rect 5644 8676 5700 8678
rect 5906 8744 5962 8800
rect 5630 7964 5632 7984
rect 5632 7964 5684 7984
rect 5684 7964 5686 7984
rect 5630 7928 5686 7964
rect 5404 7642 5460 7644
rect 5484 7642 5540 7644
rect 5564 7642 5620 7644
rect 5644 7642 5700 7644
rect 5404 7590 5450 7642
rect 5450 7590 5460 7642
rect 5484 7590 5514 7642
rect 5514 7590 5526 7642
rect 5526 7590 5540 7642
rect 5564 7590 5578 7642
rect 5578 7590 5590 7642
rect 5590 7590 5620 7642
rect 5644 7590 5654 7642
rect 5654 7590 5700 7642
rect 5404 7588 5460 7590
rect 5484 7588 5540 7590
rect 5564 7588 5620 7590
rect 5644 7588 5700 7590
rect 5170 7384 5226 7440
rect 5630 7404 5686 7440
rect 5630 7384 5632 7404
rect 5632 7384 5684 7404
rect 5684 7384 5686 7404
rect 5630 7112 5686 7168
rect 5538 6976 5594 7032
rect 5404 6554 5460 6556
rect 5484 6554 5540 6556
rect 5564 6554 5620 6556
rect 5644 6554 5700 6556
rect 5404 6502 5450 6554
rect 5450 6502 5460 6554
rect 5484 6502 5514 6554
rect 5514 6502 5526 6554
rect 5526 6502 5540 6554
rect 5564 6502 5578 6554
rect 5578 6502 5590 6554
rect 5590 6502 5620 6554
rect 5644 6502 5654 6554
rect 5654 6502 5700 6554
rect 5404 6500 5460 6502
rect 5484 6500 5540 6502
rect 5564 6500 5620 6502
rect 5644 6500 5700 6502
rect 5404 5466 5460 5468
rect 5484 5466 5540 5468
rect 5564 5466 5620 5468
rect 5644 5466 5700 5468
rect 5404 5414 5450 5466
rect 5450 5414 5460 5466
rect 5484 5414 5514 5466
rect 5514 5414 5526 5466
rect 5526 5414 5540 5466
rect 5564 5414 5578 5466
rect 5578 5414 5590 5466
rect 5590 5414 5620 5466
rect 5644 5414 5654 5466
rect 5654 5414 5700 5466
rect 5404 5412 5460 5414
rect 5484 5412 5540 5414
rect 5564 5412 5620 5414
rect 5644 5412 5700 5414
rect 6366 11736 6422 11772
rect 6458 11056 6514 11112
rect 6274 9696 6330 9752
rect 6090 5616 6146 5672
rect 5404 4378 5460 4380
rect 5484 4378 5540 4380
rect 5564 4378 5620 4380
rect 5644 4378 5700 4380
rect 5404 4326 5450 4378
rect 5450 4326 5460 4378
rect 5484 4326 5514 4378
rect 5514 4326 5526 4378
rect 5526 4326 5540 4378
rect 5564 4326 5578 4378
rect 5578 4326 5590 4378
rect 5590 4326 5620 4378
rect 5644 4326 5654 4378
rect 5654 4326 5700 4378
rect 5404 4324 5460 4326
rect 5484 4324 5540 4326
rect 5564 4324 5620 4326
rect 5644 4324 5700 4326
rect 6734 9560 6790 9616
rect 7628 13626 7684 13628
rect 7708 13626 7764 13628
rect 7788 13626 7844 13628
rect 7868 13626 7924 13628
rect 7628 13574 7674 13626
rect 7674 13574 7684 13626
rect 7708 13574 7738 13626
rect 7738 13574 7750 13626
rect 7750 13574 7764 13626
rect 7788 13574 7802 13626
rect 7802 13574 7814 13626
rect 7814 13574 7844 13626
rect 7868 13574 7878 13626
rect 7878 13574 7924 13626
rect 7628 13572 7684 13574
rect 7708 13572 7764 13574
rect 7788 13572 7844 13574
rect 7868 13572 7924 13574
rect 7194 11464 7250 11520
rect 6826 8608 6882 8664
rect 6458 3984 6514 4040
rect 6274 3440 6330 3496
rect 5404 3290 5460 3292
rect 5484 3290 5540 3292
rect 5564 3290 5620 3292
rect 5644 3290 5700 3292
rect 5404 3238 5450 3290
rect 5450 3238 5460 3290
rect 5484 3238 5514 3290
rect 5514 3238 5526 3290
rect 5526 3238 5540 3290
rect 5564 3238 5578 3290
rect 5578 3238 5590 3290
rect 5590 3238 5620 3290
rect 5644 3238 5654 3290
rect 5654 3238 5700 3290
rect 5404 3236 5460 3238
rect 5484 3236 5540 3238
rect 5564 3236 5620 3238
rect 5644 3236 5700 3238
rect 4802 2352 4858 2408
rect 6090 3052 6146 3088
rect 6090 3032 6092 3052
rect 6092 3032 6144 3052
rect 6144 3032 6146 3052
rect 6918 7112 6974 7168
rect 6826 6296 6882 6352
rect 7562 12688 7618 12744
rect 7628 12538 7684 12540
rect 7708 12538 7764 12540
rect 7788 12538 7844 12540
rect 7868 12538 7924 12540
rect 7628 12486 7674 12538
rect 7674 12486 7684 12538
rect 7708 12486 7738 12538
rect 7738 12486 7750 12538
rect 7750 12486 7764 12538
rect 7788 12486 7802 12538
rect 7802 12486 7814 12538
rect 7814 12486 7844 12538
rect 7868 12486 7878 12538
rect 7878 12486 7924 12538
rect 7628 12484 7684 12486
rect 7708 12484 7764 12486
rect 7788 12484 7844 12486
rect 7868 12484 7924 12486
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9898 14170
rect 9898 14118 9908 14170
rect 9932 14118 9962 14170
rect 9962 14118 9974 14170
rect 9974 14118 9988 14170
rect 10012 14118 10026 14170
rect 10026 14118 10038 14170
rect 10038 14118 10068 14170
rect 10092 14118 10102 14170
rect 10102 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 8114 13232 8170 13288
rect 8022 12416 8078 12472
rect 7654 12044 7656 12064
rect 7656 12044 7708 12064
rect 7708 12044 7710 12064
rect 7654 12008 7710 12044
rect 7194 10376 7250 10432
rect 7194 10240 7250 10296
rect 7286 8608 7342 8664
rect 7746 11600 7802 11656
rect 7628 11450 7684 11452
rect 7708 11450 7764 11452
rect 7788 11450 7844 11452
rect 7868 11450 7924 11452
rect 7628 11398 7674 11450
rect 7674 11398 7684 11450
rect 7708 11398 7738 11450
rect 7738 11398 7750 11450
rect 7750 11398 7764 11450
rect 7788 11398 7802 11450
rect 7802 11398 7814 11450
rect 7814 11398 7844 11450
rect 7868 11398 7878 11450
rect 7878 11398 7924 11450
rect 7628 11396 7684 11398
rect 7708 11396 7764 11398
rect 7788 11396 7844 11398
rect 7868 11396 7924 11398
rect 8022 11092 8024 11112
rect 8024 11092 8076 11112
rect 8076 11092 8078 11112
rect 8022 11056 8078 11092
rect 7628 10362 7684 10364
rect 7708 10362 7764 10364
rect 7788 10362 7844 10364
rect 7868 10362 7924 10364
rect 7628 10310 7674 10362
rect 7674 10310 7684 10362
rect 7708 10310 7738 10362
rect 7738 10310 7750 10362
rect 7750 10310 7764 10362
rect 7788 10310 7802 10362
rect 7802 10310 7814 10362
rect 7814 10310 7844 10362
rect 7868 10310 7878 10362
rect 7878 10310 7924 10362
rect 7628 10308 7684 10310
rect 7708 10308 7764 10310
rect 7788 10308 7844 10310
rect 7868 10308 7924 10310
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9898 13082
rect 9898 13030 9908 13082
rect 9932 13030 9962 13082
rect 9962 13030 9974 13082
rect 9974 13030 9988 13082
rect 10012 13030 10026 13082
rect 10026 13030 10038 13082
rect 10038 13030 10068 13082
rect 10092 13030 10102 13082
rect 10102 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 10230 12300 10286 12336
rect 10230 12280 10232 12300
rect 10232 12280 10284 12300
rect 10284 12280 10286 12300
rect 10506 12144 10562 12200
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9898 11994
rect 9898 11942 9908 11994
rect 9932 11942 9962 11994
rect 9962 11942 9974 11994
rect 9974 11942 9988 11994
rect 10012 11942 10026 11994
rect 10026 11942 10038 11994
rect 10038 11942 10068 11994
rect 10092 11942 10102 11994
rect 10102 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 8022 9832 8078 9888
rect 7654 9580 7710 9616
rect 7654 9560 7656 9580
rect 7656 9560 7708 9580
rect 7708 9560 7710 9580
rect 7628 9274 7684 9276
rect 7708 9274 7764 9276
rect 7788 9274 7844 9276
rect 7868 9274 7924 9276
rect 7628 9222 7674 9274
rect 7674 9222 7684 9274
rect 7708 9222 7738 9274
rect 7738 9222 7750 9274
rect 7750 9222 7764 9274
rect 7788 9222 7802 9274
rect 7802 9222 7814 9274
rect 7814 9222 7844 9274
rect 7868 9222 7878 9274
rect 7878 9222 7924 9274
rect 7628 9220 7684 9222
rect 7708 9220 7764 9222
rect 7788 9220 7844 9222
rect 7868 9220 7924 9222
rect 7562 8608 7618 8664
rect 7562 8336 7618 8392
rect 7628 8186 7684 8188
rect 7708 8186 7764 8188
rect 7788 8186 7844 8188
rect 7868 8186 7924 8188
rect 7628 8134 7674 8186
rect 7674 8134 7684 8186
rect 7708 8134 7738 8186
rect 7738 8134 7750 8186
rect 7750 8134 7764 8186
rect 7788 8134 7802 8186
rect 7802 8134 7814 8186
rect 7814 8134 7844 8186
rect 7868 8134 7878 8186
rect 7878 8134 7924 8186
rect 7628 8132 7684 8134
rect 7708 8132 7764 8134
rect 7788 8132 7844 8134
rect 7868 8132 7924 8134
rect 7628 7098 7684 7100
rect 7708 7098 7764 7100
rect 7788 7098 7844 7100
rect 7868 7098 7924 7100
rect 7628 7046 7674 7098
rect 7674 7046 7684 7098
rect 7708 7046 7738 7098
rect 7738 7046 7750 7098
rect 7750 7046 7764 7098
rect 7788 7046 7802 7098
rect 7802 7046 7814 7098
rect 7814 7046 7844 7098
rect 7868 7046 7878 7098
rect 7878 7046 7924 7098
rect 7628 7044 7684 7046
rect 7708 7044 7764 7046
rect 7788 7044 7844 7046
rect 7868 7044 7924 7046
rect 8298 9324 8300 9344
rect 8300 9324 8352 9344
rect 8352 9324 8354 9344
rect 8298 9288 8354 9324
rect 7628 6010 7684 6012
rect 7708 6010 7764 6012
rect 7788 6010 7844 6012
rect 7868 6010 7924 6012
rect 7628 5958 7674 6010
rect 7674 5958 7684 6010
rect 7708 5958 7738 6010
rect 7738 5958 7750 6010
rect 7750 5958 7764 6010
rect 7788 5958 7802 6010
rect 7802 5958 7814 6010
rect 7814 5958 7844 6010
rect 7868 5958 7878 6010
rect 7878 5958 7924 6010
rect 7628 5956 7684 5958
rect 7708 5956 7764 5958
rect 7788 5956 7844 5958
rect 7868 5956 7924 5958
rect 7628 4922 7684 4924
rect 7708 4922 7764 4924
rect 7788 4922 7844 4924
rect 7868 4922 7924 4924
rect 7628 4870 7674 4922
rect 7674 4870 7684 4922
rect 7708 4870 7738 4922
rect 7738 4870 7750 4922
rect 7750 4870 7764 4922
rect 7788 4870 7802 4922
rect 7802 4870 7814 4922
rect 7814 4870 7844 4922
rect 7868 4870 7878 4922
rect 7878 4870 7924 4922
rect 7628 4868 7684 4870
rect 7708 4868 7764 4870
rect 7788 4868 7844 4870
rect 7868 4868 7924 4870
rect 6550 3032 6606 3088
rect 5404 2202 5460 2204
rect 5484 2202 5540 2204
rect 5564 2202 5620 2204
rect 5644 2202 5700 2204
rect 5404 2150 5450 2202
rect 5450 2150 5460 2202
rect 5484 2150 5514 2202
rect 5514 2150 5526 2202
rect 5526 2150 5540 2202
rect 5564 2150 5578 2202
rect 5578 2150 5590 2202
rect 5590 2150 5620 2202
rect 5644 2150 5654 2202
rect 5654 2150 5700 2202
rect 5404 2148 5460 2150
rect 5484 2148 5540 2150
rect 5564 2148 5620 2150
rect 5644 2148 5700 2150
rect 6458 2624 6514 2680
rect 7628 3834 7684 3836
rect 7708 3834 7764 3836
rect 7788 3834 7844 3836
rect 7868 3834 7924 3836
rect 7628 3782 7674 3834
rect 7674 3782 7684 3834
rect 7708 3782 7738 3834
rect 7738 3782 7750 3834
rect 7750 3782 7764 3834
rect 7788 3782 7802 3834
rect 7802 3782 7814 3834
rect 7814 3782 7844 3834
rect 7868 3782 7878 3834
rect 7878 3782 7924 3834
rect 7628 3780 7684 3782
rect 7708 3780 7764 3782
rect 7788 3780 7844 3782
rect 7868 3780 7924 3782
rect 7628 2746 7684 2748
rect 7708 2746 7764 2748
rect 7788 2746 7844 2748
rect 7868 2746 7924 2748
rect 7628 2694 7674 2746
rect 7674 2694 7684 2746
rect 7708 2694 7738 2746
rect 7738 2694 7750 2746
rect 7750 2694 7764 2746
rect 7788 2694 7802 2746
rect 7802 2694 7814 2746
rect 7814 2694 7844 2746
rect 7868 2694 7878 2746
rect 7878 2694 7924 2746
rect 7628 2692 7684 2694
rect 7708 2692 7764 2694
rect 7788 2692 7844 2694
rect 7868 2692 7924 2694
rect 8666 10920 8722 10976
rect 8666 10784 8722 10840
rect 8942 9152 8998 9208
rect 9034 9016 9090 9072
rect 8850 8608 8906 8664
rect 8758 8472 8814 8528
rect 8942 6704 8998 6760
rect 8482 3576 8538 3632
rect 7930 2372 7986 2408
rect 7930 2352 7932 2372
rect 7932 2352 7984 2372
rect 7984 2352 7986 2372
rect 9402 10104 9458 10160
rect 9218 9596 9220 9616
rect 9220 9596 9272 9616
rect 9272 9596 9274 9616
rect 9218 9560 9274 9596
rect 9218 9152 9274 9208
rect 9218 8744 9274 8800
rect 9586 10104 9642 10160
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9898 10906
rect 9898 10854 9908 10906
rect 9932 10854 9962 10906
rect 9962 10854 9974 10906
rect 9974 10854 9988 10906
rect 10012 10854 10026 10906
rect 10026 10854 10038 10906
rect 10038 10854 10068 10906
rect 10092 10854 10102 10906
rect 10102 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9586 9696 9642 9752
rect 9586 9288 9642 9344
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9898 9818
rect 9898 9766 9908 9818
rect 9932 9766 9962 9818
rect 9962 9766 9974 9818
rect 9974 9766 9988 9818
rect 10012 9766 10026 9818
rect 10026 9766 10038 9818
rect 10038 9766 10068 9818
rect 10092 9766 10102 9818
rect 10102 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9770 9288 9826 9344
rect 9586 8608 9642 8664
rect 9494 8472 9550 8528
rect 10506 11056 10562 11112
rect 10690 11600 10746 11656
rect 10506 9968 10562 10024
rect 10230 9424 10286 9480
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9898 8730
rect 9898 8678 9908 8730
rect 9932 8678 9962 8730
rect 9962 8678 9974 8730
rect 9974 8678 9988 8730
rect 10012 8678 10026 8730
rect 10026 8678 10038 8730
rect 10038 8678 10068 8730
rect 10092 8678 10102 8730
rect 10102 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9898 7642
rect 9898 7590 9908 7642
rect 9932 7590 9962 7642
rect 9962 7590 9974 7642
rect 9974 7590 9988 7642
rect 10012 7590 10026 7642
rect 10026 7590 10038 7642
rect 10038 7590 10068 7642
rect 10092 7590 10102 7642
rect 10102 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9898 6554
rect 9898 6502 9908 6554
rect 9932 6502 9962 6554
rect 9962 6502 9974 6554
rect 9974 6502 9988 6554
rect 10012 6502 10026 6554
rect 10026 6502 10038 6554
rect 10038 6502 10068 6554
rect 10092 6502 10102 6554
rect 10102 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9898 5466
rect 9898 5414 9908 5466
rect 9932 5414 9962 5466
rect 9962 5414 9974 5466
rect 9974 5414 9988 5466
rect 10012 5414 10026 5466
rect 10026 5414 10038 5466
rect 10038 5414 10068 5466
rect 10092 5414 10102 5466
rect 10102 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9678 5344 9734 5400
rect 9310 3984 9366 4040
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9898 4378
rect 9898 4326 9908 4378
rect 9932 4326 9962 4378
rect 9962 4326 9974 4378
rect 9974 4326 9988 4378
rect 10012 4326 10026 4378
rect 10026 4326 10038 4378
rect 10038 4326 10068 4378
rect 10092 4326 10102 4378
rect 10102 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 9586 3168 9642 3224
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9898 3290
rect 9898 3238 9908 3290
rect 9932 3238 9962 3290
rect 9962 3238 9974 3290
rect 9974 3238 9988 3290
rect 10012 3238 10026 3290
rect 10026 3238 10038 3290
rect 10038 3238 10068 3290
rect 10092 3238 10102 3290
rect 10102 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 10414 9152 10470 9208
rect 10414 8780 10416 8800
rect 10416 8780 10468 8800
rect 10468 8780 10470 8800
rect 10414 8744 10470 8780
rect 10690 8472 10746 8528
rect 10414 6160 10470 6216
rect 10966 12144 11022 12200
rect 11150 11500 11152 11520
rect 11152 11500 11204 11520
rect 11204 11500 11206 11520
rect 11150 11464 11206 11500
rect 12076 14714 12132 14716
rect 12156 14714 12212 14716
rect 12236 14714 12292 14716
rect 12316 14714 12372 14716
rect 12076 14662 12122 14714
rect 12122 14662 12132 14714
rect 12156 14662 12186 14714
rect 12186 14662 12198 14714
rect 12198 14662 12212 14714
rect 12236 14662 12250 14714
rect 12250 14662 12262 14714
rect 12262 14662 12292 14714
rect 12316 14662 12326 14714
rect 12326 14662 12372 14714
rect 12076 14660 12132 14662
rect 12156 14660 12212 14662
rect 12236 14660 12292 14662
rect 12316 14660 12372 14662
rect 12076 13626 12132 13628
rect 12156 13626 12212 13628
rect 12236 13626 12292 13628
rect 12316 13626 12372 13628
rect 12076 13574 12122 13626
rect 12122 13574 12132 13626
rect 12156 13574 12186 13626
rect 12186 13574 12198 13626
rect 12198 13574 12212 13626
rect 12236 13574 12250 13626
rect 12250 13574 12262 13626
rect 12262 13574 12292 13626
rect 12316 13574 12326 13626
rect 12326 13574 12372 13626
rect 12076 13572 12132 13574
rect 12156 13572 12212 13574
rect 12236 13572 12292 13574
rect 12316 13572 12372 13574
rect 12076 12538 12132 12540
rect 12156 12538 12212 12540
rect 12236 12538 12292 12540
rect 12316 12538 12372 12540
rect 12076 12486 12122 12538
rect 12122 12486 12132 12538
rect 12156 12486 12186 12538
rect 12186 12486 12198 12538
rect 12198 12486 12212 12538
rect 12236 12486 12250 12538
rect 12250 12486 12262 12538
rect 12262 12486 12292 12538
rect 12316 12486 12326 12538
rect 12326 12486 12372 12538
rect 12076 12484 12132 12486
rect 12156 12484 12212 12486
rect 12236 12484 12292 12486
rect 12316 12484 12372 12486
rect 11794 11464 11850 11520
rect 12076 11450 12132 11452
rect 12156 11450 12212 11452
rect 12236 11450 12292 11452
rect 12316 11450 12372 11452
rect 12076 11398 12122 11450
rect 12122 11398 12132 11450
rect 12156 11398 12186 11450
rect 12186 11398 12198 11450
rect 12198 11398 12212 11450
rect 12236 11398 12250 11450
rect 12250 11398 12262 11450
rect 12262 11398 12292 11450
rect 12316 11398 12326 11450
rect 12326 11398 12372 11450
rect 12076 11396 12132 11398
rect 12156 11396 12212 11398
rect 12236 11396 12292 11398
rect 12316 11396 12372 11398
rect 11242 4664 11298 4720
rect 11610 7420 11612 7440
rect 11612 7420 11664 7440
rect 11664 7420 11666 7440
rect 11610 7384 11666 7420
rect 11518 3984 11574 4040
rect 12076 10362 12132 10364
rect 12156 10362 12212 10364
rect 12236 10362 12292 10364
rect 12316 10362 12372 10364
rect 12076 10310 12122 10362
rect 12122 10310 12132 10362
rect 12156 10310 12186 10362
rect 12186 10310 12198 10362
rect 12198 10310 12212 10362
rect 12236 10310 12250 10362
rect 12250 10310 12262 10362
rect 12262 10310 12292 10362
rect 12316 10310 12326 10362
rect 12326 10310 12372 10362
rect 12076 10308 12132 10310
rect 12156 10308 12212 10310
rect 12236 10308 12292 10310
rect 12316 10308 12372 10310
rect 15014 15680 15070 15736
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14540 14170 14596 14172
rect 14300 14118 14346 14170
rect 14346 14118 14356 14170
rect 14380 14118 14410 14170
rect 14410 14118 14422 14170
rect 14422 14118 14436 14170
rect 14460 14118 14474 14170
rect 14474 14118 14486 14170
rect 14486 14118 14516 14170
rect 14540 14118 14550 14170
rect 14550 14118 14596 14170
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 14540 14116 14596 14118
rect 13726 13812 13728 13832
rect 13728 13812 13780 13832
rect 13780 13812 13782 13832
rect 13726 13776 13782 13812
rect 14922 14048 14978 14104
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14540 13082 14596 13084
rect 14300 13030 14346 13082
rect 14346 13030 14356 13082
rect 14380 13030 14410 13082
rect 14410 13030 14422 13082
rect 14422 13030 14436 13082
rect 14460 13030 14474 13082
rect 14474 13030 14486 13082
rect 14486 13030 14516 13082
rect 14540 13030 14550 13082
rect 14550 13030 14596 13082
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 14540 13028 14596 13030
rect 15198 15408 15254 15464
rect 15290 15272 15346 15328
rect 15290 14864 15346 14920
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16764 14714 16820 14716
rect 16524 14662 16570 14714
rect 16570 14662 16580 14714
rect 16604 14662 16634 14714
rect 16634 14662 16646 14714
rect 16646 14662 16660 14714
rect 16684 14662 16698 14714
rect 16698 14662 16710 14714
rect 16710 14662 16740 14714
rect 16764 14662 16774 14714
rect 16774 14662 16820 14714
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16764 14660 16820 14662
rect 15198 14456 15254 14512
rect 15290 13232 15346 13288
rect 15198 13132 15200 13152
rect 15200 13132 15252 13152
rect 15252 13132 15254 13152
rect 15198 13096 15254 13132
rect 14922 12316 14924 12336
rect 14924 12316 14976 12336
rect 14976 12316 14978 12336
rect 14922 12280 14978 12316
rect 12070 9460 12072 9480
rect 12072 9460 12124 9480
rect 12124 9460 12126 9480
rect 12070 9424 12126 9460
rect 12076 9274 12132 9276
rect 12156 9274 12212 9276
rect 12236 9274 12292 9276
rect 12316 9274 12372 9276
rect 12076 9222 12122 9274
rect 12122 9222 12132 9274
rect 12156 9222 12186 9274
rect 12186 9222 12198 9274
rect 12198 9222 12212 9274
rect 12236 9222 12250 9274
rect 12250 9222 12262 9274
rect 12262 9222 12292 9274
rect 12316 9222 12326 9274
rect 12326 9222 12372 9274
rect 12076 9220 12132 9222
rect 12156 9220 12212 9222
rect 12236 9220 12292 9222
rect 12316 9220 12372 9222
rect 12438 9052 12440 9072
rect 12440 9052 12492 9072
rect 12492 9052 12494 9072
rect 12438 9016 12494 9052
rect 12076 8186 12132 8188
rect 12156 8186 12212 8188
rect 12236 8186 12292 8188
rect 12316 8186 12372 8188
rect 12076 8134 12122 8186
rect 12122 8134 12132 8186
rect 12156 8134 12186 8186
rect 12186 8134 12198 8186
rect 12198 8134 12212 8186
rect 12236 8134 12250 8186
rect 12250 8134 12262 8186
rect 12262 8134 12292 8186
rect 12316 8134 12326 8186
rect 12326 8134 12372 8186
rect 12076 8132 12132 8134
rect 12156 8132 12212 8134
rect 12236 8132 12292 8134
rect 12316 8132 12372 8134
rect 12076 7098 12132 7100
rect 12156 7098 12212 7100
rect 12236 7098 12292 7100
rect 12316 7098 12372 7100
rect 12076 7046 12122 7098
rect 12122 7046 12132 7098
rect 12156 7046 12186 7098
rect 12186 7046 12198 7098
rect 12198 7046 12212 7098
rect 12236 7046 12250 7098
rect 12250 7046 12262 7098
rect 12262 7046 12292 7098
rect 12316 7046 12326 7098
rect 12326 7046 12372 7098
rect 12076 7044 12132 7046
rect 12156 7044 12212 7046
rect 12236 7044 12292 7046
rect 12316 7044 12372 7046
rect 12898 9696 12954 9752
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14540 11994 14596 11996
rect 14300 11942 14346 11994
rect 14346 11942 14356 11994
rect 14380 11942 14410 11994
rect 14410 11942 14422 11994
rect 14422 11942 14436 11994
rect 14460 11942 14474 11994
rect 14474 11942 14486 11994
rect 14486 11942 14516 11994
rect 14540 11942 14550 11994
rect 14550 11942 14596 11994
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14540 11940 14596 11942
rect 13358 9052 13360 9072
rect 13360 9052 13412 9072
rect 13412 9052 13414 9072
rect 13358 9016 13414 9052
rect 12898 7792 12954 7848
rect 13266 7656 13322 7712
rect 12076 6010 12132 6012
rect 12156 6010 12212 6012
rect 12236 6010 12292 6012
rect 12316 6010 12372 6012
rect 12076 5958 12122 6010
rect 12122 5958 12132 6010
rect 12156 5958 12186 6010
rect 12186 5958 12198 6010
rect 12198 5958 12212 6010
rect 12236 5958 12250 6010
rect 12250 5958 12262 6010
rect 12262 5958 12292 6010
rect 12316 5958 12326 6010
rect 12326 5958 12372 6010
rect 12076 5956 12132 5958
rect 12156 5956 12212 5958
rect 12236 5956 12292 5958
rect 12316 5956 12372 5958
rect 12076 4922 12132 4924
rect 12156 4922 12212 4924
rect 12236 4922 12292 4924
rect 12316 4922 12372 4924
rect 12076 4870 12122 4922
rect 12122 4870 12132 4922
rect 12156 4870 12186 4922
rect 12186 4870 12198 4922
rect 12198 4870 12212 4922
rect 12236 4870 12250 4922
rect 12250 4870 12262 4922
rect 12262 4870 12292 4922
rect 12316 4870 12326 4922
rect 12326 4870 12372 4922
rect 12076 4868 12132 4870
rect 12156 4868 12212 4870
rect 12236 4868 12292 4870
rect 12316 4868 12372 4870
rect 12076 3834 12132 3836
rect 12156 3834 12212 3836
rect 12236 3834 12292 3836
rect 12316 3834 12372 3836
rect 12076 3782 12122 3834
rect 12122 3782 12132 3834
rect 12156 3782 12186 3834
rect 12186 3782 12198 3834
rect 12198 3782 12212 3834
rect 12236 3782 12250 3834
rect 12250 3782 12262 3834
rect 12262 3782 12292 3834
rect 12316 3782 12326 3834
rect 12326 3782 12372 3834
rect 12076 3780 12132 3782
rect 12156 3780 12212 3782
rect 12236 3780 12292 3782
rect 12316 3780 12372 3782
rect 9678 2372 9734 2408
rect 9678 2352 9680 2372
rect 9680 2352 9732 2372
rect 9732 2352 9734 2372
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9898 2202
rect 9898 2150 9908 2202
rect 9932 2150 9962 2202
rect 9962 2150 9974 2202
rect 9974 2150 9988 2202
rect 10012 2150 10026 2202
rect 10026 2150 10038 2202
rect 10038 2150 10068 2202
rect 10092 2150 10102 2202
rect 10102 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 12076 2746 12132 2748
rect 12156 2746 12212 2748
rect 12236 2746 12292 2748
rect 12316 2746 12372 2748
rect 12076 2694 12122 2746
rect 12122 2694 12132 2746
rect 12156 2694 12186 2746
rect 12186 2694 12198 2746
rect 12198 2694 12212 2746
rect 12236 2694 12250 2746
rect 12250 2694 12262 2746
rect 12262 2694 12292 2746
rect 12316 2694 12326 2746
rect 12326 2694 12372 2746
rect 12076 2692 12132 2694
rect 12156 2692 12212 2694
rect 12236 2692 12292 2694
rect 12316 2692 12372 2694
rect 12346 2488 12402 2544
rect 14830 11600 14886 11656
rect 14462 11328 14518 11384
rect 14186 11228 14188 11248
rect 14188 11228 14240 11248
rect 14240 11228 14242 11248
rect 14186 11192 14242 11228
rect 13542 8744 13598 8800
rect 13266 6704 13322 6760
rect 14738 11192 14794 11248
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14540 10906 14596 10908
rect 14300 10854 14346 10906
rect 14346 10854 14356 10906
rect 14380 10854 14410 10906
rect 14410 10854 14422 10906
rect 14422 10854 14436 10906
rect 14460 10854 14474 10906
rect 14474 10854 14486 10906
rect 14486 10854 14516 10906
rect 14540 10854 14550 10906
rect 14550 10854 14596 10906
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14540 10852 14596 10854
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14540 9818 14596 9820
rect 14300 9766 14346 9818
rect 14346 9766 14356 9818
rect 14380 9766 14410 9818
rect 14410 9766 14422 9818
rect 14422 9766 14436 9818
rect 14460 9766 14474 9818
rect 14474 9766 14486 9818
rect 14486 9766 14516 9818
rect 14540 9766 14550 9818
rect 14550 9766 14596 9818
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14540 9764 14596 9766
rect 15106 12280 15162 12336
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14540 8730 14596 8732
rect 14300 8678 14346 8730
rect 14346 8678 14356 8730
rect 14380 8678 14410 8730
rect 14410 8678 14422 8730
rect 14422 8678 14436 8730
rect 14460 8678 14474 8730
rect 14474 8678 14486 8730
rect 14486 8678 14516 8730
rect 14540 8678 14550 8730
rect 14550 8678 14596 8730
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14540 8676 14596 8678
rect 14830 8780 14832 8800
rect 14832 8780 14884 8800
rect 14884 8780 14886 8800
rect 14830 8744 14886 8780
rect 14922 8356 14978 8392
rect 14922 8336 14924 8356
rect 14924 8336 14976 8356
rect 14976 8336 14978 8356
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14540 7642 14596 7644
rect 14300 7590 14346 7642
rect 14346 7590 14356 7642
rect 14380 7590 14410 7642
rect 14410 7590 14422 7642
rect 14422 7590 14436 7642
rect 14460 7590 14474 7642
rect 14474 7590 14486 7642
rect 14486 7590 14516 7642
rect 14540 7590 14550 7642
rect 14550 7590 14596 7642
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14540 7588 14596 7590
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14540 6554 14596 6556
rect 14300 6502 14346 6554
rect 14346 6502 14356 6554
rect 14380 6502 14410 6554
rect 14410 6502 14422 6554
rect 14422 6502 14436 6554
rect 14460 6502 14474 6554
rect 14474 6502 14486 6554
rect 14486 6502 14516 6554
rect 14540 6502 14550 6554
rect 14550 6502 14596 6554
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 14540 6500 14596 6502
rect 17958 16496 18014 16552
rect 16302 13812 16304 13832
rect 16304 13812 16356 13832
rect 16356 13812 16358 13832
rect 16302 13776 16358 13812
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16764 13626 16820 13628
rect 16524 13574 16570 13626
rect 16570 13574 16580 13626
rect 16604 13574 16634 13626
rect 16634 13574 16646 13626
rect 16646 13574 16660 13626
rect 16684 13574 16698 13626
rect 16698 13574 16710 13626
rect 16710 13574 16740 13626
rect 16764 13574 16774 13626
rect 16774 13574 16820 13626
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16764 13572 16820 13574
rect 17866 13096 17922 13152
rect 16026 12824 16082 12880
rect 15290 9968 15346 10024
rect 15474 7928 15530 7984
rect 15750 7928 15806 7984
rect 15658 7384 15714 7440
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16764 12538 16820 12540
rect 16524 12486 16570 12538
rect 16570 12486 16580 12538
rect 16604 12486 16634 12538
rect 16634 12486 16646 12538
rect 16646 12486 16660 12538
rect 16684 12486 16698 12538
rect 16698 12486 16710 12538
rect 16710 12486 16740 12538
rect 16764 12486 16774 12538
rect 16774 12486 16820 12538
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 16764 12484 16820 12486
rect 16854 11600 16910 11656
rect 15934 8608 15990 8664
rect 15934 8200 15990 8256
rect 15934 7928 15990 7984
rect 15658 6976 15714 7032
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14540 5466 14596 5468
rect 14300 5414 14346 5466
rect 14346 5414 14356 5466
rect 14380 5414 14410 5466
rect 14410 5414 14422 5466
rect 14422 5414 14436 5466
rect 14460 5414 14474 5466
rect 14474 5414 14486 5466
rect 14486 5414 14516 5466
rect 14540 5414 14550 5466
rect 14550 5414 14596 5466
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 14540 5412 14596 5414
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14540 4378 14596 4380
rect 14300 4326 14346 4378
rect 14346 4326 14356 4378
rect 14380 4326 14410 4378
rect 14410 4326 14422 4378
rect 14422 4326 14436 4378
rect 14460 4326 14474 4378
rect 14474 4326 14486 4378
rect 14486 4326 14516 4378
rect 14540 4326 14550 4378
rect 14550 4326 14596 4378
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 14540 4324 14596 4326
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14540 3290 14596 3292
rect 14300 3238 14346 3290
rect 14346 3238 14356 3290
rect 14380 3238 14410 3290
rect 14410 3238 14422 3290
rect 14422 3238 14436 3290
rect 14460 3238 14474 3290
rect 14474 3238 14486 3290
rect 14486 3238 14516 3290
rect 14540 3238 14550 3290
rect 14550 3238 14596 3290
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 14540 3236 14596 3238
rect 14462 3032 14518 3088
rect 14370 2916 14426 2952
rect 14370 2896 14372 2916
rect 14372 2896 14424 2916
rect 14424 2896 14426 2916
rect 15198 5616 15254 5672
rect 15290 3984 15346 4040
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14540 2202 14596 2204
rect 14300 2150 14346 2202
rect 14346 2150 14356 2202
rect 14380 2150 14410 2202
rect 14410 2150 14422 2202
rect 14422 2150 14436 2202
rect 14460 2150 14474 2202
rect 14474 2150 14486 2202
rect 14486 2150 14516 2202
rect 14540 2150 14550 2202
rect 14550 2150 14596 2202
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 14540 2148 14596 2150
rect 16210 10548 16212 10568
rect 16212 10548 16264 10568
rect 16264 10548 16266 10568
rect 16210 10512 16266 10548
rect 16210 10104 16266 10160
rect 16210 8880 16266 8936
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16764 11450 16820 11452
rect 16524 11398 16570 11450
rect 16570 11398 16580 11450
rect 16604 11398 16634 11450
rect 16634 11398 16646 11450
rect 16646 11398 16660 11450
rect 16684 11398 16698 11450
rect 16698 11398 16710 11450
rect 16710 11398 16740 11450
rect 16764 11398 16774 11450
rect 16774 11398 16820 11450
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16764 11396 16820 11398
rect 17130 11736 17186 11792
rect 16946 11056 17002 11112
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16764 10362 16820 10364
rect 16524 10310 16570 10362
rect 16570 10310 16580 10362
rect 16604 10310 16634 10362
rect 16634 10310 16646 10362
rect 16646 10310 16660 10362
rect 16684 10310 16698 10362
rect 16698 10310 16710 10362
rect 16710 10310 16740 10362
rect 16764 10310 16774 10362
rect 16774 10310 16820 10362
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16764 10308 16820 10310
rect 16394 9968 16450 10024
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16764 9274 16820 9276
rect 16524 9222 16570 9274
rect 16570 9222 16580 9274
rect 16604 9222 16634 9274
rect 16634 9222 16646 9274
rect 16646 9222 16660 9274
rect 16684 9222 16698 9274
rect 16698 9222 16710 9274
rect 16710 9222 16740 9274
rect 16764 9222 16774 9274
rect 16774 9222 16820 9274
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16764 9220 16820 9222
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16764 8186 16820 8188
rect 16524 8134 16570 8186
rect 16570 8134 16580 8186
rect 16604 8134 16634 8186
rect 16634 8134 16646 8186
rect 16646 8134 16660 8186
rect 16684 8134 16698 8186
rect 16698 8134 16710 8186
rect 16710 8134 16740 8186
rect 16764 8134 16774 8186
rect 16774 8134 16820 8186
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16764 8132 16820 8134
rect 17038 10376 17094 10432
rect 17038 9288 17094 9344
rect 17222 9424 17278 9480
rect 17130 8608 17186 8664
rect 17038 8336 17094 8392
rect 16302 7248 16358 7304
rect 16854 7792 16910 7848
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16764 7098 16820 7100
rect 16524 7046 16570 7098
rect 16570 7046 16580 7098
rect 16604 7046 16634 7098
rect 16634 7046 16646 7098
rect 16646 7046 16660 7098
rect 16684 7046 16698 7098
rect 16698 7046 16710 7098
rect 16710 7046 16740 7098
rect 16764 7046 16774 7098
rect 16774 7046 16820 7098
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16764 7044 16820 7046
rect 16486 6704 16542 6760
rect 16210 5616 16266 5672
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16764 6010 16820 6012
rect 16524 5958 16570 6010
rect 16570 5958 16580 6010
rect 16604 5958 16634 6010
rect 16634 5958 16646 6010
rect 16646 5958 16660 6010
rect 16684 5958 16698 6010
rect 16698 5958 16710 6010
rect 16710 5958 16740 6010
rect 16764 5958 16774 6010
rect 16774 5958 16820 6010
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 16764 5956 16820 5958
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16764 4922 16820 4924
rect 16524 4870 16570 4922
rect 16570 4870 16580 4922
rect 16604 4870 16634 4922
rect 16634 4870 16646 4922
rect 16646 4870 16660 4922
rect 16684 4870 16698 4922
rect 16698 4870 16710 4922
rect 16710 4870 16740 4922
rect 16764 4870 16774 4922
rect 16774 4870 16820 4922
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16764 4868 16820 4870
rect 16118 3848 16174 3904
rect 4066 720 4122 776
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16764 3834 16820 3836
rect 16524 3782 16570 3834
rect 16570 3782 16580 3834
rect 16604 3782 16634 3834
rect 16634 3782 16646 3834
rect 16646 3782 16660 3834
rect 16684 3782 16698 3834
rect 16698 3782 16710 3834
rect 16710 3782 16740 3834
rect 16764 3782 16774 3834
rect 16774 3782 16820 3834
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 16764 3780 16820 3782
rect 17222 6740 17224 6760
rect 17224 6740 17276 6760
rect 17276 6740 17278 6760
rect 17222 6704 17278 6740
rect 16946 3576 17002 3632
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16764 2746 16820 2748
rect 16524 2694 16570 2746
rect 16570 2694 16580 2746
rect 16604 2694 16634 2746
rect 16634 2694 16646 2746
rect 16646 2694 16660 2746
rect 16684 2694 16698 2746
rect 16698 2694 16710 2746
rect 16710 2694 16740 2746
rect 16764 2694 16774 2746
rect 16774 2694 16820 2746
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16764 2692 16820 2694
rect 17866 10920 17922 10976
rect 17682 9152 17738 9208
rect 17682 8780 17684 8800
rect 17684 8780 17736 8800
rect 17736 8780 17738 8800
rect 17682 8744 17738 8780
rect 17590 8336 17646 8392
rect 17866 9016 17922 9072
rect 17866 8744 17922 8800
rect 17498 7248 17554 7304
rect 17498 5616 17554 5672
rect 17406 4020 17408 4040
rect 17408 4020 17460 4040
rect 17460 4020 17462 4040
rect 17406 3984 17462 4020
rect 17314 1400 17370 1456
rect 17866 7928 17922 7984
rect 17682 1808 17738 1864
rect 17406 992 17462 1048
rect 18142 9560 18198 9616
rect 18050 8356 18106 8392
rect 18050 8336 18052 8356
rect 18052 8336 18104 8356
rect 18104 8336 18106 8356
rect 18050 7964 18052 7984
rect 18052 7964 18104 7984
rect 18104 7964 18106 7984
rect 18050 7928 18106 7964
rect 18050 7112 18106 7168
rect 18050 6432 18106 6488
rect 17958 5480 18014 5536
rect 18418 7520 18474 7576
rect 18418 6704 18474 6760
rect 18510 6296 18566 6352
rect 18142 4664 18198 4720
rect 18234 3440 18290 3496
rect 18602 5888 18658 5944
rect 18694 5072 18750 5128
rect 18050 3032 18106 3088
rect 17866 2932 17868 2952
rect 17868 2932 17920 2952
rect 17920 2932 17922 2952
rect 17866 2896 17922 2932
rect 18418 2252 18420 2272
rect 18420 2252 18472 2272
rect 18472 2252 18474 2272
rect 18418 2216 18474 2252
rect 18970 10532 19026 10568
rect 18970 10512 18972 10532
rect 18972 10512 19024 10532
rect 19024 10512 19026 10532
rect 18878 4256 18934 4312
rect 18970 3848 19026 3904
rect 18786 2624 18842 2680
rect 16302 584 16358 640
<< metal3 >>
rect 0 16690 800 16720
rect 4429 16690 4495 16693
rect 0 16688 4495 16690
rect 0 16632 4434 16688
rect 4490 16632 4495 16688
rect 0 16630 4495 16632
rect 0 16600 800 16630
rect 4429 16627 4495 16630
rect 17953 16554 18019 16557
rect 19200 16554 20000 16584
rect 17953 16552 20000 16554
rect 17953 16496 17958 16552
rect 18014 16496 20000 16552
rect 17953 16494 20000 16496
rect 17953 16491 18019 16494
rect 19200 16464 20000 16494
rect 0 16282 800 16312
rect 3969 16282 4035 16285
rect 0 16280 4035 16282
rect 0 16224 3974 16280
rect 4030 16224 4035 16280
rect 0 16222 4035 16224
rect 0 16192 800 16222
rect 3969 16219 4035 16222
rect 17718 16084 17724 16148
rect 17788 16146 17794 16148
rect 19200 16146 20000 16176
rect 17788 16086 20000 16146
rect 17788 16084 17794 16086
rect 19200 16056 20000 16086
rect 0 15874 800 15904
rect 4061 15874 4127 15877
rect 0 15872 4127 15874
rect 0 15816 4066 15872
rect 4122 15816 4127 15872
rect 0 15814 4127 15816
rect 0 15784 800 15814
rect 4061 15811 4127 15814
rect 15009 15738 15075 15741
rect 19200 15738 20000 15768
rect 15009 15736 20000 15738
rect 15009 15680 15014 15736
rect 15070 15680 20000 15736
rect 15009 15678 20000 15680
rect 15009 15675 15075 15678
rect 19200 15648 20000 15678
rect 0 15466 800 15496
rect 3417 15466 3483 15469
rect 0 15464 3483 15466
rect 0 15408 3422 15464
rect 3478 15408 3483 15464
rect 0 15406 3483 15408
rect 0 15376 800 15406
rect 3417 15403 3483 15406
rect 15193 15466 15259 15469
rect 17718 15466 17724 15468
rect 15193 15464 17724 15466
rect 15193 15408 15198 15464
rect 15254 15408 17724 15464
rect 15193 15406 17724 15408
rect 15193 15403 15259 15406
rect 17718 15404 17724 15406
rect 17788 15404 17794 15468
rect 15285 15330 15351 15333
rect 19200 15330 20000 15360
rect 15285 15328 20000 15330
rect 15285 15272 15290 15328
rect 15346 15272 20000 15328
rect 15285 15270 20000 15272
rect 15285 15267 15351 15270
rect 19200 15240 20000 15270
rect 0 15058 800 15088
rect 3734 15058 3740 15060
rect 0 14998 3740 15058
rect 0 14968 800 14998
rect 3734 14996 3740 14998
rect 3804 14996 3810 15060
rect 15285 14922 15351 14925
rect 19200 14922 20000 14952
rect 15285 14920 20000 14922
rect 15285 14864 15290 14920
rect 15346 14864 20000 14920
rect 15285 14862 20000 14864
rect 15285 14859 15351 14862
rect 19200 14832 20000 14862
rect 3170 14720 3486 14721
rect 0 14650 800 14680
rect 3170 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3486 14720
rect 3170 14655 3486 14656
rect 7618 14720 7934 14721
rect 7618 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7934 14720
rect 7618 14655 7934 14656
rect 12066 14720 12382 14721
rect 12066 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12382 14720
rect 12066 14655 12382 14656
rect 16514 14720 16830 14721
rect 16514 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16830 14720
rect 16514 14655 16830 14656
rect 2773 14650 2839 14653
rect 0 14648 2839 14650
rect 0 14592 2778 14648
rect 2834 14592 2839 14648
rect 0 14590 2839 14592
rect 0 14560 800 14590
rect 2773 14587 2839 14590
rect 15193 14514 15259 14517
rect 19200 14514 20000 14544
rect 15193 14512 20000 14514
rect 15193 14456 15198 14512
rect 15254 14456 20000 14512
rect 15193 14454 20000 14456
rect 15193 14451 15259 14454
rect 19200 14424 20000 14454
rect 0 14242 800 14272
rect 3509 14242 3575 14245
rect 0 14240 3575 14242
rect 0 14184 3514 14240
rect 3570 14184 3575 14240
rect 0 14182 3575 14184
rect 0 14152 800 14182
rect 3509 14179 3575 14182
rect 5394 14176 5710 14177
rect 5394 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5710 14176
rect 5394 14111 5710 14112
rect 9842 14176 10158 14177
rect 9842 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10158 14176
rect 9842 14111 10158 14112
rect 14290 14176 14606 14177
rect 14290 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14606 14176
rect 14290 14111 14606 14112
rect 14917 14106 14983 14109
rect 19200 14106 20000 14136
rect 14917 14104 20000 14106
rect 14917 14048 14922 14104
rect 14978 14048 20000 14104
rect 14917 14046 20000 14048
rect 14917 14043 14983 14046
rect 19200 14016 20000 14046
rect 4654 13908 4660 13972
rect 4724 13970 4730 13972
rect 4724 13910 6930 13970
rect 4724 13908 4730 13910
rect 0 13834 800 13864
rect 3417 13834 3483 13837
rect 0 13832 3483 13834
rect 0 13776 3422 13832
rect 3478 13776 3483 13832
rect 0 13774 3483 13776
rect 6870 13834 6930 13910
rect 13721 13834 13787 13837
rect 16297 13836 16363 13837
rect 14958 13834 14964 13836
rect 6870 13832 14964 13834
rect 6870 13776 13726 13832
rect 13782 13776 14964 13832
rect 6870 13774 14964 13776
rect 0 13744 800 13774
rect 3417 13771 3483 13774
rect 13721 13771 13787 13774
rect 14958 13772 14964 13774
rect 15028 13772 15034 13836
rect 16246 13772 16252 13836
rect 16316 13834 16363 13836
rect 16316 13832 16408 13834
rect 16358 13776 16408 13832
rect 16316 13774 16408 13776
rect 16316 13772 16363 13774
rect 16297 13771 16363 13772
rect 19200 13698 20000 13728
rect 17910 13638 20000 13698
rect 3170 13632 3486 13633
rect 3170 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3486 13632
rect 3170 13567 3486 13568
rect 7618 13632 7934 13633
rect 7618 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7934 13632
rect 7618 13567 7934 13568
rect 12066 13632 12382 13633
rect 12066 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12382 13632
rect 12066 13567 12382 13568
rect 16514 13632 16830 13633
rect 16514 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16830 13632
rect 16514 13567 16830 13568
rect 0 13426 800 13456
rect 4153 13426 4219 13429
rect 0 13424 4219 13426
rect 0 13368 4158 13424
rect 4214 13368 4219 13424
rect 0 13366 4219 13368
rect 0 13336 800 13366
rect 4153 13363 4219 13366
rect 8109 13290 8175 13293
rect 15285 13290 15351 13293
rect 17910 13290 17970 13638
rect 19200 13608 20000 13638
rect 19200 13290 20000 13320
rect 8109 13288 17970 13290
rect 8109 13232 8114 13288
rect 8170 13232 15290 13288
rect 15346 13232 17970 13288
rect 8109 13230 17970 13232
rect 18278 13230 20000 13290
rect 8109 13227 8175 13230
rect 15285 13227 15351 13230
rect 15193 13156 15259 13157
rect 15142 13092 15148 13156
rect 15212 13154 15259 13156
rect 17861 13154 17927 13157
rect 18278 13154 18338 13230
rect 19200 13200 20000 13230
rect 15212 13152 15304 13154
rect 15254 13096 15304 13152
rect 15212 13094 15304 13096
rect 17861 13152 18338 13154
rect 17861 13096 17866 13152
rect 17922 13096 18338 13152
rect 17861 13094 18338 13096
rect 15212 13092 15259 13094
rect 15193 13091 15259 13092
rect 17861 13091 17927 13094
rect 5394 13088 5710 13089
rect 0 13018 800 13048
rect 5394 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5710 13088
rect 5394 13023 5710 13024
rect 9842 13088 10158 13089
rect 9842 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10158 13088
rect 9842 13023 10158 13024
rect 14290 13088 14606 13089
rect 14290 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14606 13088
rect 14290 13023 14606 13024
rect 1853 13018 1919 13021
rect 0 13016 1919 13018
rect 0 12960 1858 13016
rect 1914 12960 1919 13016
rect 0 12958 1919 12960
rect 0 12928 800 12958
rect 1853 12955 1919 12958
rect 16021 12882 16087 12885
rect 19200 12882 20000 12912
rect 16021 12880 20000 12882
rect 16021 12824 16026 12880
rect 16082 12824 20000 12880
rect 16021 12822 20000 12824
rect 16021 12819 16087 12822
rect 19200 12792 20000 12822
rect 2221 12746 2287 12749
rect 7557 12746 7623 12749
rect 2221 12744 7623 12746
rect 2221 12688 2226 12744
rect 2282 12688 7562 12744
rect 7618 12688 7623 12744
rect 2221 12686 7623 12688
rect 2221 12683 2287 12686
rect 7557 12683 7623 12686
rect 0 12610 800 12640
rect 2773 12610 2839 12613
rect 0 12608 2839 12610
rect 0 12552 2778 12608
rect 2834 12552 2839 12608
rect 0 12550 2839 12552
rect 0 12520 800 12550
rect 2773 12547 2839 12550
rect 3170 12544 3486 12545
rect 3170 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3486 12544
rect 3170 12479 3486 12480
rect 7618 12544 7934 12545
rect 7618 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7934 12544
rect 7618 12479 7934 12480
rect 12066 12544 12382 12545
rect 12066 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12382 12544
rect 12066 12479 12382 12480
rect 16514 12544 16830 12545
rect 16514 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16830 12544
rect 16514 12479 16830 12480
rect 5809 12474 5875 12477
rect 5942 12474 5948 12476
rect 5809 12472 5948 12474
rect 5809 12416 5814 12472
rect 5870 12416 5948 12472
rect 5809 12414 5948 12416
rect 5809 12411 5875 12414
rect 5942 12412 5948 12414
rect 6012 12412 6018 12476
rect 8017 12474 8083 12477
rect 8150 12474 8156 12476
rect 8017 12472 8156 12474
rect 8017 12416 8022 12472
rect 8078 12416 8156 12472
rect 8017 12414 8156 12416
rect 8017 12411 8083 12414
rect 8150 12412 8156 12414
rect 8220 12412 8226 12476
rect 19200 12474 20000 12504
rect 16944 12414 20000 12474
rect 2313 12338 2379 12341
rect 10225 12338 10291 12341
rect 14917 12338 14983 12341
rect 2313 12336 14983 12338
rect 2313 12280 2318 12336
rect 2374 12280 10230 12336
rect 10286 12280 14922 12336
rect 14978 12280 14983 12336
rect 2313 12278 14983 12280
rect 2313 12275 2379 12278
rect 10225 12275 10291 12278
rect 14917 12275 14983 12278
rect 15101 12338 15167 12341
rect 16944 12338 17004 12414
rect 19200 12384 20000 12414
rect 15101 12336 17004 12338
rect 15101 12280 15106 12336
rect 15162 12280 17004 12336
rect 15101 12278 17004 12280
rect 15101 12275 15167 12278
rect 0 12202 800 12232
rect 3233 12202 3299 12205
rect 0 12200 3299 12202
rect 0 12144 3238 12200
rect 3294 12144 3299 12200
rect 0 12142 3299 12144
rect 0 12112 800 12142
rect 3233 12139 3299 12142
rect 3734 12140 3740 12204
rect 3804 12202 3810 12204
rect 4797 12202 4863 12205
rect 3804 12200 4863 12202
rect 3804 12144 4802 12200
rect 4858 12144 4863 12200
rect 3804 12142 4863 12144
rect 3804 12140 3810 12142
rect 4797 12139 4863 12142
rect 4981 12202 5047 12205
rect 10501 12202 10567 12205
rect 4981 12200 10567 12202
rect 4981 12144 4986 12200
rect 5042 12144 10506 12200
rect 10562 12144 10567 12200
rect 4981 12142 10567 12144
rect 4981 12139 5047 12142
rect 10501 12139 10567 12142
rect 10961 12202 11027 12205
rect 10961 12200 15946 12202
rect 10961 12144 10966 12200
rect 11022 12144 15946 12200
rect 10961 12142 15946 12144
rect 10961 12139 11027 12142
rect 6269 12066 6335 12069
rect 7649 12066 7715 12069
rect 15886 12066 15946 12142
rect 19200 12066 20000 12096
rect 6269 12064 9690 12066
rect 6269 12008 6274 12064
rect 6330 12008 7654 12064
rect 7710 12008 9690 12064
rect 6269 12006 9690 12008
rect 15886 12006 20000 12066
rect 6269 12003 6335 12006
rect 7649 12003 7715 12006
rect 5394 12000 5710 12001
rect 5394 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5710 12000
rect 5394 11935 5710 11936
rect 2446 11868 2452 11932
rect 2516 11930 2522 11932
rect 2516 11870 5274 11930
rect 2516 11868 2522 11870
rect 0 11794 800 11824
rect 4061 11794 4127 11797
rect 0 11792 4127 11794
rect 0 11736 4066 11792
rect 4122 11736 4127 11792
rect 0 11734 4127 11736
rect 5214 11794 5274 11870
rect 6361 11794 6427 11797
rect 5214 11792 6427 11794
rect 5214 11736 6366 11792
rect 6422 11736 6427 11792
rect 5214 11734 6427 11736
rect 9630 11794 9690 12006
rect 9842 12000 10158 12001
rect 9842 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10158 12000
rect 9842 11935 10158 11936
rect 14290 12000 14606 12001
rect 14290 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14606 12000
rect 19200 11976 20000 12006
rect 14290 11935 14606 11936
rect 17125 11794 17191 11797
rect 9630 11792 17191 11794
rect 9630 11736 17130 11792
rect 17186 11736 17191 11792
rect 9630 11734 17191 11736
rect 0 11704 800 11734
rect 4061 11731 4127 11734
rect 6361 11731 6427 11734
rect 17125 11731 17191 11734
rect 2497 11658 2563 11661
rect 7741 11658 7807 11661
rect 2497 11656 7807 11658
rect 2497 11600 2502 11656
rect 2558 11600 7746 11656
rect 7802 11600 7807 11656
rect 2497 11598 7807 11600
rect 2497 11595 2563 11598
rect 7741 11595 7807 11598
rect 10685 11658 10751 11661
rect 14825 11658 14891 11661
rect 10685 11656 14891 11658
rect 10685 11600 10690 11656
rect 10746 11600 14830 11656
rect 14886 11600 14891 11656
rect 10685 11598 14891 11600
rect 10685 11595 10751 11598
rect 14825 11595 14891 11598
rect 16849 11658 16915 11661
rect 19200 11658 20000 11688
rect 16849 11656 20000 11658
rect 16849 11600 16854 11656
rect 16910 11600 20000 11656
rect 16849 11598 20000 11600
rect 16849 11595 16915 11598
rect 19200 11568 20000 11598
rect 3877 11522 3943 11525
rect 7189 11522 7255 11525
rect 3877 11520 7255 11522
rect 3877 11464 3882 11520
rect 3938 11464 7194 11520
rect 7250 11464 7255 11520
rect 3877 11462 7255 11464
rect 3877 11459 3943 11462
rect 7189 11459 7255 11462
rect 11145 11522 11211 11525
rect 11789 11522 11855 11525
rect 11145 11520 11898 11522
rect 11145 11464 11150 11520
rect 11206 11464 11794 11520
rect 11850 11464 11898 11520
rect 11145 11462 11898 11464
rect 11145 11459 11211 11462
rect 11789 11459 11898 11462
rect 3170 11456 3486 11457
rect 0 11386 800 11416
rect 3170 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3486 11456
rect 3170 11391 3486 11392
rect 7618 11456 7934 11457
rect 7618 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7934 11456
rect 7618 11391 7934 11392
rect 1209 11386 1275 11389
rect 0 11384 1275 11386
rect 0 11328 1214 11384
rect 1270 11328 1275 11384
rect 0 11326 1275 11328
rect 0 11296 800 11326
rect 1209 11323 1275 11326
rect 3049 11250 3115 11253
rect 3049 11248 7298 11250
rect 3049 11192 3054 11248
rect 3110 11192 7298 11248
rect 3049 11190 7298 11192
rect 3049 11187 3115 11190
rect 2865 11116 2931 11117
rect 2814 11114 2820 11116
rect 2774 11054 2820 11114
rect 2884 11112 2931 11116
rect 6453 11116 6519 11117
rect 2926 11056 2931 11112
rect 2814 11052 2820 11054
rect 2884 11052 2931 11056
rect 2865 11051 2931 11052
rect 5214 11054 5872 11114
rect 0 10978 800 11008
rect 2773 10978 2839 10981
rect 3417 10978 3483 10981
rect 0 10976 3483 10978
rect 0 10920 2778 10976
rect 2834 10920 3422 10976
rect 3478 10920 3483 10976
rect 0 10918 3483 10920
rect 0 10888 800 10918
rect 2773 10915 2839 10918
rect 3417 10915 3483 10918
rect 4061 10978 4127 10981
rect 5214 10978 5274 11054
rect 4061 10976 5274 10978
rect 4061 10920 4066 10976
rect 4122 10920 5274 10976
rect 4061 10918 5274 10920
rect 4061 10915 4127 10918
rect 5394 10912 5710 10913
rect 5394 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5710 10912
rect 5394 10847 5710 10848
rect 5812 10842 5872 11054
rect 6453 11112 6500 11116
rect 6564 11114 6570 11116
rect 7238 11114 7298 11190
rect 7414 11188 7420 11252
rect 7484 11250 7490 11252
rect 8150 11250 8156 11252
rect 7484 11190 8156 11250
rect 7484 11188 7490 11190
rect 8150 11188 8156 11190
rect 8220 11188 8226 11252
rect 11838 11250 11898 11459
rect 12066 11456 12382 11457
rect 12066 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12382 11456
rect 12066 11391 12382 11392
rect 16514 11456 16830 11457
rect 16514 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16830 11456
rect 16514 11391 16830 11392
rect 14457 11386 14523 11389
rect 14774 11386 14780 11388
rect 14457 11384 14780 11386
rect 14457 11328 14462 11384
rect 14518 11328 14780 11384
rect 14457 11326 14780 11328
rect 14457 11323 14523 11326
rect 14774 11324 14780 11326
rect 14844 11324 14850 11388
rect 14181 11250 14247 11253
rect 11838 11248 14247 11250
rect 11838 11192 14186 11248
rect 14242 11192 14247 11248
rect 11838 11190 14247 11192
rect 14181 11187 14247 11190
rect 14733 11250 14799 11253
rect 19200 11250 20000 11280
rect 14733 11248 20000 11250
rect 14733 11192 14738 11248
rect 14794 11192 20000 11248
rect 14733 11190 20000 11192
rect 14733 11187 14799 11190
rect 19200 11160 20000 11190
rect 8017 11114 8083 11117
rect 8150 11114 8156 11116
rect 6453 11056 6458 11112
rect 6453 11052 6500 11056
rect 6564 11054 6610 11114
rect 7238 11054 7850 11114
rect 6564 11052 6570 11054
rect 6453 11051 6519 11052
rect 7790 10978 7850 11054
rect 8017 11112 8156 11114
rect 8017 11056 8022 11112
rect 8078 11056 8156 11112
rect 8017 11054 8156 11056
rect 8017 11051 8083 11054
rect 8150 11052 8156 11054
rect 8220 11052 8226 11116
rect 10501 11114 10567 11117
rect 16941 11114 17007 11117
rect 10501 11112 17007 11114
rect 10501 11056 10506 11112
rect 10562 11056 16946 11112
rect 17002 11056 17007 11112
rect 10501 11054 17007 11056
rect 10501 11051 10567 11054
rect 16941 11051 17007 11054
rect 8661 10978 8727 10981
rect 17861 10978 17927 10981
rect 7790 10976 8727 10978
rect 7790 10920 8666 10976
rect 8722 10920 8727 10976
rect 7790 10918 8727 10920
rect 8661 10915 8727 10918
rect 15702 10976 17927 10978
rect 15702 10920 17866 10976
rect 17922 10920 17927 10976
rect 15702 10918 17927 10920
rect 9842 10912 10158 10913
rect 9842 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10158 10912
rect 9842 10847 10158 10848
rect 14290 10912 14606 10913
rect 14290 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14606 10912
rect 14290 10847 14606 10848
rect 8661 10842 8727 10845
rect 5812 10840 8727 10842
rect 5812 10784 8666 10840
rect 8722 10784 8727 10840
rect 5812 10782 8727 10784
rect 8661 10779 8727 10782
rect 4705 10706 4771 10709
rect 15702 10706 15762 10918
rect 17861 10915 17927 10918
rect 19200 10842 20000 10872
rect 4705 10704 15762 10706
rect 4705 10648 4710 10704
rect 4766 10648 15762 10704
rect 4705 10646 15762 10648
rect 15886 10782 20000 10842
rect 4705 10643 4771 10646
rect 0 10570 800 10600
rect 1761 10570 1827 10573
rect 0 10568 1827 10570
rect 0 10512 1766 10568
rect 1822 10512 1827 10568
rect 0 10510 1827 10512
rect 0 10480 800 10510
rect 1761 10507 1827 10510
rect 5349 10570 5415 10573
rect 15886 10570 15946 10782
rect 19200 10752 20000 10782
rect 5349 10568 15946 10570
rect 5349 10512 5354 10568
rect 5410 10512 15946 10568
rect 5349 10510 15946 10512
rect 16205 10570 16271 10573
rect 18965 10570 19031 10573
rect 16205 10568 19031 10570
rect 16205 10512 16210 10568
rect 16266 10512 18970 10568
rect 19026 10512 19031 10568
rect 16205 10510 19031 10512
rect 5349 10507 5415 10510
rect 16205 10507 16271 10510
rect 18965 10507 19031 10510
rect 4705 10434 4771 10437
rect 7189 10434 7255 10437
rect 4705 10432 7255 10434
rect 4705 10376 4710 10432
rect 4766 10376 7194 10432
rect 7250 10376 7255 10432
rect 4705 10374 7255 10376
rect 4705 10371 4771 10374
rect 7189 10371 7255 10374
rect 17033 10434 17099 10437
rect 19200 10434 20000 10464
rect 17033 10432 20000 10434
rect 17033 10376 17038 10432
rect 17094 10376 20000 10432
rect 17033 10374 20000 10376
rect 17033 10371 17099 10374
rect 3170 10368 3486 10369
rect 3170 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3486 10368
rect 3170 10303 3486 10304
rect 7618 10368 7934 10369
rect 7618 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7934 10368
rect 7618 10303 7934 10304
rect 12066 10368 12382 10369
rect 12066 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12382 10368
rect 12066 10303 12382 10304
rect 16514 10368 16830 10369
rect 16514 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16830 10368
rect 19200 10344 20000 10374
rect 16514 10303 16830 10304
rect 5533 10298 5599 10301
rect 7189 10298 7255 10301
rect 5533 10296 7255 10298
rect 5533 10240 5538 10296
rect 5594 10240 7194 10296
rect 7250 10240 7255 10296
rect 5533 10238 7255 10240
rect 5533 10235 5599 10238
rect 7189 10235 7255 10238
rect 0 10162 800 10192
rect 1117 10162 1183 10165
rect 3049 10162 3115 10165
rect 0 10160 3115 10162
rect 0 10104 1122 10160
rect 1178 10104 3054 10160
rect 3110 10104 3115 10160
rect 0 10102 3115 10104
rect 0 10072 800 10102
rect 1117 10099 1183 10102
rect 3049 10099 3115 10102
rect 4889 10162 4955 10165
rect 9397 10162 9463 10165
rect 4889 10160 9463 10162
rect 4889 10104 4894 10160
rect 4950 10104 9402 10160
rect 9458 10104 9463 10160
rect 4889 10102 9463 10104
rect 4889 10099 4955 10102
rect 9397 10099 9463 10102
rect 9581 10162 9647 10165
rect 16205 10162 16271 10165
rect 9581 10160 16271 10162
rect 9581 10104 9586 10160
rect 9642 10104 16210 10160
rect 16266 10104 16271 10160
rect 9581 10102 16271 10104
rect 9581 10099 9647 10102
rect 16205 10099 16271 10102
rect 1761 10026 1827 10029
rect 2313 10026 2379 10029
rect 5441 10026 5507 10029
rect 10501 10026 10567 10029
rect 1761 10024 2790 10026
rect 1761 9968 1766 10024
rect 1822 9968 2318 10024
rect 2374 9968 2790 10024
rect 1761 9966 2790 9968
rect 1761 9963 1827 9966
rect 2313 9963 2379 9966
rect 2730 9890 2790 9966
rect 5441 10024 10567 10026
rect 5441 9968 5446 10024
rect 5502 9968 10506 10024
rect 10562 9968 10567 10024
rect 5441 9966 10567 9968
rect 5441 9963 5507 9966
rect 10501 9963 10567 9966
rect 15285 10026 15351 10029
rect 16389 10026 16455 10029
rect 19200 10026 20000 10056
rect 15285 10024 20000 10026
rect 15285 9968 15290 10024
rect 15346 9968 16394 10024
rect 16450 9968 20000 10024
rect 15285 9966 20000 9968
rect 15285 9963 15351 9966
rect 16389 9963 16455 9966
rect 19200 9936 20000 9966
rect 8017 9890 8083 9893
rect 2730 9830 5274 9890
rect 0 9754 800 9784
rect 2773 9754 2839 9757
rect 0 9752 2839 9754
rect 0 9696 2778 9752
rect 2834 9696 2839 9752
rect 0 9694 2839 9696
rect 0 9664 800 9694
rect 2773 9691 2839 9694
rect 3550 9692 3556 9756
rect 3620 9754 3626 9756
rect 3693 9754 3759 9757
rect 3620 9752 3759 9754
rect 3620 9696 3698 9752
rect 3754 9696 3759 9752
rect 3620 9694 3759 9696
rect 3620 9692 3626 9694
rect 3693 9691 3759 9694
rect 4061 9756 4127 9757
rect 4061 9752 4108 9756
rect 4172 9754 4178 9756
rect 4061 9696 4066 9752
rect 4061 9692 4108 9696
rect 4172 9694 4218 9754
rect 4172 9692 4178 9694
rect 4061 9691 4127 9692
rect 5214 9618 5274 9830
rect 5812 9888 8083 9890
rect 5812 9832 8022 9888
rect 8078 9832 8083 9888
rect 5812 9830 8083 9832
rect 5394 9824 5710 9825
rect 5394 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5710 9824
rect 5394 9759 5710 9760
rect 5812 9618 5872 9830
rect 8017 9827 8083 9830
rect 9842 9824 10158 9825
rect 9842 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10158 9824
rect 9842 9759 10158 9760
rect 14290 9824 14606 9825
rect 14290 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14606 9824
rect 14290 9759 14606 9760
rect 6269 9754 6335 9757
rect 9581 9754 9647 9757
rect 6269 9752 9647 9754
rect 6269 9696 6274 9752
rect 6330 9696 9586 9752
rect 9642 9696 9647 9752
rect 6269 9694 9647 9696
rect 6269 9691 6335 9694
rect 9581 9691 9647 9694
rect 12893 9756 12959 9757
rect 12893 9752 12940 9756
rect 13004 9754 13010 9756
rect 12893 9696 12898 9752
rect 12893 9692 12940 9696
rect 13004 9694 13050 9754
rect 13004 9692 13010 9694
rect 12893 9691 12959 9692
rect 5214 9558 5872 9618
rect 6729 9618 6795 9621
rect 7649 9618 7715 9621
rect 9213 9618 9279 9621
rect 18137 9618 18203 9621
rect 19200 9618 20000 9648
rect 6729 9616 18203 9618
rect 6729 9560 6734 9616
rect 6790 9560 7654 9616
rect 7710 9560 9218 9616
rect 9274 9560 18142 9616
rect 18198 9560 18203 9616
rect 6729 9558 18203 9560
rect 6729 9555 6795 9558
rect 7649 9555 7715 9558
rect 9213 9555 9279 9558
rect 18137 9555 18203 9558
rect 18278 9558 20000 9618
rect 3141 9482 3207 9485
rect 4981 9482 5047 9485
rect 10225 9482 10291 9485
rect 12065 9482 12131 9485
rect 3141 9480 10291 9482
rect 3141 9424 3146 9480
rect 3202 9424 4986 9480
rect 5042 9424 10230 9480
rect 10286 9424 10291 9480
rect 3141 9422 10291 9424
rect 3141 9419 3207 9422
rect 4981 9419 5047 9422
rect 10225 9419 10291 9422
rect 11838 9480 12131 9482
rect 11838 9424 12070 9480
rect 12126 9424 12131 9480
rect 11838 9422 12131 9424
rect 0 9346 800 9376
rect 2865 9346 2931 9349
rect 0 9344 2931 9346
rect 0 9288 2870 9344
rect 2926 9288 2931 9344
rect 0 9286 2931 9288
rect 0 9256 800 9286
rect 2865 9283 2931 9286
rect 8293 9346 8359 9349
rect 8293 9344 9276 9346
rect 8293 9288 8298 9344
rect 8354 9288 9276 9344
rect 8293 9286 9276 9288
rect 8293 9283 8359 9286
rect 3170 9280 3486 9281
rect 3170 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3486 9280
rect 3170 9215 3486 9216
rect 7618 9280 7934 9281
rect 7618 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7934 9280
rect 7618 9215 7934 9216
rect 9216 9213 9276 9286
rect 9438 9284 9444 9348
rect 9508 9346 9514 9348
rect 9581 9346 9647 9349
rect 9508 9344 9647 9346
rect 9508 9288 9586 9344
rect 9642 9288 9647 9344
rect 9508 9286 9647 9288
rect 9508 9284 9514 9286
rect 9581 9283 9647 9286
rect 9765 9346 9831 9349
rect 11838 9346 11898 9422
rect 12065 9419 12131 9422
rect 17217 9482 17283 9485
rect 18278 9482 18338 9558
rect 19200 9528 20000 9558
rect 17217 9480 18338 9482
rect 17217 9424 17222 9480
rect 17278 9424 18338 9480
rect 17217 9422 18338 9424
rect 17217 9419 17283 9422
rect 9765 9344 11898 9346
rect 9765 9288 9770 9344
rect 9826 9288 11898 9344
rect 9765 9286 11898 9288
rect 17033 9346 17099 9349
rect 17166 9346 17172 9348
rect 17033 9344 17172 9346
rect 17033 9288 17038 9344
rect 17094 9288 17172 9344
rect 17033 9286 17172 9288
rect 9765 9283 9831 9286
rect 17033 9283 17099 9286
rect 17166 9284 17172 9286
rect 17236 9284 17242 9348
rect 12066 9280 12382 9281
rect 12066 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12382 9280
rect 12066 9215 12382 9216
rect 16514 9280 16830 9281
rect 16514 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16830 9280
rect 16514 9215 16830 9216
rect 8937 9210 9003 9213
rect 8020 9208 9003 9210
rect 8020 9152 8942 9208
rect 8998 9152 9003 9208
rect 8020 9150 9003 9152
rect 5993 9074 6059 9077
rect 8020 9074 8080 9150
rect 8937 9147 9003 9150
rect 9213 9210 9279 9213
rect 10409 9210 10475 9213
rect 9213 9208 10475 9210
rect 9213 9152 9218 9208
rect 9274 9152 10414 9208
rect 10470 9152 10475 9208
rect 9213 9150 10475 9152
rect 9213 9147 9279 9150
rect 10409 9147 10475 9150
rect 17677 9210 17743 9213
rect 19200 9210 20000 9240
rect 17677 9208 20000 9210
rect 17677 9152 17682 9208
rect 17738 9152 20000 9208
rect 17677 9150 20000 9152
rect 17677 9147 17743 9150
rect 19200 9120 20000 9150
rect 5993 9072 8080 9074
rect 5993 9016 5998 9072
rect 6054 9016 8080 9072
rect 5993 9014 8080 9016
rect 9029 9074 9095 9077
rect 12433 9074 12499 9077
rect 9029 9072 12499 9074
rect 9029 9016 9034 9072
rect 9090 9016 12438 9072
rect 12494 9016 12499 9072
rect 9029 9014 12499 9016
rect 5993 9011 6059 9014
rect 9029 9011 9095 9014
rect 12433 9011 12499 9014
rect 13353 9074 13419 9077
rect 17861 9074 17927 9077
rect 13353 9072 17927 9074
rect 13353 9016 13358 9072
rect 13414 9016 17866 9072
rect 17922 9016 17927 9072
rect 13353 9014 17927 9016
rect 13353 9011 13419 9014
rect 17861 9011 17927 9014
rect 0 8938 800 8968
rect 3969 8938 4035 8941
rect 0 8936 4035 8938
rect 0 8880 3974 8936
rect 4030 8880 4035 8936
rect 0 8878 4035 8880
rect 0 8848 800 8878
rect 3969 8875 4035 8878
rect 4838 8876 4844 8940
rect 4908 8938 4914 8940
rect 5533 8938 5599 8941
rect 4908 8936 5599 8938
rect 4908 8880 5538 8936
rect 5594 8880 5599 8936
rect 4908 8878 5599 8880
rect 4908 8876 4914 8878
rect 5533 8875 5599 8878
rect 5809 8938 5875 8941
rect 16205 8938 16271 8941
rect 5809 8936 16271 8938
rect 5809 8880 5814 8936
rect 5870 8880 16210 8936
rect 16266 8880 16271 8936
rect 5809 8878 16271 8880
rect 5809 8875 5875 8878
rect 16205 8875 16271 8878
rect 2957 8804 3023 8805
rect 2957 8802 3004 8804
rect 2912 8800 3004 8802
rect 2912 8744 2962 8800
rect 2912 8742 3004 8744
rect 2957 8740 3004 8742
rect 3068 8740 3074 8804
rect 5073 8802 5139 8805
rect 5206 8802 5212 8804
rect 5073 8800 5212 8802
rect 5073 8744 5078 8800
rect 5134 8744 5212 8800
rect 5073 8742 5212 8744
rect 2957 8739 3023 8740
rect 5073 8739 5139 8742
rect 5206 8740 5212 8742
rect 5276 8740 5282 8804
rect 5901 8802 5967 8805
rect 9213 8802 9279 8805
rect 5901 8800 9279 8802
rect 5901 8744 5906 8800
rect 5962 8744 9218 8800
rect 9274 8744 9279 8800
rect 5901 8742 9279 8744
rect 5901 8739 5967 8742
rect 9213 8739 9279 8742
rect 10409 8802 10475 8805
rect 13537 8802 13603 8805
rect 10409 8800 13603 8802
rect 10409 8744 10414 8800
rect 10470 8744 13542 8800
rect 13598 8744 13603 8800
rect 10409 8742 13603 8744
rect 10409 8739 10475 8742
rect 13537 8739 13603 8742
rect 14825 8802 14891 8805
rect 17677 8802 17743 8805
rect 14825 8800 17743 8802
rect 14825 8744 14830 8800
rect 14886 8744 17682 8800
rect 17738 8744 17743 8800
rect 14825 8742 17743 8744
rect 14825 8739 14891 8742
rect 17677 8739 17743 8742
rect 17861 8802 17927 8805
rect 19200 8802 20000 8832
rect 17861 8800 20000 8802
rect 17861 8744 17866 8800
rect 17922 8744 20000 8800
rect 17861 8742 20000 8744
rect 17861 8739 17927 8742
rect 5394 8736 5710 8737
rect 5394 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5710 8736
rect 5394 8671 5710 8672
rect 9842 8736 10158 8737
rect 9842 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10158 8736
rect 9842 8671 10158 8672
rect 14290 8736 14606 8737
rect 14290 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14606 8736
rect 19200 8712 20000 8742
rect 14290 8671 14606 8672
rect 4981 8666 5047 8669
rect 6821 8666 6887 8669
rect 7281 8666 7347 8669
rect 4981 8664 5090 8666
rect 4981 8608 4986 8664
rect 5042 8608 5090 8664
rect 4981 8603 5090 8608
rect 6821 8664 7347 8666
rect 6821 8608 6826 8664
rect 6882 8608 7286 8664
rect 7342 8608 7347 8664
rect 6821 8606 7347 8608
rect 6821 8603 6887 8606
rect 7281 8603 7347 8606
rect 7557 8666 7623 8669
rect 8845 8666 8911 8669
rect 9581 8666 9647 8669
rect 7557 8664 9647 8666
rect 7557 8608 7562 8664
rect 7618 8608 8850 8664
rect 8906 8608 9586 8664
rect 9642 8608 9647 8664
rect 7557 8606 9647 8608
rect 7557 8603 7623 8606
rect 8845 8603 8911 8606
rect 9581 8603 9647 8606
rect 15929 8666 15995 8669
rect 17125 8666 17191 8669
rect 15929 8664 17191 8666
rect 15929 8608 15934 8664
rect 15990 8608 17130 8664
rect 17186 8608 17191 8664
rect 15929 8606 17191 8608
rect 15929 8603 15995 8606
rect 17125 8603 17191 8606
rect 0 8530 800 8560
rect 1669 8530 1735 8533
rect 0 8528 1735 8530
rect 0 8472 1674 8528
rect 1730 8472 1735 8528
rect 0 8470 1735 8472
rect 0 8440 800 8470
rect 1669 8467 1735 8470
rect 1945 8530 2011 8533
rect 5030 8530 5090 8603
rect 8753 8530 8819 8533
rect 9254 8530 9260 8532
rect 1945 8528 4308 8530
rect 1945 8472 1950 8528
rect 2006 8472 4308 8528
rect 1945 8470 4308 8472
rect 5030 8470 8402 8530
rect 1945 8467 2011 8470
rect 2630 8332 2636 8396
rect 2700 8394 2706 8396
rect 3417 8394 3483 8397
rect 2700 8392 3483 8394
rect 2700 8336 3422 8392
rect 3478 8336 3483 8392
rect 2700 8334 3483 8336
rect 4248 8394 4308 8470
rect 7557 8394 7623 8397
rect 4248 8392 7623 8394
rect 4248 8336 7562 8392
rect 7618 8336 7623 8392
rect 4248 8334 7623 8336
rect 2700 8332 2706 8334
rect 3417 8331 3483 8334
rect 7557 8331 7623 8334
rect 3601 8258 3667 8261
rect 4429 8258 4495 8261
rect 3601 8256 4495 8258
rect 3601 8200 3606 8256
rect 3662 8200 4434 8256
rect 4490 8200 4495 8256
rect 3601 8198 4495 8200
rect 8342 8258 8402 8470
rect 8753 8528 9260 8530
rect 8753 8472 8758 8528
rect 8814 8472 9260 8528
rect 8753 8470 9260 8472
rect 8753 8467 8819 8470
rect 9254 8468 9260 8470
rect 9324 8468 9330 8532
rect 9489 8530 9555 8533
rect 10685 8530 10751 8533
rect 9489 8528 10751 8530
rect 9489 8472 9494 8528
rect 9550 8472 10690 8528
rect 10746 8472 10751 8528
rect 9489 8470 10751 8472
rect 9489 8467 9555 8470
rect 10685 8467 10751 8470
rect 14774 8468 14780 8532
rect 14844 8530 14850 8532
rect 14844 8470 17234 8530
rect 14844 8468 14850 8470
rect 14917 8394 14983 8397
rect 17033 8394 17099 8397
rect 11838 8334 12634 8394
rect 11838 8258 11898 8334
rect 8342 8198 11898 8258
rect 12574 8258 12634 8334
rect 14917 8392 17099 8394
rect 14917 8336 14922 8392
rect 14978 8336 17038 8392
rect 17094 8336 17099 8392
rect 14917 8334 17099 8336
rect 17174 8394 17234 8470
rect 17585 8394 17651 8397
rect 17174 8392 17651 8394
rect 17174 8336 17590 8392
rect 17646 8336 17651 8392
rect 17174 8334 17651 8336
rect 14917 8331 14983 8334
rect 17033 8331 17099 8334
rect 17585 8331 17651 8334
rect 18045 8394 18111 8397
rect 19200 8394 20000 8424
rect 18045 8392 20000 8394
rect 18045 8336 18050 8392
rect 18106 8336 20000 8392
rect 18045 8334 20000 8336
rect 18045 8331 18111 8334
rect 19200 8304 20000 8334
rect 15929 8258 15995 8261
rect 12574 8256 15995 8258
rect 12574 8200 15934 8256
rect 15990 8200 15995 8256
rect 12574 8198 15995 8200
rect 3601 8195 3667 8198
rect 4429 8195 4495 8198
rect 15929 8195 15995 8198
rect 3170 8192 3486 8193
rect 0 8122 800 8152
rect 3170 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3486 8192
rect 3170 8127 3486 8128
rect 7618 8192 7934 8193
rect 7618 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7934 8192
rect 7618 8127 7934 8128
rect 12066 8192 12382 8193
rect 12066 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12382 8192
rect 12066 8127 12382 8128
rect 16514 8192 16830 8193
rect 16514 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16830 8192
rect 16514 8127 16830 8128
rect 2221 8122 2287 8125
rect 0 8120 2287 8122
rect 0 8064 2226 8120
rect 2282 8064 2287 8120
rect 0 8062 2287 8064
rect 0 8032 800 8062
rect 2221 8059 2287 8062
rect 3417 7986 3483 7989
rect 3734 7986 3740 7988
rect 3417 7984 3740 7986
rect 3417 7928 3422 7984
rect 3478 7928 3740 7984
rect 3417 7926 3740 7928
rect 3417 7923 3483 7926
rect 3734 7924 3740 7926
rect 3804 7924 3810 7988
rect 5625 7986 5691 7989
rect 15469 7986 15535 7989
rect 15745 7986 15811 7989
rect 5625 7984 12818 7986
rect 5625 7928 5630 7984
rect 5686 7928 12818 7984
rect 5625 7926 12818 7928
rect 5625 7923 5691 7926
rect 1669 7850 1735 7853
rect 12758 7850 12818 7926
rect 15469 7984 15811 7986
rect 15469 7928 15474 7984
rect 15530 7928 15750 7984
rect 15806 7928 15811 7984
rect 15469 7926 15811 7928
rect 15469 7923 15535 7926
rect 15745 7923 15811 7926
rect 15929 7986 15995 7989
rect 17861 7986 17927 7989
rect 15929 7984 17927 7986
rect 15929 7928 15934 7984
rect 15990 7928 17866 7984
rect 17922 7928 17927 7984
rect 15929 7926 17927 7928
rect 15929 7923 15995 7926
rect 17861 7923 17927 7926
rect 18045 7986 18111 7989
rect 19200 7986 20000 8016
rect 18045 7984 20000 7986
rect 18045 7928 18050 7984
rect 18106 7928 20000 7984
rect 18045 7926 20000 7928
rect 18045 7923 18111 7926
rect 19200 7896 20000 7926
rect 12893 7850 12959 7853
rect 16849 7850 16915 7853
rect 1669 7848 12634 7850
rect 1669 7792 1674 7848
rect 1730 7792 12634 7848
rect 1669 7790 12634 7792
rect 12758 7848 16915 7850
rect 12758 7792 12898 7848
rect 12954 7792 16854 7848
rect 16910 7792 16915 7848
rect 12758 7790 16915 7792
rect 1669 7787 1735 7790
rect 0 7714 800 7744
rect 1485 7714 1551 7717
rect 0 7712 1551 7714
rect 0 7656 1490 7712
rect 1546 7656 1551 7712
rect 0 7654 1551 7656
rect 0 7624 800 7654
rect 1485 7651 1551 7654
rect 2221 7714 2287 7717
rect 4245 7714 4311 7717
rect 2221 7712 4311 7714
rect 2221 7656 2226 7712
rect 2282 7656 4250 7712
rect 4306 7656 4311 7712
rect 2221 7654 4311 7656
rect 12574 7714 12634 7790
rect 12893 7787 12959 7790
rect 16849 7787 16915 7790
rect 13261 7714 13327 7717
rect 12574 7712 13327 7714
rect 12574 7656 13266 7712
rect 13322 7656 13327 7712
rect 12574 7654 13327 7656
rect 2221 7651 2287 7654
rect 4245 7651 4311 7654
rect 13261 7651 13327 7654
rect 5394 7648 5710 7649
rect 5394 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5710 7648
rect 5394 7583 5710 7584
rect 9842 7648 10158 7649
rect 9842 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10158 7648
rect 9842 7583 10158 7584
rect 14290 7648 14606 7649
rect 14290 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14606 7648
rect 14290 7583 14606 7584
rect 2589 7578 2655 7581
rect 3785 7578 3851 7581
rect 2589 7576 3851 7578
rect 2589 7520 2594 7576
rect 2650 7520 3790 7576
rect 3846 7520 3851 7576
rect 2589 7518 3851 7520
rect 2589 7515 2655 7518
rect 3785 7515 3851 7518
rect 4286 7516 4292 7580
rect 4356 7578 4362 7580
rect 4521 7578 4587 7581
rect 4654 7578 4660 7580
rect 4356 7576 4660 7578
rect 4356 7520 4526 7576
rect 4582 7520 4660 7576
rect 4356 7518 4660 7520
rect 4356 7516 4362 7518
rect 4521 7515 4587 7518
rect 4654 7516 4660 7518
rect 4724 7516 4730 7580
rect 18413 7578 18479 7581
rect 19200 7578 20000 7608
rect 18413 7576 20000 7578
rect 18413 7520 18418 7576
rect 18474 7520 20000 7576
rect 18413 7518 20000 7520
rect 18413 7515 18479 7518
rect 19200 7488 20000 7518
rect 2221 7442 2287 7445
rect 3417 7442 3483 7445
rect 5165 7442 5231 7445
rect 2221 7440 2790 7442
rect 2221 7384 2226 7440
rect 2282 7384 2790 7440
rect 2221 7382 2790 7384
rect 2221 7379 2287 7382
rect 0 7306 800 7336
rect 1485 7306 1551 7309
rect 0 7304 1551 7306
rect 0 7248 1490 7304
rect 1546 7248 1551 7304
rect 0 7246 1551 7248
rect 2730 7306 2790 7382
rect 3417 7440 5231 7442
rect 3417 7384 3422 7440
rect 3478 7384 5170 7440
rect 5226 7384 5231 7440
rect 3417 7382 5231 7384
rect 3417 7379 3483 7382
rect 5165 7379 5231 7382
rect 5625 7442 5691 7445
rect 5942 7442 5948 7444
rect 5625 7440 5948 7442
rect 5625 7384 5630 7440
rect 5686 7384 5948 7440
rect 5625 7382 5948 7384
rect 5625 7379 5691 7382
rect 5942 7380 5948 7382
rect 6012 7380 6018 7444
rect 11605 7442 11671 7445
rect 15653 7442 15719 7445
rect 11605 7440 15719 7442
rect 11605 7384 11610 7440
rect 11666 7384 15658 7440
rect 15714 7384 15719 7440
rect 11605 7382 15719 7384
rect 11605 7379 11671 7382
rect 15653 7379 15719 7382
rect 3325 7306 3391 7309
rect 16297 7306 16363 7309
rect 17493 7306 17559 7309
rect 2730 7304 17559 7306
rect 2730 7248 3330 7304
rect 3386 7248 16302 7304
rect 16358 7248 17498 7304
rect 17554 7248 17559 7304
rect 2730 7246 17559 7248
rect 0 7216 800 7246
rect 1485 7243 1551 7246
rect 3325 7243 3391 7246
rect 16297 7243 16363 7246
rect 17493 7243 17559 7246
rect 2589 7170 2655 7173
rect 2589 7168 3020 7170
rect 2589 7112 2594 7168
rect 2650 7112 3020 7168
rect 2589 7110 3020 7112
rect 2589 7107 2655 7110
rect 2960 7037 3020 7110
rect 4838 7108 4844 7172
rect 4908 7170 4914 7172
rect 5625 7170 5691 7173
rect 6913 7170 6979 7173
rect 4908 7168 6979 7170
rect 4908 7112 5630 7168
rect 5686 7112 6918 7168
rect 6974 7112 6979 7168
rect 4908 7110 6979 7112
rect 4908 7108 4914 7110
rect 5625 7107 5691 7110
rect 6913 7107 6979 7110
rect 18045 7170 18111 7173
rect 19200 7170 20000 7200
rect 18045 7168 20000 7170
rect 18045 7112 18050 7168
rect 18106 7112 20000 7168
rect 18045 7110 20000 7112
rect 18045 7107 18111 7110
rect 3170 7104 3486 7105
rect 3170 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3486 7104
rect 3170 7039 3486 7040
rect 7618 7104 7934 7105
rect 7618 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7934 7104
rect 7618 7039 7934 7040
rect 12066 7104 12382 7105
rect 12066 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12382 7104
rect 12066 7039 12382 7040
rect 16514 7104 16830 7105
rect 16514 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16830 7104
rect 19200 7080 20000 7110
rect 16514 7039 16830 7040
rect 2446 6972 2452 7036
rect 2516 7034 2522 7036
rect 2589 7034 2655 7037
rect 2516 7032 2655 7034
rect 2516 6976 2594 7032
rect 2650 6976 2655 7032
rect 2516 6974 2655 6976
rect 2516 6972 2522 6974
rect 2589 6971 2655 6974
rect 2957 7032 3023 7037
rect 2957 6976 2962 7032
rect 3018 6976 3023 7032
rect 2957 6971 3023 6976
rect 5206 6972 5212 7036
rect 5276 7034 5282 7036
rect 5533 7034 5599 7037
rect 15653 7034 15719 7037
rect 5276 7032 7482 7034
rect 5276 6976 5538 7032
rect 5594 6976 7482 7032
rect 5276 6974 7482 6976
rect 5276 6972 5282 6974
rect 5533 6971 5599 6974
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 4061 6900 4127 6901
rect 4061 6898 4108 6900
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 2730 6896 4108 6898
rect 2730 6840 4066 6896
rect 2730 6838 4108 6840
rect 2589 6762 2655 6765
rect 2730 6762 2790 6838
rect 4061 6836 4108 6838
rect 4172 6836 4178 6900
rect 4613 6898 4679 6901
rect 4797 6898 4863 6901
rect 4613 6896 4863 6898
rect 4613 6840 4618 6896
rect 4674 6840 4802 6896
rect 4858 6840 4863 6896
rect 4613 6838 4863 6840
rect 7422 6898 7482 6974
rect 8020 6974 11898 7034
rect 8020 6898 8080 6974
rect 7422 6838 8080 6898
rect 11838 6898 11898 6974
rect 12574 7032 15719 7034
rect 12574 6976 15658 7032
rect 15714 6976 15719 7032
rect 12574 6974 15719 6976
rect 12574 6898 12634 6974
rect 15653 6971 15719 6974
rect 11838 6838 12634 6898
rect 4061 6835 4127 6836
rect 4613 6835 4679 6838
rect 4797 6835 4863 6838
rect 2589 6760 2790 6762
rect 2589 6704 2594 6760
rect 2650 6704 2790 6760
rect 2589 6702 2790 6704
rect 2589 6699 2655 6702
rect 2998 6700 3004 6764
rect 3068 6762 3074 6764
rect 4337 6762 4403 6765
rect 8937 6762 9003 6765
rect 3068 6760 9003 6762
rect 3068 6704 4342 6760
rect 4398 6704 8942 6760
rect 8998 6704 9003 6760
rect 3068 6702 9003 6704
rect 3068 6700 3074 6702
rect 2037 6626 2103 6629
rect 3006 6626 3066 6700
rect 4337 6699 4403 6702
rect 8937 6699 9003 6702
rect 13261 6762 13327 6765
rect 16481 6762 16547 6765
rect 17217 6762 17283 6765
rect 13261 6760 17283 6762
rect 13261 6704 13266 6760
rect 13322 6704 16486 6760
rect 16542 6704 17222 6760
rect 17278 6704 17283 6760
rect 13261 6702 17283 6704
rect 13261 6699 13327 6702
rect 16481 6699 16547 6702
rect 17217 6699 17283 6702
rect 18413 6762 18479 6765
rect 19200 6762 20000 6792
rect 18413 6760 20000 6762
rect 18413 6704 18418 6760
rect 18474 6704 20000 6760
rect 18413 6702 20000 6704
rect 18413 6699 18479 6702
rect 19200 6672 20000 6702
rect 2037 6624 3066 6626
rect 2037 6568 2042 6624
rect 2098 6568 3066 6624
rect 2037 6566 3066 6568
rect 2037 6563 2103 6566
rect 5394 6560 5710 6561
rect 0 6490 800 6520
rect 5394 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5710 6560
rect 5394 6495 5710 6496
rect 9842 6560 10158 6561
rect 9842 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10158 6560
rect 9842 6495 10158 6496
rect 14290 6560 14606 6561
rect 14290 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14606 6560
rect 14290 6495 14606 6496
rect 1577 6490 1643 6493
rect 0 6488 1643 6490
rect 0 6432 1582 6488
rect 1638 6432 1643 6488
rect 0 6430 1643 6432
rect 0 6400 800 6430
rect 1577 6427 1643 6430
rect 2405 6490 2471 6493
rect 5206 6490 5212 6492
rect 2405 6488 5212 6490
rect 2405 6432 2410 6488
rect 2466 6432 5212 6488
rect 2405 6430 5212 6432
rect 2405 6427 2471 6430
rect 5206 6428 5212 6430
rect 5276 6428 5282 6492
rect 17718 6428 17724 6492
rect 17788 6490 17794 6492
rect 18045 6490 18111 6493
rect 17788 6488 18111 6490
rect 17788 6432 18050 6488
rect 18106 6432 18111 6488
rect 17788 6430 18111 6432
rect 17788 6428 17794 6430
rect 18045 6427 18111 6430
rect 2681 6354 2747 6357
rect 6821 6354 6887 6357
rect 2681 6352 6887 6354
rect 2681 6296 2686 6352
rect 2742 6296 6826 6352
rect 6882 6296 6887 6352
rect 2681 6294 6887 6296
rect 2681 6291 2747 6294
rect 6821 6291 6887 6294
rect 18505 6354 18571 6357
rect 19200 6354 20000 6384
rect 18505 6352 20000 6354
rect 18505 6296 18510 6352
rect 18566 6296 20000 6352
rect 18505 6294 20000 6296
rect 18505 6291 18571 6294
rect 19200 6264 20000 6294
rect 1393 6218 1459 6221
rect 1166 6216 1459 6218
rect 1166 6160 1398 6216
rect 1454 6160 1459 6216
rect 1166 6158 1459 6160
rect 0 6082 800 6112
rect 1166 6082 1226 6158
rect 1393 6155 1459 6158
rect 3417 6218 3483 6221
rect 3785 6218 3851 6221
rect 10409 6218 10475 6221
rect 3417 6216 10475 6218
rect 3417 6160 3422 6216
rect 3478 6160 3790 6216
rect 3846 6160 10414 6216
rect 10470 6160 10475 6216
rect 3417 6158 10475 6160
rect 3417 6155 3483 6158
rect 3785 6155 3851 6158
rect 10409 6155 10475 6158
rect 0 6022 1226 6082
rect 0 5992 800 6022
rect 3170 6016 3486 6017
rect 3170 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3486 6016
rect 3170 5951 3486 5952
rect 7618 6016 7934 6017
rect 7618 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7934 6016
rect 7618 5951 7934 5952
rect 12066 6016 12382 6017
rect 12066 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12382 6016
rect 12066 5951 12382 5952
rect 16514 6016 16830 6017
rect 16514 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16830 6016
rect 16514 5951 16830 5952
rect 18597 5946 18663 5949
rect 19200 5946 20000 5976
rect 18597 5944 20000 5946
rect 18597 5888 18602 5944
rect 18658 5888 20000 5944
rect 18597 5886 20000 5888
rect 18597 5883 18663 5886
rect 19200 5856 20000 5886
rect 0 5674 800 5704
rect 1761 5674 1827 5677
rect 0 5672 1827 5674
rect 0 5616 1766 5672
rect 1822 5616 1827 5672
rect 0 5614 1827 5616
rect 0 5584 800 5614
rect 1761 5611 1827 5614
rect 4429 5674 4495 5677
rect 6085 5674 6151 5677
rect 4429 5672 6151 5674
rect 4429 5616 4434 5672
rect 4490 5616 6090 5672
rect 6146 5616 6151 5672
rect 4429 5614 6151 5616
rect 4429 5611 4495 5614
rect 6085 5611 6151 5614
rect 15193 5674 15259 5677
rect 16205 5674 16271 5677
rect 17493 5674 17559 5677
rect 15193 5672 17559 5674
rect 15193 5616 15198 5672
rect 15254 5616 16210 5672
rect 16266 5616 17498 5672
rect 17554 5616 17559 5672
rect 15193 5614 17559 5616
rect 15193 5611 15259 5614
rect 16205 5611 16271 5614
rect 17493 5611 17559 5614
rect 17953 5538 18019 5541
rect 19200 5538 20000 5568
rect 17953 5536 20000 5538
rect 17953 5480 17958 5536
rect 18014 5480 20000 5536
rect 17953 5478 20000 5480
rect 17953 5475 18019 5478
rect 5394 5472 5710 5473
rect 5394 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5710 5472
rect 5394 5407 5710 5408
rect 9842 5472 10158 5473
rect 9842 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10158 5472
rect 9842 5407 10158 5408
rect 14290 5472 14606 5473
rect 14290 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14606 5472
rect 19200 5448 20000 5478
rect 14290 5407 14606 5408
rect 7414 5340 7420 5404
rect 7484 5402 7490 5404
rect 9673 5402 9739 5405
rect 7484 5400 9739 5402
rect 7484 5344 9678 5400
rect 9734 5344 9739 5400
rect 7484 5342 9739 5344
rect 7484 5340 7490 5342
rect 9673 5339 9739 5342
rect 0 5266 800 5296
rect 933 5266 999 5269
rect 0 5264 999 5266
rect 0 5208 938 5264
rect 994 5208 999 5264
rect 0 5206 999 5208
rect 0 5176 800 5206
rect 933 5203 999 5206
rect 18689 5130 18755 5133
rect 19200 5130 20000 5160
rect 18689 5128 20000 5130
rect 18689 5072 18694 5128
rect 18750 5072 20000 5128
rect 18689 5070 20000 5072
rect 18689 5067 18755 5070
rect 19200 5040 20000 5070
rect 3170 4928 3486 4929
rect 0 4858 800 4888
rect 3170 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3486 4928
rect 3170 4863 3486 4864
rect 7618 4928 7934 4929
rect 7618 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7934 4928
rect 7618 4863 7934 4864
rect 12066 4928 12382 4929
rect 12066 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12382 4928
rect 12066 4863 12382 4864
rect 16514 4928 16830 4929
rect 16514 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16830 4928
rect 16514 4863 16830 4864
rect 2957 4858 3023 4861
rect 0 4856 3023 4858
rect 0 4800 2962 4856
rect 3018 4800 3023 4856
rect 0 4798 3023 4800
rect 0 4768 800 4798
rect 2957 4795 3023 4798
rect 2129 4722 2195 4725
rect 2630 4722 2636 4724
rect 2129 4720 2636 4722
rect 2129 4664 2134 4720
rect 2190 4664 2636 4720
rect 2129 4662 2636 4664
rect 2129 4659 2195 4662
rect 2630 4660 2636 4662
rect 2700 4722 2706 4724
rect 11237 4722 11303 4725
rect 2700 4720 11303 4722
rect 2700 4664 11242 4720
rect 11298 4664 11303 4720
rect 2700 4662 11303 4664
rect 2700 4660 2706 4662
rect 11237 4659 11303 4662
rect 18137 4722 18203 4725
rect 19200 4722 20000 4752
rect 18137 4720 20000 4722
rect 18137 4664 18142 4720
rect 18198 4664 20000 4720
rect 18137 4662 20000 4664
rect 18137 4659 18203 4662
rect 19200 4632 20000 4662
rect 0 4450 800 4480
rect 2221 4450 2287 4453
rect 0 4448 2287 4450
rect 0 4392 2226 4448
rect 2282 4392 2287 4448
rect 0 4390 2287 4392
rect 0 4360 800 4390
rect 2221 4387 2287 4390
rect 5394 4384 5710 4385
rect 5394 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5710 4384
rect 5394 4319 5710 4320
rect 9842 4384 10158 4385
rect 9842 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10158 4384
rect 9842 4319 10158 4320
rect 14290 4384 14606 4385
rect 14290 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14606 4384
rect 14290 4319 14606 4320
rect 18873 4314 18939 4317
rect 19200 4314 20000 4344
rect 18873 4312 20000 4314
rect 18873 4256 18878 4312
rect 18934 4256 20000 4312
rect 18873 4254 20000 4256
rect 18873 4251 18939 4254
rect 19200 4224 20000 4254
rect 2773 4180 2839 4181
rect 2773 4176 2820 4180
rect 2884 4178 2890 4180
rect 2773 4120 2778 4176
rect 2773 4116 2820 4120
rect 2884 4118 2930 4178
rect 2884 4116 2890 4118
rect 2773 4115 2839 4116
rect 0 4042 800 4072
rect 1669 4042 1735 4045
rect 0 4040 1735 4042
rect 0 3984 1674 4040
rect 1730 3984 1735 4040
rect 0 3982 1735 3984
rect 0 3952 800 3982
rect 1669 3979 1735 3982
rect 4153 4042 4219 4045
rect 6453 4042 6519 4045
rect 4153 4040 6519 4042
rect 4153 3984 4158 4040
rect 4214 3984 6458 4040
rect 6514 3984 6519 4040
rect 4153 3982 6519 3984
rect 4153 3979 4219 3982
rect 6453 3979 6519 3982
rect 9305 4042 9371 4045
rect 11513 4042 11579 4045
rect 9305 4040 11579 4042
rect 9305 3984 9310 4040
rect 9366 3984 11518 4040
rect 11574 3984 11579 4040
rect 9305 3982 11579 3984
rect 9305 3979 9371 3982
rect 11513 3979 11579 3982
rect 15285 4042 15351 4045
rect 16246 4042 16252 4044
rect 15285 4040 16252 4042
rect 15285 3984 15290 4040
rect 15346 3984 16252 4040
rect 15285 3982 16252 3984
rect 15285 3979 15351 3982
rect 16246 3980 16252 3982
rect 16316 3980 16322 4044
rect 17166 3980 17172 4044
rect 17236 4042 17242 4044
rect 17401 4042 17467 4045
rect 17236 4040 17467 4042
rect 17236 3984 17406 4040
rect 17462 3984 17467 4040
rect 17236 3982 17467 3984
rect 17236 3980 17242 3982
rect 17401 3979 17467 3982
rect 14958 3844 14964 3908
rect 15028 3906 15034 3908
rect 16113 3906 16179 3909
rect 15028 3904 16179 3906
rect 15028 3848 16118 3904
rect 16174 3848 16179 3904
rect 15028 3846 16179 3848
rect 15028 3844 15034 3846
rect 16113 3843 16179 3846
rect 18965 3906 19031 3909
rect 19200 3906 20000 3936
rect 18965 3904 20000 3906
rect 18965 3848 18970 3904
rect 19026 3848 20000 3904
rect 18965 3846 20000 3848
rect 18965 3843 19031 3846
rect 3170 3840 3486 3841
rect 3170 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3486 3840
rect 3170 3775 3486 3776
rect 7618 3840 7934 3841
rect 7618 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7934 3840
rect 7618 3775 7934 3776
rect 12066 3840 12382 3841
rect 12066 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12382 3840
rect 12066 3775 12382 3776
rect 16514 3840 16830 3841
rect 16514 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16830 3840
rect 19200 3816 20000 3846
rect 16514 3775 16830 3776
rect 0 3634 800 3664
rect 1853 3634 1919 3637
rect 0 3632 1919 3634
rect 0 3576 1858 3632
rect 1914 3576 1919 3632
rect 0 3574 1919 3576
rect 0 3544 800 3574
rect 1853 3571 1919 3574
rect 8150 3572 8156 3636
rect 8220 3634 8226 3636
rect 8477 3634 8543 3637
rect 8220 3632 8543 3634
rect 8220 3576 8482 3632
rect 8538 3576 8543 3632
rect 8220 3574 8543 3576
rect 8220 3572 8226 3574
rect 8477 3571 8543 3574
rect 15142 3572 15148 3636
rect 15212 3634 15218 3636
rect 16941 3634 17007 3637
rect 15212 3632 17007 3634
rect 15212 3576 16946 3632
rect 17002 3576 17007 3632
rect 15212 3574 17007 3576
rect 15212 3572 15218 3574
rect 16941 3571 17007 3574
rect 3601 3498 3667 3501
rect 6269 3498 6335 3501
rect 3601 3496 6335 3498
rect 3601 3440 3606 3496
rect 3662 3440 6274 3496
rect 6330 3440 6335 3496
rect 3601 3438 6335 3440
rect 3601 3435 3667 3438
rect 6269 3435 6335 3438
rect 18229 3498 18295 3501
rect 19200 3498 20000 3528
rect 18229 3496 20000 3498
rect 18229 3440 18234 3496
rect 18290 3440 20000 3496
rect 18229 3438 20000 3440
rect 18229 3435 18295 3438
rect 19200 3408 20000 3438
rect 5394 3296 5710 3297
rect 0 3226 800 3256
rect 5394 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5710 3296
rect 5394 3231 5710 3232
rect 9842 3296 10158 3297
rect 9842 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10158 3296
rect 9842 3231 10158 3232
rect 14290 3296 14606 3297
rect 14290 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14606 3296
rect 14290 3231 14606 3232
rect 1485 3226 1551 3229
rect 0 3224 1551 3226
rect 0 3168 1490 3224
rect 1546 3168 1551 3224
rect 0 3166 1551 3168
rect 0 3136 800 3166
rect 1485 3163 1551 3166
rect 9438 3164 9444 3228
rect 9508 3226 9514 3228
rect 9581 3226 9647 3229
rect 9508 3224 9647 3226
rect 9508 3168 9586 3224
rect 9642 3168 9647 3224
rect 9508 3166 9647 3168
rect 9508 3164 9514 3166
rect 9581 3163 9647 3166
rect 3325 3090 3391 3093
rect 3550 3090 3556 3092
rect 3325 3088 3556 3090
rect 3325 3032 3330 3088
rect 3386 3032 3556 3088
rect 3325 3030 3556 3032
rect 3325 3027 3391 3030
rect 3550 3028 3556 3030
rect 3620 3028 3626 3092
rect 6085 3090 6151 3093
rect 6545 3090 6611 3093
rect 14457 3090 14523 3093
rect 6085 3088 14523 3090
rect 6085 3032 6090 3088
rect 6146 3032 6550 3088
rect 6606 3032 14462 3088
rect 14518 3032 14523 3088
rect 6085 3030 14523 3032
rect 6085 3027 6151 3030
rect 6545 3027 6611 3030
rect 14457 3027 14523 3030
rect 18045 3090 18111 3093
rect 19200 3090 20000 3120
rect 18045 3088 20000 3090
rect 18045 3032 18050 3088
rect 18106 3032 20000 3088
rect 18045 3030 20000 3032
rect 18045 3027 18111 3030
rect 19200 3000 20000 3030
rect 14365 2954 14431 2957
rect 17861 2954 17927 2957
rect 14365 2952 17927 2954
rect 14365 2896 14370 2952
rect 14426 2896 17866 2952
rect 17922 2896 17927 2952
rect 14365 2894 17927 2896
rect 14365 2891 14431 2894
rect 17861 2891 17927 2894
rect 0 2818 800 2848
rect 1945 2818 2011 2821
rect 0 2816 2011 2818
rect 0 2760 1950 2816
rect 2006 2760 2011 2816
rect 0 2758 2011 2760
rect 0 2728 800 2758
rect 1945 2755 2011 2758
rect 3170 2752 3486 2753
rect 3170 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3486 2752
rect 3170 2687 3486 2688
rect 7618 2752 7934 2753
rect 7618 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7934 2752
rect 7618 2687 7934 2688
rect 12066 2752 12382 2753
rect 12066 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12382 2752
rect 12066 2687 12382 2688
rect 16514 2752 16830 2753
rect 16514 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16830 2752
rect 16514 2687 16830 2688
rect 6453 2684 6519 2685
rect 6453 2680 6500 2684
rect 6564 2682 6570 2684
rect 18781 2682 18847 2685
rect 19200 2682 20000 2712
rect 6453 2624 6458 2680
rect 6453 2620 6500 2624
rect 6564 2622 6610 2682
rect 18781 2680 20000 2682
rect 18781 2624 18786 2680
rect 18842 2624 20000 2680
rect 18781 2622 20000 2624
rect 6564 2620 6570 2622
rect 6453 2619 6519 2620
rect 18781 2619 18847 2622
rect 19200 2592 20000 2622
rect 2497 2546 2563 2549
rect 4286 2546 4292 2548
rect 2497 2544 4292 2546
rect 2497 2488 2502 2544
rect 2558 2488 4292 2544
rect 2497 2486 4292 2488
rect 2497 2483 2563 2486
rect 4286 2484 4292 2486
rect 4356 2484 4362 2548
rect 12341 2546 12407 2549
rect 12934 2546 12940 2548
rect 12341 2544 12940 2546
rect 12341 2488 12346 2544
rect 12402 2488 12940 2544
rect 12341 2486 12940 2488
rect 12341 2483 12407 2486
rect 12934 2484 12940 2486
rect 13004 2484 13010 2548
rect 0 2410 800 2440
rect 1669 2410 1735 2413
rect 0 2408 1735 2410
rect 0 2352 1674 2408
rect 1730 2352 1735 2408
rect 0 2350 1735 2352
rect 0 2320 800 2350
rect 1669 2347 1735 2350
rect 4797 2410 4863 2413
rect 7925 2410 7991 2413
rect 4797 2408 7991 2410
rect 4797 2352 4802 2408
rect 4858 2352 7930 2408
rect 7986 2352 7991 2408
rect 4797 2350 7991 2352
rect 4797 2347 4863 2350
rect 7925 2347 7991 2350
rect 9254 2348 9260 2412
rect 9324 2410 9330 2412
rect 9673 2410 9739 2413
rect 9324 2408 9739 2410
rect 9324 2352 9678 2408
rect 9734 2352 9739 2408
rect 9324 2350 9739 2352
rect 9324 2348 9330 2350
rect 9673 2347 9739 2350
rect 18413 2274 18479 2277
rect 19200 2274 20000 2304
rect 18413 2272 20000 2274
rect 18413 2216 18418 2272
rect 18474 2216 20000 2272
rect 18413 2214 20000 2216
rect 18413 2211 18479 2214
rect 5394 2208 5710 2209
rect 5394 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5710 2208
rect 5394 2143 5710 2144
rect 9842 2208 10158 2209
rect 9842 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10158 2208
rect 9842 2143 10158 2144
rect 14290 2208 14606 2209
rect 14290 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14606 2208
rect 19200 2184 20000 2214
rect 14290 2143 14606 2144
rect 0 2002 800 2032
rect 1761 2002 1827 2005
rect 0 2000 1827 2002
rect 0 1944 1766 2000
rect 1822 1944 1827 2000
rect 0 1942 1827 1944
rect 0 1912 800 1942
rect 1761 1939 1827 1942
rect 17677 1866 17743 1869
rect 19200 1866 20000 1896
rect 17677 1864 20000 1866
rect 17677 1808 17682 1864
rect 17738 1808 20000 1864
rect 17677 1806 20000 1808
rect 17677 1803 17743 1806
rect 19200 1776 20000 1806
rect 0 1594 800 1624
rect 1485 1594 1551 1597
rect 0 1592 1551 1594
rect 0 1536 1490 1592
rect 1546 1536 1551 1592
rect 0 1534 1551 1536
rect 0 1504 800 1534
rect 1485 1531 1551 1534
rect 17309 1458 17375 1461
rect 19200 1458 20000 1488
rect 17309 1456 20000 1458
rect 17309 1400 17314 1456
rect 17370 1400 20000 1456
rect 17309 1398 20000 1400
rect 17309 1395 17375 1398
rect 19200 1368 20000 1398
rect 0 1186 800 1216
rect 1393 1186 1459 1189
rect 0 1184 1459 1186
rect 0 1128 1398 1184
rect 1454 1128 1459 1184
rect 0 1126 1459 1128
rect 0 1096 800 1126
rect 1393 1123 1459 1126
rect 17401 1050 17467 1053
rect 19200 1050 20000 1080
rect 17401 1048 20000 1050
rect 17401 992 17406 1048
rect 17462 992 20000 1048
rect 17401 990 20000 992
rect 17401 987 17467 990
rect 19200 960 20000 990
rect 0 778 800 808
rect 4061 778 4127 781
rect 0 776 4127 778
rect 0 720 4066 776
rect 4122 720 4127 776
rect 0 718 4127 720
rect 0 688 800 718
rect 4061 715 4127 718
rect 16297 642 16363 645
rect 19200 642 20000 672
rect 16297 640 20000 642
rect 16297 584 16302 640
rect 16358 584 20000 640
rect 16297 582 20000 584
rect 16297 579 16363 582
rect 19200 552 20000 582
rect 0 370 800 400
rect 2773 370 2839 373
rect 0 368 2839 370
rect 0 312 2778 368
rect 2834 312 2839 368
rect 0 310 2839 312
rect 0 280 800 310
rect 2773 307 2839 310
<< via3 >>
rect 17724 16084 17788 16148
rect 17724 15404 17788 15468
rect 3740 14996 3804 15060
rect 3176 14716 3240 14720
rect 3176 14660 3180 14716
rect 3180 14660 3236 14716
rect 3236 14660 3240 14716
rect 3176 14656 3240 14660
rect 3256 14716 3320 14720
rect 3256 14660 3260 14716
rect 3260 14660 3316 14716
rect 3316 14660 3320 14716
rect 3256 14656 3320 14660
rect 3336 14716 3400 14720
rect 3336 14660 3340 14716
rect 3340 14660 3396 14716
rect 3396 14660 3400 14716
rect 3336 14656 3400 14660
rect 3416 14716 3480 14720
rect 3416 14660 3420 14716
rect 3420 14660 3476 14716
rect 3476 14660 3480 14716
rect 3416 14656 3480 14660
rect 7624 14716 7688 14720
rect 7624 14660 7628 14716
rect 7628 14660 7684 14716
rect 7684 14660 7688 14716
rect 7624 14656 7688 14660
rect 7704 14716 7768 14720
rect 7704 14660 7708 14716
rect 7708 14660 7764 14716
rect 7764 14660 7768 14716
rect 7704 14656 7768 14660
rect 7784 14716 7848 14720
rect 7784 14660 7788 14716
rect 7788 14660 7844 14716
rect 7844 14660 7848 14716
rect 7784 14656 7848 14660
rect 7864 14716 7928 14720
rect 7864 14660 7868 14716
rect 7868 14660 7924 14716
rect 7924 14660 7928 14716
rect 7864 14656 7928 14660
rect 12072 14716 12136 14720
rect 12072 14660 12076 14716
rect 12076 14660 12132 14716
rect 12132 14660 12136 14716
rect 12072 14656 12136 14660
rect 12152 14716 12216 14720
rect 12152 14660 12156 14716
rect 12156 14660 12212 14716
rect 12212 14660 12216 14716
rect 12152 14656 12216 14660
rect 12232 14716 12296 14720
rect 12232 14660 12236 14716
rect 12236 14660 12292 14716
rect 12292 14660 12296 14716
rect 12232 14656 12296 14660
rect 12312 14716 12376 14720
rect 12312 14660 12316 14716
rect 12316 14660 12372 14716
rect 12372 14660 12376 14716
rect 12312 14656 12376 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 16760 14716 16824 14720
rect 16760 14660 16764 14716
rect 16764 14660 16820 14716
rect 16820 14660 16824 14716
rect 16760 14656 16824 14660
rect 5400 14172 5464 14176
rect 5400 14116 5404 14172
rect 5404 14116 5460 14172
rect 5460 14116 5464 14172
rect 5400 14112 5464 14116
rect 5480 14172 5544 14176
rect 5480 14116 5484 14172
rect 5484 14116 5540 14172
rect 5540 14116 5544 14172
rect 5480 14112 5544 14116
rect 5560 14172 5624 14176
rect 5560 14116 5564 14172
rect 5564 14116 5620 14172
rect 5620 14116 5624 14172
rect 5560 14112 5624 14116
rect 5640 14172 5704 14176
rect 5640 14116 5644 14172
rect 5644 14116 5700 14172
rect 5700 14116 5704 14172
rect 5640 14112 5704 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 14536 14172 14600 14176
rect 14536 14116 14540 14172
rect 14540 14116 14596 14172
rect 14596 14116 14600 14172
rect 14536 14112 14600 14116
rect 4660 13908 4724 13972
rect 14964 13772 15028 13836
rect 16252 13832 16316 13836
rect 16252 13776 16302 13832
rect 16302 13776 16316 13832
rect 16252 13772 16316 13776
rect 3176 13628 3240 13632
rect 3176 13572 3180 13628
rect 3180 13572 3236 13628
rect 3236 13572 3240 13628
rect 3176 13568 3240 13572
rect 3256 13628 3320 13632
rect 3256 13572 3260 13628
rect 3260 13572 3316 13628
rect 3316 13572 3320 13628
rect 3256 13568 3320 13572
rect 3336 13628 3400 13632
rect 3336 13572 3340 13628
rect 3340 13572 3396 13628
rect 3396 13572 3400 13628
rect 3336 13568 3400 13572
rect 3416 13628 3480 13632
rect 3416 13572 3420 13628
rect 3420 13572 3476 13628
rect 3476 13572 3480 13628
rect 3416 13568 3480 13572
rect 7624 13628 7688 13632
rect 7624 13572 7628 13628
rect 7628 13572 7684 13628
rect 7684 13572 7688 13628
rect 7624 13568 7688 13572
rect 7704 13628 7768 13632
rect 7704 13572 7708 13628
rect 7708 13572 7764 13628
rect 7764 13572 7768 13628
rect 7704 13568 7768 13572
rect 7784 13628 7848 13632
rect 7784 13572 7788 13628
rect 7788 13572 7844 13628
rect 7844 13572 7848 13628
rect 7784 13568 7848 13572
rect 7864 13628 7928 13632
rect 7864 13572 7868 13628
rect 7868 13572 7924 13628
rect 7924 13572 7928 13628
rect 7864 13568 7928 13572
rect 12072 13628 12136 13632
rect 12072 13572 12076 13628
rect 12076 13572 12132 13628
rect 12132 13572 12136 13628
rect 12072 13568 12136 13572
rect 12152 13628 12216 13632
rect 12152 13572 12156 13628
rect 12156 13572 12212 13628
rect 12212 13572 12216 13628
rect 12152 13568 12216 13572
rect 12232 13628 12296 13632
rect 12232 13572 12236 13628
rect 12236 13572 12292 13628
rect 12292 13572 12296 13628
rect 12232 13568 12296 13572
rect 12312 13628 12376 13632
rect 12312 13572 12316 13628
rect 12316 13572 12372 13628
rect 12372 13572 12376 13628
rect 12312 13568 12376 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 16760 13628 16824 13632
rect 16760 13572 16764 13628
rect 16764 13572 16820 13628
rect 16820 13572 16824 13628
rect 16760 13568 16824 13572
rect 15148 13152 15212 13156
rect 15148 13096 15198 13152
rect 15198 13096 15212 13152
rect 15148 13092 15212 13096
rect 5400 13084 5464 13088
rect 5400 13028 5404 13084
rect 5404 13028 5460 13084
rect 5460 13028 5464 13084
rect 5400 13024 5464 13028
rect 5480 13084 5544 13088
rect 5480 13028 5484 13084
rect 5484 13028 5540 13084
rect 5540 13028 5544 13084
rect 5480 13024 5544 13028
rect 5560 13084 5624 13088
rect 5560 13028 5564 13084
rect 5564 13028 5620 13084
rect 5620 13028 5624 13084
rect 5560 13024 5624 13028
rect 5640 13084 5704 13088
rect 5640 13028 5644 13084
rect 5644 13028 5700 13084
rect 5700 13028 5704 13084
rect 5640 13024 5704 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 14536 13084 14600 13088
rect 14536 13028 14540 13084
rect 14540 13028 14596 13084
rect 14596 13028 14600 13084
rect 14536 13024 14600 13028
rect 3176 12540 3240 12544
rect 3176 12484 3180 12540
rect 3180 12484 3236 12540
rect 3236 12484 3240 12540
rect 3176 12480 3240 12484
rect 3256 12540 3320 12544
rect 3256 12484 3260 12540
rect 3260 12484 3316 12540
rect 3316 12484 3320 12540
rect 3256 12480 3320 12484
rect 3336 12540 3400 12544
rect 3336 12484 3340 12540
rect 3340 12484 3396 12540
rect 3396 12484 3400 12540
rect 3336 12480 3400 12484
rect 3416 12540 3480 12544
rect 3416 12484 3420 12540
rect 3420 12484 3476 12540
rect 3476 12484 3480 12540
rect 3416 12480 3480 12484
rect 7624 12540 7688 12544
rect 7624 12484 7628 12540
rect 7628 12484 7684 12540
rect 7684 12484 7688 12540
rect 7624 12480 7688 12484
rect 7704 12540 7768 12544
rect 7704 12484 7708 12540
rect 7708 12484 7764 12540
rect 7764 12484 7768 12540
rect 7704 12480 7768 12484
rect 7784 12540 7848 12544
rect 7784 12484 7788 12540
rect 7788 12484 7844 12540
rect 7844 12484 7848 12540
rect 7784 12480 7848 12484
rect 7864 12540 7928 12544
rect 7864 12484 7868 12540
rect 7868 12484 7924 12540
rect 7924 12484 7928 12540
rect 7864 12480 7928 12484
rect 12072 12540 12136 12544
rect 12072 12484 12076 12540
rect 12076 12484 12132 12540
rect 12132 12484 12136 12540
rect 12072 12480 12136 12484
rect 12152 12540 12216 12544
rect 12152 12484 12156 12540
rect 12156 12484 12212 12540
rect 12212 12484 12216 12540
rect 12152 12480 12216 12484
rect 12232 12540 12296 12544
rect 12232 12484 12236 12540
rect 12236 12484 12292 12540
rect 12292 12484 12296 12540
rect 12232 12480 12296 12484
rect 12312 12540 12376 12544
rect 12312 12484 12316 12540
rect 12316 12484 12372 12540
rect 12372 12484 12376 12540
rect 12312 12480 12376 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 16760 12540 16824 12544
rect 16760 12484 16764 12540
rect 16764 12484 16820 12540
rect 16820 12484 16824 12540
rect 16760 12480 16824 12484
rect 5948 12412 6012 12476
rect 8156 12412 8220 12476
rect 3740 12140 3804 12204
rect 5400 11996 5464 12000
rect 5400 11940 5404 11996
rect 5404 11940 5460 11996
rect 5460 11940 5464 11996
rect 5400 11936 5464 11940
rect 5480 11996 5544 12000
rect 5480 11940 5484 11996
rect 5484 11940 5540 11996
rect 5540 11940 5544 11996
rect 5480 11936 5544 11940
rect 5560 11996 5624 12000
rect 5560 11940 5564 11996
rect 5564 11940 5620 11996
rect 5620 11940 5624 11996
rect 5560 11936 5624 11940
rect 5640 11996 5704 12000
rect 5640 11940 5644 11996
rect 5644 11940 5700 11996
rect 5700 11940 5704 11996
rect 5640 11936 5704 11940
rect 2452 11868 2516 11932
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 14536 11996 14600 12000
rect 14536 11940 14540 11996
rect 14540 11940 14596 11996
rect 14596 11940 14600 11996
rect 14536 11936 14600 11940
rect 3176 11452 3240 11456
rect 3176 11396 3180 11452
rect 3180 11396 3236 11452
rect 3236 11396 3240 11452
rect 3176 11392 3240 11396
rect 3256 11452 3320 11456
rect 3256 11396 3260 11452
rect 3260 11396 3316 11452
rect 3316 11396 3320 11452
rect 3256 11392 3320 11396
rect 3336 11452 3400 11456
rect 3336 11396 3340 11452
rect 3340 11396 3396 11452
rect 3396 11396 3400 11452
rect 3336 11392 3400 11396
rect 3416 11452 3480 11456
rect 3416 11396 3420 11452
rect 3420 11396 3476 11452
rect 3476 11396 3480 11452
rect 3416 11392 3480 11396
rect 7624 11452 7688 11456
rect 7624 11396 7628 11452
rect 7628 11396 7684 11452
rect 7684 11396 7688 11452
rect 7624 11392 7688 11396
rect 7704 11452 7768 11456
rect 7704 11396 7708 11452
rect 7708 11396 7764 11452
rect 7764 11396 7768 11452
rect 7704 11392 7768 11396
rect 7784 11452 7848 11456
rect 7784 11396 7788 11452
rect 7788 11396 7844 11452
rect 7844 11396 7848 11452
rect 7784 11392 7848 11396
rect 7864 11452 7928 11456
rect 7864 11396 7868 11452
rect 7868 11396 7924 11452
rect 7924 11396 7928 11452
rect 7864 11392 7928 11396
rect 2820 11112 2884 11116
rect 2820 11056 2870 11112
rect 2870 11056 2884 11112
rect 2820 11052 2884 11056
rect 5400 10908 5464 10912
rect 5400 10852 5404 10908
rect 5404 10852 5460 10908
rect 5460 10852 5464 10908
rect 5400 10848 5464 10852
rect 5480 10908 5544 10912
rect 5480 10852 5484 10908
rect 5484 10852 5540 10908
rect 5540 10852 5544 10908
rect 5480 10848 5544 10852
rect 5560 10908 5624 10912
rect 5560 10852 5564 10908
rect 5564 10852 5620 10908
rect 5620 10852 5624 10908
rect 5560 10848 5624 10852
rect 5640 10908 5704 10912
rect 5640 10852 5644 10908
rect 5644 10852 5700 10908
rect 5700 10852 5704 10908
rect 5640 10848 5704 10852
rect 6500 11112 6564 11116
rect 7420 11188 7484 11252
rect 8156 11188 8220 11252
rect 12072 11452 12136 11456
rect 12072 11396 12076 11452
rect 12076 11396 12132 11452
rect 12132 11396 12136 11452
rect 12072 11392 12136 11396
rect 12152 11452 12216 11456
rect 12152 11396 12156 11452
rect 12156 11396 12212 11452
rect 12212 11396 12216 11452
rect 12152 11392 12216 11396
rect 12232 11452 12296 11456
rect 12232 11396 12236 11452
rect 12236 11396 12292 11452
rect 12292 11396 12296 11452
rect 12232 11392 12296 11396
rect 12312 11452 12376 11456
rect 12312 11396 12316 11452
rect 12316 11396 12372 11452
rect 12372 11396 12376 11452
rect 12312 11392 12376 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 16760 11452 16824 11456
rect 16760 11396 16764 11452
rect 16764 11396 16820 11452
rect 16820 11396 16824 11452
rect 16760 11392 16824 11396
rect 14780 11324 14844 11388
rect 6500 11056 6514 11112
rect 6514 11056 6564 11112
rect 6500 11052 6564 11056
rect 8156 11052 8220 11116
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 14536 10908 14600 10912
rect 14536 10852 14540 10908
rect 14540 10852 14596 10908
rect 14596 10852 14600 10908
rect 14536 10848 14600 10852
rect 3176 10364 3240 10368
rect 3176 10308 3180 10364
rect 3180 10308 3236 10364
rect 3236 10308 3240 10364
rect 3176 10304 3240 10308
rect 3256 10364 3320 10368
rect 3256 10308 3260 10364
rect 3260 10308 3316 10364
rect 3316 10308 3320 10364
rect 3256 10304 3320 10308
rect 3336 10364 3400 10368
rect 3336 10308 3340 10364
rect 3340 10308 3396 10364
rect 3396 10308 3400 10364
rect 3336 10304 3400 10308
rect 3416 10364 3480 10368
rect 3416 10308 3420 10364
rect 3420 10308 3476 10364
rect 3476 10308 3480 10364
rect 3416 10304 3480 10308
rect 7624 10364 7688 10368
rect 7624 10308 7628 10364
rect 7628 10308 7684 10364
rect 7684 10308 7688 10364
rect 7624 10304 7688 10308
rect 7704 10364 7768 10368
rect 7704 10308 7708 10364
rect 7708 10308 7764 10364
rect 7764 10308 7768 10364
rect 7704 10304 7768 10308
rect 7784 10364 7848 10368
rect 7784 10308 7788 10364
rect 7788 10308 7844 10364
rect 7844 10308 7848 10364
rect 7784 10304 7848 10308
rect 7864 10364 7928 10368
rect 7864 10308 7868 10364
rect 7868 10308 7924 10364
rect 7924 10308 7928 10364
rect 7864 10304 7928 10308
rect 12072 10364 12136 10368
rect 12072 10308 12076 10364
rect 12076 10308 12132 10364
rect 12132 10308 12136 10364
rect 12072 10304 12136 10308
rect 12152 10364 12216 10368
rect 12152 10308 12156 10364
rect 12156 10308 12212 10364
rect 12212 10308 12216 10364
rect 12152 10304 12216 10308
rect 12232 10364 12296 10368
rect 12232 10308 12236 10364
rect 12236 10308 12292 10364
rect 12292 10308 12296 10364
rect 12232 10304 12296 10308
rect 12312 10364 12376 10368
rect 12312 10308 12316 10364
rect 12316 10308 12372 10364
rect 12372 10308 12376 10364
rect 12312 10304 12376 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 16760 10364 16824 10368
rect 16760 10308 16764 10364
rect 16764 10308 16820 10364
rect 16820 10308 16824 10364
rect 16760 10304 16824 10308
rect 3556 9692 3620 9756
rect 4108 9752 4172 9756
rect 4108 9696 4122 9752
rect 4122 9696 4172 9752
rect 4108 9692 4172 9696
rect 5400 9820 5464 9824
rect 5400 9764 5404 9820
rect 5404 9764 5460 9820
rect 5460 9764 5464 9820
rect 5400 9760 5464 9764
rect 5480 9820 5544 9824
rect 5480 9764 5484 9820
rect 5484 9764 5540 9820
rect 5540 9764 5544 9820
rect 5480 9760 5544 9764
rect 5560 9820 5624 9824
rect 5560 9764 5564 9820
rect 5564 9764 5620 9820
rect 5620 9764 5624 9820
rect 5560 9760 5624 9764
rect 5640 9820 5704 9824
rect 5640 9764 5644 9820
rect 5644 9764 5700 9820
rect 5700 9764 5704 9820
rect 5640 9760 5704 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 14536 9820 14600 9824
rect 14536 9764 14540 9820
rect 14540 9764 14596 9820
rect 14596 9764 14600 9820
rect 14536 9760 14600 9764
rect 12940 9752 13004 9756
rect 12940 9696 12954 9752
rect 12954 9696 13004 9752
rect 12940 9692 13004 9696
rect 3176 9276 3240 9280
rect 3176 9220 3180 9276
rect 3180 9220 3236 9276
rect 3236 9220 3240 9276
rect 3176 9216 3240 9220
rect 3256 9276 3320 9280
rect 3256 9220 3260 9276
rect 3260 9220 3316 9276
rect 3316 9220 3320 9276
rect 3256 9216 3320 9220
rect 3336 9276 3400 9280
rect 3336 9220 3340 9276
rect 3340 9220 3396 9276
rect 3396 9220 3400 9276
rect 3336 9216 3400 9220
rect 3416 9276 3480 9280
rect 3416 9220 3420 9276
rect 3420 9220 3476 9276
rect 3476 9220 3480 9276
rect 3416 9216 3480 9220
rect 7624 9276 7688 9280
rect 7624 9220 7628 9276
rect 7628 9220 7684 9276
rect 7684 9220 7688 9276
rect 7624 9216 7688 9220
rect 7704 9276 7768 9280
rect 7704 9220 7708 9276
rect 7708 9220 7764 9276
rect 7764 9220 7768 9276
rect 7704 9216 7768 9220
rect 7784 9276 7848 9280
rect 7784 9220 7788 9276
rect 7788 9220 7844 9276
rect 7844 9220 7848 9276
rect 7784 9216 7848 9220
rect 7864 9276 7928 9280
rect 7864 9220 7868 9276
rect 7868 9220 7924 9276
rect 7924 9220 7928 9276
rect 7864 9216 7928 9220
rect 9444 9284 9508 9348
rect 17172 9284 17236 9348
rect 12072 9276 12136 9280
rect 12072 9220 12076 9276
rect 12076 9220 12132 9276
rect 12132 9220 12136 9276
rect 12072 9216 12136 9220
rect 12152 9276 12216 9280
rect 12152 9220 12156 9276
rect 12156 9220 12212 9276
rect 12212 9220 12216 9276
rect 12152 9216 12216 9220
rect 12232 9276 12296 9280
rect 12232 9220 12236 9276
rect 12236 9220 12292 9276
rect 12292 9220 12296 9276
rect 12232 9216 12296 9220
rect 12312 9276 12376 9280
rect 12312 9220 12316 9276
rect 12316 9220 12372 9276
rect 12372 9220 12376 9276
rect 12312 9216 12376 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 16760 9276 16824 9280
rect 16760 9220 16764 9276
rect 16764 9220 16820 9276
rect 16820 9220 16824 9276
rect 16760 9216 16824 9220
rect 4844 8876 4908 8940
rect 3004 8800 3068 8804
rect 3004 8744 3018 8800
rect 3018 8744 3068 8800
rect 3004 8740 3068 8744
rect 5212 8740 5276 8804
rect 5400 8732 5464 8736
rect 5400 8676 5404 8732
rect 5404 8676 5460 8732
rect 5460 8676 5464 8732
rect 5400 8672 5464 8676
rect 5480 8732 5544 8736
rect 5480 8676 5484 8732
rect 5484 8676 5540 8732
rect 5540 8676 5544 8732
rect 5480 8672 5544 8676
rect 5560 8732 5624 8736
rect 5560 8676 5564 8732
rect 5564 8676 5620 8732
rect 5620 8676 5624 8732
rect 5560 8672 5624 8676
rect 5640 8732 5704 8736
rect 5640 8676 5644 8732
rect 5644 8676 5700 8732
rect 5700 8676 5704 8732
rect 5640 8672 5704 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 14536 8732 14600 8736
rect 14536 8676 14540 8732
rect 14540 8676 14596 8732
rect 14596 8676 14600 8732
rect 14536 8672 14600 8676
rect 2636 8332 2700 8396
rect 9260 8468 9324 8532
rect 14780 8468 14844 8532
rect 3176 8188 3240 8192
rect 3176 8132 3180 8188
rect 3180 8132 3236 8188
rect 3236 8132 3240 8188
rect 3176 8128 3240 8132
rect 3256 8188 3320 8192
rect 3256 8132 3260 8188
rect 3260 8132 3316 8188
rect 3316 8132 3320 8188
rect 3256 8128 3320 8132
rect 3336 8188 3400 8192
rect 3336 8132 3340 8188
rect 3340 8132 3396 8188
rect 3396 8132 3400 8188
rect 3336 8128 3400 8132
rect 3416 8188 3480 8192
rect 3416 8132 3420 8188
rect 3420 8132 3476 8188
rect 3476 8132 3480 8188
rect 3416 8128 3480 8132
rect 7624 8188 7688 8192
rect 7624 8132 7628 8188
rect 7628 8132 7684 8188
rect 7684 8132 7688 8188
rect 7624 8128 7688 8132
rect 7704 8188 7768 8192
rect 7704 8132 7708 8188
rect 7708 8132 7764 8188
rect 7764 8132 7768 8188
rect 7704 8128 7768 8132
rect 7784 8188 7848 8192
rect 7784 8132 7788 8188
rect 7788 8132 7844 8188
rect 7844 8132 7848 8188
rect 7784 8128 7848 8132
rect 7864 8188 7928 8192
rect 7864 8132 7868 8188
rect 7868 8132 7924 8188
rect 7924 8132 7928 8188
rect 7864 8128 7928 8132
rect 12072 8188 12136 8192
rect 12072 8132 12076 8188
rect 12076 8132 12132 8188
rect 12132 8132 12136 8188
rect 12072 8128 12136 8132
rect 12152 8188 12216 8192
rect 12152 8132 12156 8188
rect 12156 8132 12212 8188
rect 12212 8132 12216 8188
rect 12152 8128 12216 8132
rect 12232 8188 12296 8192
rect 12232 8132 12236 8188
rect 12236 8132 12292 8188
rect 12292 8132 12296 8188
rect 12232 8128 12296 8132
rect 12312 8188 12376 8192
rect 12312 8132 12316 8188
rect 12316 8132 12372 8188
rect 12372 8132 12376 8188
rect 12312 8128 12376 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 16760 8188 16824 8192
rect 16760 8132 16764 8188
rect 16764 8132 16820 8188
rect 16820 8132 16824 8188
rect 16760 8128 16824 8132
rect 3740 7924 3804 7988
rect 5400 7644 5464 7648
rect 5400 7588 5404 7644
rect 5404 7588 5460 7644
rect 5460 7588 5464 7644
rect 5400 7584 5464 7588
rect 5480 7644 5544 7648
rect 5480 7588 5484 7644
rect 5484 7588 5540 7644
rect 5540 7588 5544 7644
rect 5480 7584 5544 7588
rect 5560 7644 5624 7648
rect 5560 7588 5564 7644
rect 5564 7588 5620 7644
rect 5620 7588 5624 7644
rect 5560 7584 5624 7588
rect 5640 7644 5704 7648
rect 5640 7588 5644 7644
rect 5644 7588 5700 7644
rect 5700 7588 5704 7644
rect 5640 7584 5704 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 14536 7644 14600 7648
rect 14536 7588 14540 7644
rect 14540 7588 14596 7644
rect 14596 7588 14600 7644
rect 14536 7584 14600 7588
rect 4292 7516 4356 7580
rect 4660 7516 4724 7580
rect 5948 7380 6012 7444
rect 4844 7108 4908 7172
rect 3176 7100 3240 7104
rect 3176 7044 3180 7100
rect 3180 7044 3236 7100
rect 3236 7044 3240 7100
rect 3176 7040 3240 7044
rect 3256 7100 3320 7104
rect 3256 7044 3260 7100
rect 3260 7044 3316 7100
rect 3316 7044 3320 7100
rect 3256 7040 3320 7044
rect 3336 7100 3400 7104
rect 3336 7044 3340 7100
rect 3340 7044 3396 7100
rect 3396 7044 3400 7100
rect 3336 7040 3400 7044
rect 3416 7100 3480 7104
rect 3416 7044 3420 7100
rect 3420 7044 3476 7100
rect 3476 7044 3480 7100
rect 3416 7040 3480 7044
rect 7624 7100 7688 7104
rect 7624 7044 7628 7100
rect 7628 7044 7684 7100
rect 7684 7044 7688 7100
rect 7624 7040 7688 7044
rect 7704 7100 7768 7104
rect 7704 7044 7708 7100
rect 7708 7044 7764 7100
rect 7764 7044 7768 7100
rect 7704 7040 7768 7044
rect 7784 7100 7848 7104
rect 7784 7044 7788 7100
rect 7788 7044 7844 7100
rect 7844 7044 7848 7100
rect 7784 7040 7848 7044
rect 7864 7100 7928 7104
rect 7864 7044 7868 7100
rect 7868 7044 7924 7100
rect 7924 7044 7928 7100
rect 7864 7040 7928 7044
rect 12072 7100 12136 7104
rect 12072 7044 12076 7100
rect 12076 7044 12132 7100
rect 12132 7044 12136 7100
rect 12072 7040 12136 7044
rect 12152 7100 12216 7104
rect 12152 7044 12156 7100
rect 12156 7044 12212 7100
rect 12212 7044 12216 7100
rect 12152 7040 12216 7044
rect 12232 7100 12296 7104
rect 12232 7044 12236 7100
rect 12236 7044 12292 7100
rect 12292 7044 12296 7100
rect 12232 7040 12296 7044
rect 12312 7100 12376 7104
rect 12312 7044 12316 7100
rect 12316 7044 12372 7100
rect 12372 7044 12376 7100
rect 12312 7040 12376 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 16760 7100 16824 7104
rect 16760 7044 16764 7100
rect 16764 7044 16820 7100
rect 16820 7044 16824 7100
rect 16760 7040 16824 7044
rect 2452 6972 2516 7036
rect 5212 6972 5276 7036
rect 4108 6896 4172 6900
rect 4108 6840 4122 6896
rect 4122 6840 4172 6896
rect 4108 6836 4172 6840
rect 3004 6700 3068 6764
rect 5400 6556 5464 6560
rect 5400 6500 5404 6556
rect 5404 6500 5460 6556
rect 5460 6500 5464 6556
rect 5400 6496 5464 6500
rect 5480 6556 5544 6560
rect 5480 6500 5484 6556
rect 5484 6500 5540 6556
rect 5540 6500 5544 6556
rect 5480 6496 5544 6500
rect 5560 6556 5624 6560
rect 5560 6500 5564 6556
rect 5564 6500 5620 6556
rect 5620 6500 5624 6556
rect 5560 6496 5624 6500
rect 5640 6556 5704 6560
rect 5640 6500 5644 6556
rect 5644 6500 5700 6556
rect 5700 6500 5704 6556
rect 5640 6496 5704 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 14536 6556 14600 6560
rect 14536 6500 14540 6556
rect 14540 6500 14596 6556
rect 14596 6500 14600 6556
rect 14536 6496 14600 6500
rect 5212 6428 5276 6492
rect 17724 6428 17788 6492
rect 3176 6012 3240 6016
rect 3176 5956 3180 6012
rect 3180 5956 3236 6012
rect 3236 5956 3240 6012
rect 3176 5952 3240 5956
rect 3256 6012 3320 6016
rect 3256 5956 3260 6012
rect 3260 5956 3316 6012
rect 3316 5956 3320 6012
rect 3256 5952 3320 5956
rect 3336 6012 3400 6016
rect 3336 5956 3340 6012
rect 3340 5956 3396 6012
rect 3396 5956 3400 6012
rect 3336 5952 3400 5956
rect 3416 6012 3480 6016
rect 3416 5956 3420 6012
rect 3420 5956 3476 6012
rect 3476 5956 3480 6012
rect 3416 5952 3480 5956
rect 7624 6012 7688 6016
rect 7624 5956 7628 6012
rect 7628 5956 7684 6012
rect 7684 5956 7688 6012
rect 7624 5952 7688 5956
rect 7704 6012 7768 6016
rect 7704 5956 7708 6012
rect 7708 5956 7764 6012
rect 7764 5956 7768 6012
rect 7704 5952 7768 5956
rect 7784 6012 7848 6016
rect 7784 5956 7788 6012
rect 7788 5956 7844 6012
rect 7844 5956 7848 6012
rect 7784 5952 7848 5956
rect 7864 6012 7928 6016
rect 7864 5956 7868 6012
rect 7868 5956 7924 6012
rect 7924 5956 7928 6012
rect 7864 5952 7928 5956
rect 12072 6012 12136 6016
rect 12072 5956 12076 6012
rect 12076 5956 12132 6012
rect 12132 5956 12136 6012
rect 12072 5952 12136 5956
rect 12152 6012 12216 6016
rect 12152 5956 12156 6012
rect 12156 5956 12212 6012
rect 12212 5956 12216 6012
rect 12152 5952 12216 5956
rect 12232 6012 12296 6016
rect 12232 5956 12236 6012
rect 12236 5956 12292 6012
rect 12292 5956 12296 6012
rect 12232 5952 12296 5956
rect 12312 6012 12376 6016
rect 12312 5956 12316 6012
rect 12316 5956 12372 6012
rect 12372 5956 12376 6012
rect 12312 5952 12376 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 16760 6012 16824 6016
rect 16760 5956 16764 6012
rect 16764 5956 16820 6012
rect 16820 5956 16824 6012
rect 16760 5952 16824 5956
rect 5400 5468 5464 5472
rect 5400 5412 5404 5468
rect 5404 5412 5460 5468
rect 5460 5412 5464 5468
rect 5400 5408 5464 5412
rect 5480 5468 5544 5472
rect 5480 5412 5484 5468
rect 5484 5412 5540 5468
rect 5540 5412 5544 5468
rect 5480 5408 5544 5412
rect 5560 5468 5624 5472
rect 5560 5412 5564 5468
rect 5564 5412 5620 5468
rect 5620 5412 5624 5468
rect 5560 5408 5624 5412
rect 5640 5468 5704 5472
rect 5640 5412 5644 5468
rect 5644 5412 5700 5468
rect 5700 5412 5704 5468
rect 5640 5408 5704 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 14536 5468 14600 5472
rect 14536 5412 14540 5468
rect 14540 5412 14596 5468
rect 14596 5412 14600 5468
rect 14536 5408 14600 5412
rect 7420 5340 7484 5404
rect 3176 4924 3240 4928
rect 3176 4868 3180 4924
rect 3180 4868 3236 4924
rect 3236 4868 3240 4924
rect 3176 4864 3240 4868
rect 3256 4924 3320 4928
rect 3256 4868 3260 4924
rect 3260 4868 3316 4924
rect 3316 4868 3320 4924
rect 3256 4864 3320 4868
rect 3336 4924 3400 4928
rect 3336 4868 3340 4924
rect 3340 4868 3396 4924
rect 3396 4868 3400 4924
rect 3336 4864 3400 4868
rect 3416 4924 3480 4928
rect 3416 4868 3420 4924
rect 3420 4868 3476 4924
rect 3476 4868 3480 4924
rect 3416 4864 3480 4868
rect 7624 4924 7688 4928
rect 7624 4868 7628 4924
rect 7628 4868 7684 4924
rect 7684 4868 7688 4924
rect 7624 4864 7688 4868
rect 7704 4924 7768 4928
rect 7704 4868 7708 4924
rect 7708 4868 7764 4924
rect 7764 4868 7768 4924
rect 7704 4864 7768 4868
rect 7784 4924 7848 4928
rect 7784 4868 7788 4924
rect 7788 4868 7844 4924
rect 7844 4868 7848 4924
rect 7784 4864 7848 4868
rect 7864 4924 7928 4928
rect 7864 4868 7868 4924
rect 7868 4868 7924 4924
rect 7924 4868 7928 4924
rect 7864 4864 7928 4868
rect 12072 4924 12136 4928
rect 12072 4868 12076 4924
rect 12076 4868 12132 4924
rect 12132 4868 12136 4924
rect 12072 4864 12136 4868
rect 12152 4924 12216 4928
rect 12152 4868 12156 4924
rect 12156 4868 12212 4924
rect 12212 4868 12216 4924
rect 12152 4864 12216 4868
rect 12232 4924 12296 4928
rect 12232 4868 12236 4924
rect 12236 4868 12292 4924
rect 12292 4868 12296 4924
rect 12232 4864 12296 4868
rect 12312 4924 12376 4928
rect 12312 4868 12316 4924
rect 12316 4868 12372 4924
rect 12372 4868 12376 4924
rect 12312 4864 12376 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 16760 4924 16824 4928
rect 16760 4868 16764 4924
rect 16764 4868 16820 4924
rect 16820 4868 16824 4924
rect 16760 4864 16824 4868
rect 2636 4660 2700 4724
rect 5400 4380 5464 4384
rect 5400 4324 5404 4380
rect 5404 4324 5460 4380
rect 5460 4324 5464 4380
rect 5400 4320 5464 4324
rect 5480 4380 5544 4384
rect 5480 4324 5484 4380
rect 5484 4324 5540 4380
rect 5540 4324 5544 4380
rect 5480 4320 5544 4324
rect 5560 4380 5624 4384
rect 5560 4324 5564 4380
rect 5564 4324 5620 4380
rect 5620 4324 5624 4380
rect 5560 4320 5624 4324
rect 5640 4380 5704 4384
rect 5640 4324 5644 4380
rect 5644 4324 5700 4380
rect 5700 4324 5704 4380
rect 5640 4320 5704 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 14536 4380 14600 4384
rect 14536 4324 14540 4380
rect 14540 4324 14596 4380
rect 14596 4324 14600 4380
rect 14536 4320 14600 4324
rect 2820 4176 2884 4180
rect 2820 4120 2834 4176
rect 2834 4120 2884 4176
rect 2820 4116 2884 4120
rect 16252 3980 16316 4044
rect 17172 3980 17236 4044
rect 14964 3844 15028 3908
rect 3176 3836 3240 3840
rect 3176 3780 3180 3836
rect 3180 3780 3236 3836
rect 3236 3780 3240 3836
rect 3176 3776 3240 3780
rect 3256 3836 3320 3840
rect 3256 3780 3260 3836
rect 3260 3780 3316 3836
rect 3316 3780 3320 3836
rect 3256 3776 3320 3780
rect 3336 3836 3400 3840
rect 3336 3780 3340 3836
rect 3340 3780 3396 3836
rect 3396 3780 3400 3836
rect 3336 3776 3400 3780
rect 3416 3836 3480 3840
rect 3416 3780 3420 3836
rect 3420 3780 3476 3836
rect 3476 3780 3480 3836
rect 3416 3776 3480 3780
rect 7624 3836 7688 3840
rect 7624 3780 7628 3836
rect 7628 3780 7684 3836
rect 7684 3780 7688 3836
rect 7624 3776 7688 3780
rect 7704 3836 7768 3840
rect 7704 3780 7708 3836
rect 7708 3780 7764 3836
rect 7764 3780 7768 3836
rect 7704 3776 7768 3780
rect 7784 3836 7848 3840
rect 7784 3780 7788 3836
rect 7788 3780 7844 3836
rect 7844 3780 7848 3836
rect 7784 3776 7848 3780
rect 7864 3836 7928 3840
rect 7864 3780 7868 3836
rect 7868 3780 7924 3836
rect 7924 3780 7928 3836
rect 7864 3776 7928 3780
rect 12072 3836 12136 3840
rect 12072 3780 12076 3836
rect 12076 3780 12132 3836
rect 12132 3780 12136 3836
rect 12072 3776 12136 3780
rect 12152 3836 12216 3840
rect 12152 3780 12156 3836
rect 12156 3780 12212 3836
rect 12212 3780 12216 3836
rect 12152 3776 12216 3780
rect 12232 3836 12296 3840
rect 12232 3780 12236 3836
rect 12236 3780 12292 3836
rect 12292 3780 12296 3836
rect 12232 3776 12296 3780
rect 12312 3836 12376 3840
rect 12312 3780 12316 3836
rect 12316 3780 12372 3836
rect 12372 3780 12376 3836
rect 12312 3776 12376 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 16760 3836 16824 3840
rect 16760 3780 16764 3836
rect 16764 3780 16820 3836
rect 16820 3780 16824 3836
rect 16760 3776 16824 3780
rect 8156 3572 8220 3636
rect 15148 3572 15212 3636
rect 5400 3292 5464 3296
rect 5400 3236 5404 3292
rect 5404 3236 5460 3292
rect 5460 3236 5464 3292
rect 5400 3232 5464 3236
rect 5480 3292 5544 3296
rect 5480 3236 5484 3292
rect 5484 3236 5540 3292
rect 5540 3236 5544 3292
rect 5480 3232 5544 3236
rect 5560 3292 5624 3296
rect 5560 3236 5564 3292
rect 5564 3236 5620 3292
rect 5620 3236 5624 3292
rect 5560 3232 5624 3236
rect 5640 3292 5704 3296
rect 5640 3236 5644 3292
rect 5644 3236 5700 3292
rect 5700 3236 5704 3292
rect 5640 3232 5704 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 14536 3292 14600 3296
rect 14536 3236 14540 3292
rect 14540 3236 14596 3292
rect 14596 3236 14600 3292
rect 14536 3232 14600 3236
rect 9444 3164 9508 3228
rect 3556 3028 3620 3092
rect 3176 2748 3240 2752
rect 3176 2692 3180 2748
rect 3180 2692 3236 2748
rect 3236 2692 3240 2748
rect 3176 2688 3240 2692
rect 3256 2748 3320 2752
rect 3256 2692 3260 2748
rect 3260 2692 3316 2748
rect 3316 2692 3320 2748
rect 3256 2688 3320 2692
rect 3336 2748 3400 2752
rect 3336 2692 3340 2748
rect 3340 2692 3396 2748
rect 3396 2692 3400 2748
rect 3336 2688 3400 2692
rect 3416 2748 3480 2752
rect 3416 2692 3420 2748
rect 3420 2692 3476 2748
rect 3476 2692 3480 2748
rect 3416 2688 3480 2692
rect 7624 2748 7688 2752
rect 7624 2692 7628 2748
rect 7628 2692 7684 2748
rect 7684 2692 7688 2748
rect 7624 2688 7688 2692
rect 7704 2748 7768 2752
rect 7704 2692 7708 2748
rect 7708 2692 7764 2748
rect 7764 2692 7768 2748
rect 7704 2688 7768 2692
rect 7784 2748 7848 2752
rect 7784 2692 7788 2748
rect 7788 2692 7844 2748
rect 7844 2692 7848 2748
rect 7784 2688 7848 2692
rect 7864 2748 7928 2752
rect 7864 2692 7868 2748
rect 7868 2692 7924 2748
rect 7924 2692 7928 2748
rect 7864 2688 7928 2692
rect 12072 2748 12136 2752
rect 12072 2692 12076 2748
rect 12076 2692 12132 2748
rect 12132 2692 12136 2748
rect 12072 2688 12136 2692
rect 12152 2748 12216 2752
rect 12152 2692 12156 2748
rect 12156 2692 12212 2748
rect 12212 2692 12216 2748
rect 12152 2688 12216 2692
rect 12232 2748 12296 2752
rect 12232 2692 12236 2748
rect 12236 2692 12292 2748
rect 12292 2692 12296 2748
rect 12232 2688 12296 2692
rect 12312 2748 12376 2752
rect 12312 2692 12316 2748
rect 12316 2692 12372 2748
rect 12372 2692 12376 2748
rect 12312 2688 12376 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 16760 2748 16824 2752
rect 16760 2692 16764 2748
rect 16764 2692 16820 2748
rect 16820 2692 16824 2748
rect 16760 2688 16824 2692
rect 6500 2680 6564 2684
rect 6500 2624 6514 2680
rect 6514 2624 6564 2680
rect 6500 2620 6564 2624
rect 4292 2484 4356 2548
rect 12940 2484 13004 2548
rect 9260 2348 9324 2412
rect 5400 2204 5464 2208
rect 5400 2148 5404 2204
rect 5404 2148 5460 2204
rect 5460 2148 5464 2204
rect 5400 2144 5464 2148
rect 5480 2204 5544 2208
rect 5480 2148 5484 2204
rect 5484 2148 5540 2204
rect 5540 2148 5544 2204
rect 5480 2144 5544 2148
rect 5560 2204 5624 2208
rect 5560 2148 5564 2204
rect 5564 2148 5620 2204
rect 5620 2148 5624 2204
rect 5560 2144 5624 2148
rect 5640 2204 5704 2208
rect 5640 2148 5644 2204
rect 5644 2148 5700 2204
rect 5700 2148 5704 2204
rect 5640 2144 5704 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 14536 2204 14600 2208
rect 14536 2148 14540 2204
rect 14540 2148 14596 2204
rect 14596 2148 14600 2204
rect 14536 2144 14600 2148
<< metal4 >>
rect 17723 16148 17789 16149
rect 17723 16084 17724 16148
rect 17788 16084 17789 16148
rect 17723 16083 17789 16084
rect 17726 15469 17786 16083
rect 17723 15468 17789 15469
rect 17723 15404 17724 15468
rect 17788 15404 17789 15468
rect 17723 15403 17789 15404
rect 3739 15060 3805 15061
rect 3739 14996 3740 15060
rect 3804 14996 3805 15060
rect 3739 14995 3805 14996
rect 3168 14720 3488 14736
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3168 13632 3488 14656
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 3168 12544 3488 13568
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 2451 11932 2517 11933
rect 2451 11868 2452 11932
rect 2516 11868 2517 11932
rect 2451 11867 2517 11868
rect 2454 7037 2514 11867
rect 3168 11456 3488 12480
rect 3742 12205 3802 14995
rect 5392 14176 5712 14736
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 4659 13972 4725 13973
rect 4659 13908 4660 13972
rect 4724 13908 4725 13972
rect 4659 13907 4725 13908
rect 3739 12204 3805 12205
rect 3739 12140 3740 12204
rect 3804 12140 3805 12204
rect 3739 12139 3805 12140
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 2819 11116 2885 11117
rect 2819 11052 2820 11116
rect 2884 11052 2885 11116
rect 2819 11051 2885 11052
rect 2635 8396 2701 8397
rect 2635 8332 2636 8396
rect 2700 8332 2701 8396
rect 2635 8331 2701 8332
rect 2451 7036 2517 7037
rect 2451 6972 2452 7036
rect 2516 6972 2517 7036
rect 2451 6971 2517 6972
rect 2638 4725 2698 8331
rect 2635 4724 2701 4725
rect 2635 4660 2636 4724
rect 2700 4660 2701 4724
rect 2635 4659 2701 4660
rect 2822 4181 2882 11051
rect 3168 10368 3488 11392
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3168 9280 3488 10304
rect 3555 9756 3621 9757
rect 3555 9692 3556 9756
rect 3620 9692 3621 9756
rect 3555 9691 3621 9692
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 3003 8804 3069 8805
rect 3003 8740 3004 8804
rect 3068 8740 3069 8804
rect 3003 8739 3069 8740
rect 3006 6765 3066 8739
rect 3168 8192 3488 9216
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 3168 7104 3488 8128
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3003 6764 3069 6765
rect 3003 6700 3004 6764
rect 3068 6700 3069 6764
rect 3003 6699 3069 6700
rect 3168 6016 3488 7040
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 3168 4928 3488 5952
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 2819 4180 2885 4181
rect 2819 4116 2820 4180
rect 2884 4116 2885 4180
rect 2819 4115 2885 4116
rect 3168 3840 3488 4864
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 3168 2752 3488 3776
rect 3558 3093 3618 9691
rect 3742 7989 3802 12139
rect 4107 9756 4173 9757
rect 4107 9692 4108 9756
rect 4172 9692 4173 9756
rect 4107 9691 4173 9692
rect 3739 7988 3805 7989
rect 3739 7924 3740 7988
rect 3804 7924 3805 7988
rect 3739 7923 3805 7924
rect 4110 6901 4170 9691
rect 4662 7581 4722 13907
rect 5392 13088 5712 14112
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 5392 12000 5712 13024
rect 7616 14720 7936 14736
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 7616 13632 7936 14656
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 7616 12544 7936 13568
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 5947 12476 6013 12477
rect 5947 12412 5948 12476
rect 6012 12412 6013 12476
rect 5947 12411 6013 12412
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5392 10912 5712 11936
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 9824 5712 10848
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 4843 8940 4909 8941
rect 4843 8876 4844 8940
rect 4908 8876 4909 8940
rect 4843 8875 4909 8876
rect 4291 7580 4357 7581
rect 4291 7516 4292 7580
rect 4356 7516 4357 7580
rect 4291 7515 4357 7516
rect 4659 7580 4725 7581
rect 4659 7516 4660 7580
rect 4724 7516 4725 7580
rect 4659 7515 4725 7516
rect 4107 6900 4173 6901
rect 4107 6836 4108 6900
rect 4172 6836 4173 6900
rect 4107 6835 4173 6836
rect 3555 3092 3621 3093
rect 3555 3028 3556 3092
rect 3620 3028 3621 3092
rect 3555 3027 3621 3028
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2128 3488 2688
rect 4294 2549 4354 7515
rect 4846 7173 4906 8875
rect 5211 8804 5277 8805
rect 5211 8740 5212 8804
rect 5276 8740 5277 8804
rect 5211 8739 5277 8740
rect 4843 7172 4909 7173
rect 4843 7108 4844 7172
rect 4908 7108 4909 7172
rect 4843 7107 4909 7108
rect 5214 7037 5274 8739
rect 5392 8736 5712 9760
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 7648 5712 8672
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5211 7036 5277 7037
rect 5211 6972 5212 7036
rect 5276 6972 5277 7036
rect 5211 6971 5277 6972
rect 5214 6493 5274 6971
rect 5392 6560 5712 7584
rect 5950 7445 6010 12411
rect 7616 11456 7936 12480
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 8155 12476 8221 12477
rect 8155 12412 8156 12476
rect 8220 12412 8221 12476
rect 8155 12411 8221 12412
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7419 11252 7485 11253
rect 7419 11188 7420 11252
rect 7484 11188 7485 11252
rect 7419 11187 7485 11188
rect 6499 11116 6565 11117
rect 6499 11052 6500 11116
rect 6564 11052 6565 11116
rect 6499 11051 6565 11052
rect 5947 7444 6013 7445
rect 5947 7380 5948 7444
rect 6012 7380 6013 7444
rect 5947 7379 6013 7380
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5211 6492 5277 6493
rect 5211 6428 5212 6492
rect 5276 6428 5277 6492
rect 5211 6427 5277 6428
rect 5392 5472 5712 6496
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 5392 4384 5712 5408
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 5392 3296 5712 4320
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 4291 2548 4357 2549
rect 4291 2484 4292 2548
rect 4356 2484 4357 2548
rect 4291 2483 4357 2484
rect 5392 2208 5712 3232
rect 6502 2685 6562 11051
rect 7422 5405 7482 11187
rect 7616 10368 7936 11392
rect 8158 11253 8218 12411
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 8155 11252 8221 11253
rect 8155 11188 8156 11252
rect 8220 11188 8221 11252
rect 8155 11187 8221 11188
rect 8155 11116 8221 11117
rect 8155 11052 8156 11116
rect 8220 11052 8221 11116
rect 8155 11051 8221 11052
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7616 9280 7936 10304
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7616 8192 7936 9216
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7616 7104 7936 8128
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 6016 7936 7040
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7419 5404 7485 5405
rect 7419 5340 7420 5404
rect 7484 5340 7485 5404
rect 7419 5339 7485 5340
rect 7616 4928 7936 5952
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 3840 7936 4864
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 7616 2752 7936 3776
rect 8158 3637 8218 11051
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9443 9348 9509 9349
rect 9443 9284 9444 9348
rect 9508 9284 9509 9348
rect 9443 9283 9509 9284
rect 9259 8532 9325 8533
rect 9259 8468 9260 8532
rect 9324 8468 9325 8532
rect 9259 8467 9325 8468
rect 8155 3636 8221 3637
rect 8155 3572 8156 3636
rect 8220 3572 8221 3636
rect 8155 3571 8221 3572
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 6499 2684 6565 2685
rect 6499 2620 6500 2684
rect 6564 2620 6565 2684
rect 6499 2619 6565 2620
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2128 5712 2144
rect 7616 2128 7936 2688
rect 9262 2413 9322 8467
rect 9446 3229 9506 9283
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9443 3228 9509 3229
rect 9443 3164 9444 3228
rect 9508 3164 9509 3228
rect 9443 3163 9509 3164
rect 9259 2412 9325 2413
rect 9259 2348 9260 2412
rect 9324 2348 9325 2412
rect 9259 2347 9325 2348
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12064 14720 12384 14736
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 13632 12384 14656
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 12064 12544 12384 13568
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 12064 11456 12384 12480
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 10368 12384 11392
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 9280 12384 10304
rect 14288 14176 14608 14736
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 14288 13088 14608 14112
rect 16512 14720 16832 14736
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 14963 13836 15029 13837
rect 14963 13772 14964 13836
rect 15028 13772 15029 13836
rect 14963 13771 15029 13772
rect 16251 13836 16317 13837
rect 16251 13772 16252 13836
rect 16316 13772 16317 13836
rect 16251 13771 16317 13772
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 14288 12000 14608 13024
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 14288 10912 14608 11936
rect 14779 11388 14845 11389
rect 14779 11324 14780 11388
rect 14844 11324 14845 11388
rect 14779 11323 14845 11324
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 9824 14608 10848
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 12939 9756 13005 9757
rect 12939 9692 12940 9756
rect 13004 9692 13005 9756
rect 12939 9691 13005 9692
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 8192 12384 9216
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 7104 12384 8128
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 6016 12384 7040
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 4928 12384 5952
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 3840 12384 4864
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 2752 12384 3776
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 12064 2128 12384 2688
rect 12942 2549 13002 9691
rect 14288 8736 14608 9760
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 14288 7648 14608 8672
rect 14782 8533 14842 11323
rect 14779 8532 14845 8533
rect 14779 8468 14780 8532
rect 14844 8468 14845 8532
rect 14779 8467 14845 8468
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 6560 14608 7584
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 14288 5472 14608 6496
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 14288 4384 14608 5408
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 14288 3296 14608 4320
rect 14966 3909 15026 13771
rect 15147 13156 15213 13157
rect 15147 13092 15148 13156
rect 15212 13092 15213 13156
rect 15147 13091 15213 13092
rect 14963 3908 15029 3909
rect 14963 3844 14964 3908
rect 15028 3844 15029 3908
rect 14963 3843 15029 3844
rect 15150 3637 15210 13091
rect 16254 4045 16314 13771
rect 16512 13632 16832 14656
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 12544 16832 13568
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 16512 11456 16832 12480
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 10368 16832 11392
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 16512 9280 16832 10304
rect 17171 9348 17237 9349
rect 17171 9284 17172 9348
rect 17236 9284 17237 9348
rect 17171 9283 17237 9284
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 8192 16832 9216
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 16512 7104 16832 8128
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16512 6016 16832 7040
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16512 4928 16832 5952
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 16251 4044 16317 4045
rect 16251 3980 16252 4044
rect 16316 3980 16317 4044
rect 16251 3979 16317 3980
rect 16512 3840 16832 4864
rect 17174 4045 17234 9283
rect 17726 6493 17786 15403
rect 17723 6492 17789 6493
rect 17723 6428 17724 6492
rect 17788 6428 17789 6492
rect 17723 6427 17789 6428
rect 17171 4044 17237 4045
rect 17171 3980 17172 4044
rect 17236 3980 17237 4044
rect 17171 3979 17237 3980
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 15147 3636 15213 3637
rect 15147 3572 15148 3636
rect 15212 3572 15213 3636
rect 15147 3571 15213 3572
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 12939 2548 13005 2549
rect 12939 2484 12940 2548
rect 13004 2484 13005 2548
rect 12939 2483 13005 2484
rect 14288 2208 14608 3232
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 14288 2128 14608 2144
rect 16512 2752 16832 3776
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 16512 2128 16832 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17204 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1649977179
transform 1 0 15088 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform 1 0 2760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform 1 0 1564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform -1 0 1840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform -1 0 2760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform -1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform -1 0 1748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform -1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1649977179
transform 1 0 2208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform 1 0 2024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform -1 0 2024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform -1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform -1 0 1564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform 1 0 1564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1649977179
transform -1 0 1840 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1649977179
transform -1 0 1748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1649977179
transform -1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1649977179
transform -1 0 16836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1649977179
transform -1 0 16192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1649977179
transform 1 0 13248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1649977179
transform 1 0 12880 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform 1 0 11684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform -1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform -1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform 1 0 17296 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform 1 0 17664 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1649977179
transform 1 0 13064 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform 1 0 18032 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform -1 0 18492 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 18584 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform -1 0 18492 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform -1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform -1 0 18584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform -1 0 18492 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1649977179
transform -1 0 15364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 14720 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 16468 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 9936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15548 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13248 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 10580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 13984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 12052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8096 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4968 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5704 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8004 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9476 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 15824 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13248 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18492 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16836 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 17664 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 17020 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 4784 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5152 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1649977179
transform 1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 2024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 1472 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3772 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 2392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 9752 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4232 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 2576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 2760 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 2668 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 1472 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 2668 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 4232 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 3864 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 6256 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 2668 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__S
timestamp 1649977179
transform -1 0 5152 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 2576 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 2760 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 1472 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3496 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 2668 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8280 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6440 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 4232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3036 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 7452 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 8096 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7728 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11500 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8740 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 7820 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6808 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11776 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11776 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10120 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 2576 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 2760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 1472 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 2944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9936 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 4968 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 18124 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 17204 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12328 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13156 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14352 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 16652 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16100 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13892 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14076 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 16100 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 18492 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 18492 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 16468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14720 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 17020 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 18032 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 17848 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16744 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16928 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 16560 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform 1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1649977179
transform -1 0 6716 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_171
timestamp 1649977179
transform 1 0 16836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_173
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_119
timestamp 1649977179
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_140
timestamp 1649977179
transform 1 0 13984 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1649977179
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_135
timestamp 1649977179
transform 1 0 13524 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_17
timestamp 1649977179
transform 1 0 2668 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_59
timestamp 1649977179
transform 1 0 6532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_163
timestamp 1649977179
transform 1 0 16100 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1649977179
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_11
timestamp 1649977179
transform 1 0 2116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_23
timestamp 1649977179
transform 1 0 3220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7912 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_135
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_61 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_83
timestamp 1649977179
transform 1 0 8740 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_87
timestamp 1649977179
transform 1 0 9108 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1649977179
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_18
timestamp 1649977179
transform 1 0 2760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1649977179
transform 1 0 4324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_89
timestamp 1649977179
transform 1 0 9292 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_95
timestamp 1649977179
transform 1 0 9844 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_79 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8372 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1649977179
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1649977179
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_108
timestamp 1649977179
transform 1 0 11040 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_127
timestamp 1649977179
transform 1 0 12788 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_135
timestamp 1649977179
transform 1 0 13524 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1649977179
transform 1 0 1932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_82
timestamp 1649977179
transform 1 0 8648 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_109
timestamp 1649977179
transform 1 0 11132 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_130
timestamp 1649977179
transform 1 0 13064 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_20
timestamp 1649977179
transform 1 0 2944 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_56
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_100
timestamp 1649977179
transform 1 0 10304 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_103
timestamp 1649977179
transform 1 0 10580 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_115
timestamp 1649977179
transform 1 0 11684 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_119 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_124
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_128
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_143
timestamp 1649977179
transform 1 0 14260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_19
timestamp 1649977179
transform 1 0 2852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_53
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1649977179
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_13
timestamp 1649977179
transform 1 0 2300 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_17
timestamp 1649977179
transform 1 0 2668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1649977179
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_99
timestamp 1649977179
transform 1 0 10212 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_118
timestamp 1649977179
transform 1 0 11960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_175
timestamp 1649977179
transform 1 0 17204 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_28
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_49
timestamp 1649977179
transform 1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_107
timestamp 1649977179
transform 1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_126
timestamp 1649977179
transform 1 0 12696 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_14
timestamp 1649977179
transform 1 0 2392 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_47
timestamp 1649977179
transform 1 0 5428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_118
timestamp 1649977179
transform 1 0 11960 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_135
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_171
timestamp 1649977179
transform 1 0 16836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_96
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_109
timestamp 1649977179
transform 1 0 11132 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_124
timestamp 1649977179
transform 1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1649977179
transform 1 0 12972 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_141
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_147
timestamp 1649977179
transform 1 0 14628 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_178
timestamp 1649977179
transform 1 0 17480 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_186
timestamp 1649977179
transform 1 0 18216 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1649977179
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_105
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_113
timestamp 1649977179
transform 1 0 11500 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_152 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15088 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_164
timestamp 1649977179
transform 1 0 16192 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_172
timestamp 1649977179
transform 1 0 16928 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_188
timestamp 1649977179
transform 1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 1649977179
transform 1 0 1932 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_12
timestamp 1649977179
transform 1 0 2208 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_18
timestamp 1649977179
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_30
timestamp 1649977179
transform 1 0 3864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_42
timestamp 1649977179
transform 1 0 4968 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_77
timestamp 1649977179
transform 1 0 8188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_89
timestamp 1649977179
transform 1 0 9292 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_94
timestamp 1649977179
transform 1 0 9752 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_138
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_143
timestamp 1649977179
transform 1 0 14260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_155
timestamp 1649977179
transform 1 0 15364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_66
timestamp 1649977179
transform 1 0 7176 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_78
timestamp 1649977179
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_129
timestamp 1649977179
transform 1 0 12972 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1649977179
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_149
timestamp 1649977179
transform 1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_154
timestamp 1649977179
transform 1 0 15272 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_166
timestamp 1649977179
transform 1 0 16376 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_178
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_61
timestamp 1649977179
transform 1 0 6716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_73
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_85
timestamp 1649977179
transform 1 0 8924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_97
timestamp 1649977179
transform 1 0 10028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_175
timestamp 1649977179
transform 1 0 17204 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_187
timestamp 1649977179
transform 1 0 18308 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_46
timestamp 1649977179
transform 1 0 5336 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_54
timestamp 1649977179
transform 1 0 6072 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_57
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_69
timestamp 1649977179
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_113
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_125
timestamp 1649977179
transform 1 0 12604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1649977179
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_169
timestamp 1649977179
transform 1 0 16652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_181
timestamp 1649977179
transform 1 0 17756 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _17_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6900 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1649977179
transform -1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1649977179
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1649977179
transform 1 0 9384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1649977179
transform -1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1649977179
transform -1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1649977179
transform -1 0 3496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1649977179
transform 1 0 16560 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1649977179
transform -1 0 12052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1649977179
transform -1 0 17296 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1649977179
transform 1 0 2116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _34_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1649977179
transform -1 0 15088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1649977179
transform -1 0 4140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1649977179
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1649977179
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1649977179
transform -1 0 2116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1649977179
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1649977179
transform -1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1649977179
transform -1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1649977179
transform -1 0 2116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1649977179
transform -1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1649977179
transform -1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1649977179
transform -1 0 2024 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1649977179
transform -1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1649977179
transform -1 0 2392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1649977179
transform -1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1649977179
transform -1 0 2116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1649977179
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1649977179
transform -1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1649977179
transform -1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1649977179
transform 1 0 16744 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1649977179
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1649977179
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1649977179
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1649977179
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1649977179
transform 1 0 18032 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1649977179
transform 1 0 17848 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1649977179
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1649977179
transform 1 0 18216 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1649977179
transform 1 0 17848 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1649977179
transform 1 0 18216 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1649977179
transform 1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1649977179
transform 1 0 17848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1649977179
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1649977179
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13248 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14536 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10488 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 15088 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13432 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17020 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15916 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6256 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8096 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13616 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9844 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11408 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11500 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9200 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 10580 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14444 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10488 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10488 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11040 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7544 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7084 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9108 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6624 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4416 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 8372 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4784 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7360 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4600 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6532 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 5888 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8832 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8096 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8464 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9844 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4416 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6624 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9108 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13524 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 12880 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11316 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16376 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 17020 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13064 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12972 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11684 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 17020 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16376 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 14904 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15180 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15548 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15548 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17480 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17020 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15364 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13064 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 13524 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12880 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12788 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3956 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4232 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4048 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5336 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4508 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2760 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3956 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3220 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3404 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2576 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3680 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3404 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 2760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 1932 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2024 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2484 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3680 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4968 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2668 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3128 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2852 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2576 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 2576 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2668 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3496 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7268 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6348 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5428 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5520 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4784 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3404 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4784 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4600 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4600 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4784 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8096 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7268 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7176 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform -1 0 5428 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5428 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6440 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5980 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7912 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8924 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7636 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6992 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform -1 0 6256 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6900 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7176 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6440 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6440 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11960 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10120 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9292 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3956 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4784 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8740 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5980 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8832 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9476 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5152 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform -1 0 16468 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5612 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16192 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12052 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12328 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11132 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10672 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15364 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform -1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform -1 0 13616 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12420 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16928 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17296 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16376 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16100 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15824 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15732 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17204 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17020 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15088 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18032 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17112 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17756 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform -1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17020 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16928 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15732 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1649977179
transform -1 0 2208 0 1 2176
box -38 -48 590 592
<< labels >>
flabel metal2 s 1122 16400 1178 17200 0 FreeSans 224 90 0 0 IO_ISOL_N
port 0 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 SC_IN_BOT
port 1 nsew signal input
flabel metal2 s 3330 16400 3386 17200 0 FreeSans 224 90 0 0 SC_IN_TOP
port 2 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 3 nsew signal tristate
flabel metal2 s 5538 16400 5594 17200 0 FreeSans 224 90 0 0 SC_OUT_TOP
port 4 nsew signal tristate
flabel metal4 s 5392 2128 5712 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 9840 2128 10160 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 14288 2128 14608 14736 0 FreeSans 1920 90 0 0 VGND
port 5 nsew ground bidirectional
flabel metal4 s 3168 2128 3488 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 7616 2128 7936 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 12064 2128 12384 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal4 s 16512 2128 16832 14736 0 FreeSans 1920 90 0 0 VPWR
port 6 nsew power bidirectional
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 bottom_grid_pin_0_
port 7 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 bottom_grid_pin_10_
port 8 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 bottom_grid_pin_11_
port 9 nsew signal tristate
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 bottom_grid_pin_12_
port 10 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 bottom_grid_pin_13_
port 11 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 bottom_grid_pin_14_
port 12 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 bottom_grid_pin_15_
port 13 nsew signal tristate
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 bottom_grid_pin_1_
port 14 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_grid_pin_2_
port 15 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 bottom_grid_pin_3_
port 16 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 bottom_grid_pin_4_
port 17 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 bottom_grid_pin_5_
port 18 nsew signal tristate
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 bottom_grid_pin_6_
port 19 nsew signal tristate
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 bottom_grid_pin_7_
port 20 nsew signal tristate
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 bottom_grid_pin_8_
port 21 nsew signal tristate
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 bottom_grid_pin_9_
port 22 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0__pin_0_
port 23 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0__pin_1_lower
port 24 nsew signal tristate
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 bottom_width_0_height_0__pin_1_upper
port 25 nsew signal tristate
flabel metal2 s 7746 16400 7802 17200 0 FreeSans 224 90 0 0 ccff_head
port 26 nsew signal input
flabel metal2 s 9954 16400 10010 17200 0 FreeSans 224 90 0 0 ccff_tail
port 27 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 28 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 29 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 30 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 31 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 32 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 33 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 34 nsew signal input
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 35 nsew signal input
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 36 nsew signal input
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 37 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 38 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 39 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 40 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 41 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 42 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 43 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 44 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 45 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 46 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 47 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 48 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 49 nsew signal tristate
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 50 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 51 nsew signal tristate
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 52 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 53 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 54 nsew signal tristate
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 55 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 56 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 57 nsew signal tristate
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 58 nsew signal tristate
flabel metal3 s 0 1096 800 1216 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 59 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 60 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 61 nsew signal tristate
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 62 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 63 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 64 nsew signal tristate
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 65 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 66 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 67 nsew signal tristate
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 68 nsew signal input
flabel metal3 s 19200 12792 20000 12912 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 69 nsew signal input
flabel metal3 s 19200 13200 20000 13320 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 70 nsew signal input
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 71 nsew signal input
flabel metal3 s 19200 14016 20000 14136 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 72 nsew signal input
flabel metal3 s 19200 14424 20000 14544 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 73 nsew signal input
flabel metal3 s 19200 14832 20000 14952 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 74 nsew signal input
flabel metal3 s 19200 15240 20000 15360 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 75 nsew signal input
flabel metal3 s 19200 15648 20000 15768 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 76 nsew signal input
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 77 nsew signal input
flabel metal3 s 19200 16464 20000 16584 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 78 nsew signal input
flabel metal3 s 19200 9120 20000 9240 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 79 nsew signal input
flabel metal3 s 19200 9528 20000 9648 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 80 nsew signal input
flabel metal3 s 19200 9936 20000 10056 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 81 nsew signal input
flabel metal3 s 19200 10344 20000 10464 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 82 nsew signal input
flabel metal3 s 19200 10752 20000 10872 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 83 nsew signal input
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 84 nsew signal input
flabel metal3 s 19200 11568 20000 11688 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 85 nsew signal input
flabel metal3 s 19200 11976 20000 12096 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 86 nsew signal input
flabel metal3 s 19200 12384 20000 12504 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 87 nsew signal input
flabel metal3 s 19200 552 20000 672 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 88 nsew signal tristate
flabel metal3 s 19200 4632 20000 4752 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 89 nsew signal tristate
flabel metal3 s 19200 5040 20000 5160 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 90 nsew signal tristate
flabel metal3 s 19200 5448 20000 5568 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 91 nsew signal tristate
flabel metal3 s 19200 5856 20000 5976 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 92 nsew signal tristate
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 93 nsew signal tristate
flabel metal3 s 19200 6672 20000 6792 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 94 nsew signal tristate
flabel metal3 s 19200 7080 20000 7200 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 95 nsew signal tristate
flabel metal3 s 19200 7488 20000 7608 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 96 nsew signal tristate
flabel metal3 s 19200 7896 20000 8016 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 97 nsew signal tristate
flabel metal3 s 19200 8304 20000 8424 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 98 nsew signal tristate
flabel metal3 s 19200 960 20000 1080 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 99 nsew signal tristate
flabel metal3 s 19200 1368 20000 1488 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 100 nsew signal tristate
flabel metal3 s 19200 1776 20000 1896 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 101 nsew signal tristate
flabel metal3 s 19200 2184 20000 2304 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 102 nsew signal tristate
flabel metal3 s 19200 2592 20000 2712 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 103 nsew signal tristate
flabel metal3 s 19200 3000 20000 3120 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 104 nsew signal tristate
flabel metal3 s 19200 3408 20000 3528 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 105 nsew signal tristate
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 106 nsew signal tristate
flabel metal3 s 19200 4224 20000 4344 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 107 nsew signal tristate
flabel metal2 s 14370 16400 14426 17200 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 108 nsew signal tristate
flabel metal2 s 16578 16400 16634 17200 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 109 nsew signal input
flabel metal2 s 18786 16400 18842 17200 0 FreeSans 224 90 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 110 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 prog_clk_0_S_in
port 111 nsew signal input
flabel metal3 s 0 280 800 400 0 FreeSans 480 0 0 0 prog_clk_0_W_out
port 112 nsew signal tristate
flabel metal2 s 12162 16400 12218 17200 0 FreeSans 224 90 0 0 top_grid_pin_0_
port 113 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
