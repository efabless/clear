VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_core
  CLASS BLOCK ;
  FOREIGN fpga_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2540.440 BY 2899.420 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 362.430 26.930 363.030 ;
    END
  END IO_ISOL_N
  PIN Test_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 165.230 26.930 165.830 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 2702.310 2517.930 2702.910 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 66.630 26.930 67.230 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 263.830 26.930 264.430 ;
    END
  END clk
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.020 2878.630 69.300 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 554.190 2517.930 554.790 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 911.870 2517.930 912.470 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 1270.230 2517.930 1270.830 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 1628.590 2517.930 1629.190 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 1986.270 2517.930 1986.870 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 2344.630 2517.930 2345.230 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2211.700 17.630 2211.980 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2223.200 17.630 2223.480 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2234.700 17.630 2234.980 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2246.200 17.630 2246.480 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.020 2878.630 161.300 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.700 17.630 2257.980 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2269.200 17.630 2269.480 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2280.700 17.630 2280.980 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.200 17.630 2292.480 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2303.700 17.630 2303.980 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.820 17.630 1900.100 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.320 17.630 1911.600 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.820 17.630 1923.100 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1934.320 17.630 1934.600 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.820 17.630 1946.100 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.480 2878.630 253.760 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.320 17.630 1957.600 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1968.820 17.630 1969.100 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.320 17.630 1980.600 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.820 17.630 1992.100 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.940 17.630 1588.220 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.440 17.630 1599.720 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.940 17.630 1611.220 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.440 17.630 1622.720 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.940 17.630 1634.220 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.440 17.630 1645.720 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.940 2878.630 346.220 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.940 17.630 1657.220 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.440 17.630 1668.720 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.940 17.630 1680.220 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.060 17.630 1276.340 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.560 17.630 1287.840 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.060 17.630 1299.340 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.560 17.630 1310.840 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.060 17.630 1322.340 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.560 17.630 1333.840 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.060 17.630 1345.340 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.400 2878.630 438.680 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.560 17.630 1356.840 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.060 17.630 1368.340 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.180 17.630 964.460 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.680 17.630 975.960 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.180 17.630 987.460 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.680 17.630 998.960 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.180 17.630 1010.460 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.680 17.630 1021.960 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.180 17.630 1033.460 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.680 17.630 1044.960 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.860 2878.630 531.140 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.180 17.630 1056.460 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.300 17.630 652.580 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.800 17.630 664.080 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.300 17.630 675.580 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.800 17.630 687.080 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.300 17.630 698.580 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.800 17.630 710.080 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.300 17.630 721.580 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.800 17.630 733.080 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.300 17.630 744.580 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.320 2878.630 623.600 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.420 17.630 340.700 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.920 17.630 352.200 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.420 17.630 363.700 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.920 17.630 375.200 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.420 17.630 386.700 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.920 17.630 398.200 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.420 17.630 409.700 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.920 17.630 421.200 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.420 17.630 432.700 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.540 17.630 28.820 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.780 2878.630 716.060 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.040 17.630 40.320 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.540 17.630 51.820 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.040 17.630 63.320 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.540 17.630 74.820 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.040 17.630 86.320 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.540 17.630 97.820 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.040 17.630 109.320 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.540 17.630 120.820 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 461.710 26.930 462.310 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 757.510 26.930 758.110 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.240 2878.630 808.520 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 1053.990 26.930 1054.590 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 1350.470 26.930 1351.070 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 1646.950 26.930 1647.550 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 1943.430 26.930 1944.030 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 2239.910 26.930 2240.510 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 2535.710 26.930 2536.310 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 195.830 2517.930 196.430 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.700 2878.630 900.980 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 673.190 2517.930 673.790 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 1031.550 2517.930 1032.150 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 1389.230 2517.930 1389.830 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 1747.590 2517.930 1748.190 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 2105.950 2517.930 2106.550 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 2463.630 2517.930 2464.230 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.660 17.630 2315.940 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2327.160 17.630 2327.440 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2338.660 17.630 2338.940 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.160 17.630 2350.440 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.700 2878.630 992.980 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.660 17.630 2361.940 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.160 17.630 2373.440 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.660 17.630 2384.940 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.160 17.630 2396.440 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2407.660 17.630 2407.940 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.780 17.630 2004.060 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2015.280 17.630 2015.560 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2026.780 17.630 2027.060 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.280 17.630 2038.560 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2049.780 17.630 2050.060 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.160 2878.630 1085.440 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2061.280 17.630 2061.560 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.780 17.630 2073.060 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.280 17.630 2084.560 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.780 17.630 2096.060 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.900 17.630 1692.180 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.400 17.630 1703.680 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.900 17.630 1715.180 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.400 17.630 1726.680 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.900 17.630 1738.180 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.400 17.630 1749.680 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.620 2878.630 1177.900 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.900 17.630 1761.180 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.400 17.630 1772.680 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.900 17.630 1784.180 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.020 17.630 1380.300 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.520 17.630 1391.800 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.020 17.630 1403.300 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.520 17.630 1414.800 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.020 17.630 1426.300 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.520 17.630 1437.800 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.020 17.630 1449.300 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1270.080 2878.630 1270.360 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.520 17.630 1460.800 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.020 17.630 1472.300 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.140 17.630 1068.420 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.640 17.630 1079.920 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.140 17.630 1091.420 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.640 17.630 1102.920 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.140 17.630 1114.420 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.640 17.630 1125.920 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.140 17.630 1137.420 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.640 17.630 1148.920 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.540 2878.630 1362.820 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.140 17.630 1160.420 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.260 17.630 756.540 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.760 17.630 768.040 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.260 17.630 779.540 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.760 17.630 791.040 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.260 17.630 802.540 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.760 17.630 814.040 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.260 17.630 825.540 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.760 17.630 837.040 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.260 17.630 848.540 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.000 2878.630 1455.280 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.380 17.630 444.660 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.880 17.630 456.160 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.380 17.630 467.660 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.880 17.630 479.160 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.380 17.630 490.660 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.880 17.630 502.160 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.380 17.630 513.660 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.880 17.630 525.160 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.380 17.630 536.660 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.500 17.630 132.780 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.460 2878.630 1547.740 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.000 17.630 144.280 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.500 17.630 155.780 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.000 17.630 167.280 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.500 17.630 178.780 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.000 17.630 190.280 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.500 17.630 201.780 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.000 17.630 213.280 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.500 17.630 224.780 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 560.310 26.930 560.910 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 856.790 26.930 857.390 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.920 2878.630 1640.200 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 1153.270 26.930 1153.870 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 1449.070 26.930 1449.670 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 1745.550 26.930 1746.150 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 2042.030 26.930 2042.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 2338.510 26.930 2339.110 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 2634.990 26.930 2635.590 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 315.510 2517.930 316.110 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.380 2878.630 1732.660 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 792.870 2517.930 793.470 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 1150.550 2517.930 1151.150 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 1508.910 2517.930 1509.510 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 1867.270 2517.930 1867.870 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 2224.950 2517.930 2225.550 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 2583.310 2517.930 2583.910 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2419.620 17.630 2419.900 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.120 17.630 2431.400 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2442.620 17.630 2442.900 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2454.120 17.630 2454.400 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.380 2878.630 1824.660 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2465.620 17.630 2465.900 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2477.120 17.630 2477.400 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2488.620 17.630 2488.900 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.120 17.630 2500.400 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2511.620 17.630 2511.900 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.740 17.630 2108.020 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.240 17.630 2119.520 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.740 17.630 2131.020 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.240 17.630 2142.520 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2153.740 17.630 2154.020 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1916.840 2878.630 1917.120 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2165.240 17.630 2165.520 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.740 17.630 2177.020 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2188.240 17.630 2188.520 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.740 17.630 2200.020 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.860 17.630 1796.140 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1807.360 17.630 1807.640 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.860 17.630 1819.140 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.360 17.630 1830.640 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.860 17.630 1842.140 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.360 17.630 1853.640 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.300 2878.630 2009.580 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.860 17.630 1865.140 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.360 17.630 1876.640 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.860 17.630 1888.140 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.980 17.630 1484.260 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.480 17.630 1495.760 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.980 17.630 1507.260 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.480 17.630 1518.760 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.980 17.630 1530.260 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.480 17.630 1541.760 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.980 17.630 1553.260 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.760 2878.630 2102.040 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.480 17.630 1564.760 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.980 17.630 1576.260 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.100 17.630 1172.380 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.600 17.630 1183.880 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.100 17.630 1195.380 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.600 17.630 1206.880 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.100 17.630 1218.380 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.600 17.630 1229.880 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.100 17.630 1241.380 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.600 17.630 1252.880 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.220 2878.630 2194.500 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.100 17.630 1264.380 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.220 17.630 860.500 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.720 17.630 872.000 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.220 17.630 883.500 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.720 17.630 895.000 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.220 17.630 906.500 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.720 17.630 918.000 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.220 17.630 929.500 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.720 17.630 941.000 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.220 17.630 952.500 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.680 2878.630 2286.960 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.340 17.630 548.620 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.840 17.630 560.120 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.340 17.630 571.620 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.840 17.630 583.120 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.340 17.630 594.620 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.840 17.630 606.120 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.340 17.630 617.620 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.840 17.630 629.120 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.340 17.630 640.620 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.460 17.630 236.740 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2379.140 2878.630 2379.420 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.960 17.630 248.240 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.460 17.630 259.740 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.960 17.630 271.240 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.460 17.630 282.740 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.960 17.630 294.240 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.460 17.630 305.740 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.960 17.630 317.240 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.460 17.630 328.740 21.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 658.910 26.930 659.510 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 955.390 26.930 955.990 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2471.600 2878.630 2471.880 2882.630 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 1251.870 26.930 1252.470 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 1548.350 26.930 1548.950 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 1844.150 26.930 1844.750 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 2140.630 26.930 2141.230 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 2437.110 26.930 2437.710 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 2733.590 26.930 2734.190 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 434.510 2517.930 435.110 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 76.830 2517.930 77.430 ;
    END
  END prog_clk
  PIN sc_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.930 2832.190 26.930 2832.790 ;
    END
  END sc_head
  PIN sc_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2513.930 2821.990 2517.930 2822.590 ;
    END
  END sc_tail
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2529.740 6.260 2534.240 2893.160 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 6.200 6.260 10.700 2893.160 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 6.200 2888.660 2534.240 2893.160 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2861.260 2540.440 2865.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2816.260 2540.440 2820.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2771.260 2540.440 2775.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2726.260 2540.440 2730.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2681.260 2540.440 2685.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2636.260 2540.440 2640.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2591.260 2540.440 2595.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2546.260 2540.440 2550.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2501.260 2540.440 2505.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2456.260 2540.440 2460.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2411.260 2540.440 2415.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2366.260 2540.440 2370.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2321.260 2540.440 2325.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2276.260 2540.440 2280.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2231.260 2540.440 2235.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2186.260 2540.440 2190.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2141.260 2540.440 2145.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2096.260 2540.440 2100.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2051.260 2540.440 2055.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2006.260 2540.440 2010.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1961.260 2540.440 1965.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1916.260 2540.440 1920.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1871.260 2540.440 1875.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1826.260 2540.440 1830.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1781.260 2540.440 1785.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1736.260 2540.440 1740.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1691.260 2540.440 1695.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1646.260 2540.440 1650.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1601.260 2540.440 1605.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1556.260 2540.440 1560.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1511.260 2540.440 1515.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1466.260 2540.440 1470.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1421.260 2540.440 1425.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1376.260 2540.440 1380.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1331.260 2540.440 1335.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1286.260 2540.440 1290.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1241.260 2540.440 1245.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1196.260 2540.440 1200.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1151.260 2540.440 1155.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1106.260 2540.440 1110.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1061.260 2540.440 1065.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 1016.260 2540.440 1020.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 971.260 2540.440 975.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 926.260 2540.440 930.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 881.260 2540.440 885.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 836.260 2540.440 840.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 791.260 2540.440 795.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 746.260 2540.440 750.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 701.260 2540.440 705.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 656.260 2540.440 660.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 611.260 2540.440 615.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 566.260 2540.440 570.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 521.260 2540.440 525.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 476.260 2540.440 480.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 431.260 2540.440 435.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 386.260 2540.440 390.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 341.260 2540.440 345.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 296.260 2540.440 300.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 251.260 2540.440 255.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 206.260 2540.440 210.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 161.260 2540.440 165.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 116.260 2540.440 120.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 6.200 6.260 2534.240 10.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2535.940 0.060 2540.440 2899.360 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.060 4.500 2899.360 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2894.860 2540.440 2899.360 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2838.760 2540.440 2843.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2793.760 2540.440 2798.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2748.760 2540.440 2753.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2703.760 2540.440 2708.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2658.760 2540.440 2663.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2613.760 2540.440 2618.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2568.760 2540.440 2573.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2523.760 2540.440 2528.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2478.760 2540.440 2483.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2433.760 2540.440 2438.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2388.760 2540.440 2393.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2343.760 2540.440 2348.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2298.760 2540.440 2303.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2253.760 2540.440 2258.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2208.760 2540.440 2213.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2163.760 2540.440 2168.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2118.760 2540.440 2123.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2073.760 2540.440 2078.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 2028.760 2540.440 2033.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1983.760 2540.440 1988.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1938.760 2540.440 1943.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1893.760 2540.440 1898.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1848.760 2540.440 1853.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1803.760 2540.440 1808.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1758.760 2540.440 1763.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1713.760 2540.440 1718.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1668.760 2540.440 1673.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1623.760 2540.440 1628.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1578.760 2540.440 1583.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1533.760 2540.440 1538.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1488.760 2540.440 1493.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1443.760 2540.440 1448.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1398.760 2540.440 1403.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1353.760 2540.440 1358.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1308.760 2540.440 1313.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1263.760 2540.440 1268.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1218.760 2540.440 1223.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1173.760 2540.440 1178.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1128.760 2540.440 1133.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1083.760 2540.440 1088.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 1038.760 2540.440 1043.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 993.760 2540.440 998.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 948.760 2540.440 953.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 903.760 2540.440 908.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 858.760 2540.440 863.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 813.760 2540.440 818.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 768.760 2540.440 773.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 723.760 2540.440 728.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 678.760 2540.440 683.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 633.760 2540.440 638.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 588.760 2540.440 593.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 543.760 2540.440 548.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 498.760 2540.440 503.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 453.760 2540.440 458.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 408.760 2540.440 413.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 363.760 2540.440 368.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 318.760 2540.440 323.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 273.760 2540.440 278.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 228.760 2540.440 233.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 183.760 2540.440 188.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 138.760 2540.440 143.260 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.060 2540.440 4.560 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 78.450 33.355 2462.410 2867.835 ;
      LAYER met1 ;
        RECT 28.520 31.950 2511.920 2867.990 ;
      LAYER met2 ;
        RECT 28.550 2878.350 68.740 2878.630 ;
        RECT 69.580 2878.350 160.740 2878.630 ;
        RECT 161.580 2878.350 253.200 2878.630 ;
        RECT 254.040 2878.350 345.660 2878.630 ;
        RECT 346.500 2878.350 438.120 2878.630 ;
        RECT 438.960 2878.350 530.580 2878.630 ;
        RECT 531.420 2878.350 623.040 2878.630 ;
        RECT 623.880 2878.350 715.500 2878.630 ;
        RECT 716.340 2878.350 807.960 2878.630 ;
        RECT 808.800 2878.350 900.420 2878.630 ;
        RECT 901.260 2878.350 992.420 2878.630 ;
        RECT 993.260 2878.350 1084.880 2878.630 ;
        RECT 1085.720 2878.350 1177.340 2878.630 ;
        RECT 1178.180 2878.350 1269.800 2878.630 ;
        RECT 1270.640 2878.350 1362.260 2878.630 ;
        RECT 1363.100 2878.350 1454.720 2878.630 ;
        RECT 1455.560 2878.350 1547.180 2878.630 ;
        RECT 1548.020 2878.350 1639.640 2878.630 ;
        RECT 1640.480 2878.350 1732.100 2878.630 ;
        RECT 1732.940 2878.350 1824.100 2878.630 ;
        RECT 1824.940 2878.350 1916.560 2878.630 ;
        RECT 1917.400 2878.350 2009.020 2878.630 ;
        RECT 2009.860 2878.350 2101.480 2878.630 ;
        RECT 2102.320 2878.350 2193.940 2878.630 ;
        RECT 2194.780 2878.350 2286.400 2878.630 ;
        RECT 2287.240 2878.350 2378.860 2878.630 ;
        RECT 2379.700 2878.350 2471.320 2878.630 ;
        RECT 2472.160 2878.350 2511.890 2878.630 ;
        RECT 28.550 21.910 2511.890 2878.350 ;
        RECT 29.100 21.630 39.760 21.910 ;
        RECT 40.600 21.630 51.260 21.910 ;
        RECT 52.100 21.630 62.760 21.910 ;
        RECT 63.600 21.630 74.260 21.910 ;
        RECT 75.100 21.630 85.760 21.910 ;
        RECT 86.600 21.630 97.260 21.910 ;
        RECT 98.100 21.630 108.760 21.910 ;
        RECT 109.600 21.630 120.260 21.910 ;
        RECT 121.100 21.630 132.220 21.910 ;
        RECT 133.060 21.630 143.720 21.910 ;
        RECT 144.560 21.630 155.220 21.910 ;
        RECT 156.060 21.630 166.720 21.910 ;
        RECT 167.560 21.630 178.220 21.910 ;
        RECT 179.060 21.630 189.720 21.910 ;
        RECT 190.560 21.630 201.220 21.910 ;
        RECT 202.060 21.630 212.720 21.910 ;
        RECT 213.560 21.630 224.220 21.910 ;
        RECT 225.060 21.630 236.180 21.910 ;
        RECT 237.020 21.630 247.680 21.910 ;
        RECT 248.520 21.630 259.180 21.910 ;
        RECT 260.020 21.630 270.680 21.910 ;
        RECT 271.520 21.630 282.180 21.910 ;
        RECT 283.020 21.630 293.680 21.910 ;
        RECT 294.520 21.630 305.180 21.910 ;
        RECT 306.020 21.630 316.680 21.910 ;
        RECT 317.520 21.630 328.180 21.910 ;
        RECT 329.020 21.630 340.140 21.910 ;
        RECT 340.980 21.630 351.640 21.910 ;
        RECT 352.480 21.630 363.140 21.910 ;
        RECT 363.980 21.630 374.640 21.910 ;
        RECT 375.480 21.630 386.140 21.910 ;
        RECT 386.980 21.630 397.640 21.910 ;
        RECT 398.480 21.630 409.140 21.910 ;
        RECT 409.980 21.630 420.640 21.910 ;
        RECT 421.480 21.630 432.140 21.910 ;
        RECT 432.980 21.630 444.100 21.910 ;
        RECT 444.940 21.630 455.600 21.910 ;
        RECT 456.440 21.630 467.100 21.910 ;
        RECT 467.940 21.630 478.600 21.910 ;
        RECT 479.440 21.630 490.100 21.910 ;
        RECT 490.940 21.630 501.600 21.910 ;
        RECT 502.440 21.630 513.100 21.910 ;
        RECT 513.940 21.630 524.600 21.910 ;
        RECT 525.440 21.630 536.100 21.910 ;
        RECT 536.940 21.630 548.060 21.910 ;
        RECT 548.900 21.630 559.560 21.910 ;
        RECT 560.400 21.630 571.060 21.910 ;
        RECT 571.900 21.630 582.560 21.910 ;
        RECT 583.400 21.630 594.060 21.910 ;
        RECT 594.900 21.630 605.560 21.910 ;
        RECT 606.400 21.630 617.060 21.910 ;
        RECT 617.900 21.630 628.560 21.910 ;
        RECT 629.400 21.630 640.060 21.910 ;
        RECT 640.900 21.630 652.020 21.910 ;
        RECT 652.860 21.630 663.520 21.910 ;
        RECT 664.360 21.630 675.020 21.910 ;
        RECT 675.860 21.630 686.520 21.910 ;
        RECT 687.360 21.630 698.020 21.910 ;
        RECT 698.860 21.630 709.520 21.910 ;
        RECT 710.360 21.630 721.020 21.910 ;
        RECT 721.860 21.630 732.520 21.910 ;
        RECT 733.360 21.630 744.020 21.910 ;
        RECT 744.860 21.630 755.980 21.910 ;
        RECT 756.820 21.630 767.480 21.910 ;
        RECT 768.320 21.630 778.980 21.910 ;
        RECT 779.820 21.630 790.480 21.910 ;
        RECT 791.320 21.630 801.980 21.910 ;
        RECT 802.820 21.630 813.480 21.910 ;
        RECT 814.320 21.630 824.980 21.910 ;
        RECT 825.820 21.630 836.480 21.910 ;
        RECT 837.320 21.630 847.980 21.910 ;
        RECT 848.820 21.630 859.940 21.910 ;
        RECT 860.780 21.630 871.440 21.910 ;
        RECT 872.280 21.630 882.940 21.910 ;
        RECT 883.780 21.630 894.440 21.910 ;
        RECT 895.280 21.630 905.940 21.910 ;
        RECT 906.780 21.630 917.440 21.910 ;
        RECT 918.280 21.630 928.940 21.910 ;
        RECT 929.780 21.630 940.440 21.910 ;
        RECT 941.280 21.630 951.940 21.910 ;
        RECT 952.780 21.630 963.900 21.910 ;
        RECT 964.740 21.630 975.400 21.910 ;
        RECT 976.240 21.630 986.900 21.910 ;
        RECT 987.740 21.630 998.400 21.910 ;
        RECT 999.240 21.630 1009.900 21.910 ;
        RECT 1010.740 21.630 1021.400 21.910 ;
        RECT 1022.240 21.630 1032.900 21.910 ;
        RECT 1033.740 21.630 1044.400 21.910 ;
        RECT 1045.240 21.630 1055.900 21.910 ;
        RECT 1056.740 21.630 1067.860 21.910 ;
        RECT 1068.700 21.630 1079.360 21.910 ;
        RECT 1080.200 21.630 1090.860 21.910 ;
        RECT 1091.700 21.630 1102.360 21.910 ;
        RECT 1103.200 21.630 1113.860 21.910 ;
        RECT 1114.700 21.630 1125.360 21.910 ;
        RECT 1126.200 21.630 1136.860 21.910 ;
        RECT 1137.700 21.630 1148.360 21.910 ;
        RECT 1149.200 21.630 1159.860 21.910 ;
        RECT 1160.700 21.630 1171.820 21.910 ;
        RECT 1172.660 21.630 1183.320 21.910 ;
        RECT 1184.160 21.630 1194.820 21.910 ;
        RECT 1195.660 21.630 1206.320 21.910 ;
        RECT 1207.160 21.630 1217.820 21.910 ;
        RECT 1218.660 21.630 1229.320 21.910 ;
        RECT 1230.160 21.630 1240.820 21.910 ;
        RECT 1241.660 21.630 1252.320 21.910 ;
        RECT 1253.160 21.630 1263.820 21.910 ;
        RECT 1264.660 21.630 1275.780 21.910 ;
        RECT 1276.620 21.630 1287.280 21.910 ;
        RECT 1288.120 21.630 1298.780 21.910 ;
        RECT 1299.620 21.630 1310.280 21.910 ;
        RECT 1311.120 21.630 1321.780 21.910 ;
        RECT 1322.620 21.630 1333.280 21.910 ;
        RECT 1334.120 21.630 1344.780 21.910 ;
        RECT 1345.620 21.630 1356.280 21.910 ;
        RECT 1357.120 21.630 1367.780 21.910 ;
        RECT 1368.620 21.630 1379.740 21.910 ;
        RECT 1380.580 21.630 1391.240 21.910 ;
        RECT 1392.080 21.630 1402.740 21.910 ;
        RECT 1403.580 21.630 1414.240 21.910 ;
        RECT 1415.080 21.630 1425.740 21.910 ;
        RECT 1426.580 21.630 1437.240 21.910 ;
        RECT 1438.080 21.630 1448.740 21.910 ;
        RECT 1449.580 21.630 1460.240 21.910 ;
        RECT 1461.080 21.630 1471.740 21.910 ;
        RECT 1472.580 21.630 1483.700 21.910 ;
        RECT 1484.540 21.630 1495.200 21.910 ;
        RECT 1496.040 21.630 1506.700 21.910 ;
        RECT 1507.540 21.630 1518.200 21.910 ;
        RECT 1519.040 21.630 1529.700 21.910 ;
        RECT 1530.540 21.630 1541.200 21.910 ;
        RECT 1542.040 21.630 1552.700 21.910 ;
        RECT 1553.540 21.630 1564.200 21.910 ;
        RECT 1565.040 21.630 1575.700 21.910 ;
        RECT 1576.540 21.630 1587.660 21.910 ;
        RECT 1588.500 21.630 1599.160 21.910 ;
        RECT 1600.000 21.630 1610.660 21.910 ;
        RECT 1611.500 21.630 1622.160 21.910 ;
        RECT 1623.000 21.630 1633.660 21.910 ;
        RECT 1634.500 21.630 1645.160 21.910 ;
        RECT 1646.000 21.630 1656.660 21.910 ;
        RECT 1657.500 21.630 1668.160 21.910 ;
        RECT 1669.000 21.630 1679.660 21.910 ;
        RECT 1680.500 21.630 1691.620 21.910 ;
        RECT 1692.460 21.630 1703.120 21.910 ;
        RECT 1703.960 21.630 1714.620 21.910 ;
        RECT 1715.460 21.630 1726.120 21.910 ;
        RECT 1726.960 21.630 1737.620 21.910 ;
        RECT 1738.460 21.630 1749.120 21.910 ;
        RECT 1749.960 21.630 1760.620 21.910 ;
        RECT 1761.460 21.630 1772.120 21.910 ;
        RECT 1772.960 21.630 1783.620 21.910 ;
        RECT 1784.460 21.630 1795.580 21.910 ;
        RECT 1796.420 21.630 1807.080 21.910 ;
        RECT 1807.920 21.630 1818.580 21.910 ;
        RECT 1819.420 21.630 1830.080 21.910 ;
        RECT 1830.920 21.630 1841.580 21.910 ;
        RECT 1842.420 21.630 1853.080 21.910 ;
        RECT 1853.920 21.630 1864.580 21.910 ;
        RECT 1865.420 21.630 1876.080 21.910 ;
        RECT 1876.920 21.630 1887.580 21.910 ;
        RECT 1888.420 21.630 1899.540 21.910 ;
        RECT 1900.380 21.630 1911.040 21.910 ;
        RECT 1911.880 21.630 1922.540 21.910 ;
        RECT 1923.380 21.630 1934.040 21.910 ;
        RECT 1934.880 21.630 1945.540 21.910 ;
        RECT 1946.380 21.630 1957.040 21.910 ;
        RECT 1957.880 21.630 1968.540 21.910 ;
        RECT 1969.380 21.630 1980.040 21.910 ;
        RECT 1980.880 21.630 1991.540 21.910 ;
        RECT 1992.380 21.630 2003.500 21.910 ;
        RECT 2004.340 21.630 2015.000 21.910 ;
        RECT 2015.840 21.630 2026.500 21.910 ;
        RECT 2027.340 21.630 2038.000 21.910 ;
        RECT 2038.840 21.630 2049.500 21.910 ;
        RECT 2050.340 21.630 2061.000 21.910 ;
        RECT 2061.840 21.630 2072.500 21.910 ;
        RECT 2073.340 21.630 2084.000 21.910 ;
        RECT 2084.840 21.630 2095.500 21.910 ;
        RECT 2096.340 21.630 2107.460 21.910 ;
        RECT 2108.300 21.630 2118.960 21.910 ;
        RECT 2119.800 21.630 2130.460 21.910 ;
        RECT 2131.300 21.630 2141.960 21.910 ;
        RECT 2142.800 21.630 2153.460 21.910 ;
        RECT 2154.300 21.630 2164.960 21.910 ;
        RECT 2165.800 21.630 2176.460 21.910 ;
        RECT 2177.300 21.630 2187.960 21.910 ;
        RECT 2188.800 21.630 2199.460 21.910 ;
        RECT 2200.300 21.630 2211.420 21.910 ;
        RECT 2212.260 21.630 2222.920 21.910 ;
        RECT 2223.760 21.630 2234.420 21.910 ;
        RECT 2235.260 21.630 2245.920 21.910 ;
        RECT 2246.760 21.630 2257.420 21.910 ;
        RECT 2258.260 21.630 2268.920 21.910 ;
        RECT 2269.760 21.630 2280.420 21.910 ;
        RECT 2281.260 21.630 2291.920 21.910 ;
        RECT 2292.760 21.630 2303.420 21.910 ;
        RECT 2304.260 21.630 2315.380 21.910 ;
        RECT 2316.220 21.630 2326.880 21.910 ;
        RECT 2327.720 21.630 2338.380 21.910 ;
        RECT 2339.220 21.630 2349.880 21.910 ;
        RECT 2350.720 21.630 2361.380 21.910 ;
        RECT 2362.220 21.630 2372.880 21.910 ;
        RECT 2373.720 21.630 2384.380 21.910 ;
        RECT 2385.220 21.630 2395.880 21.910 ;
        RECT 2396.720 21.630 2407.380 21.910 ;
        RECT 2408.220 21.630 2419.340 21.910 ;
        RECT 2420.180 21.630 2430.840 21.910 ;
        RECT 2431.680 21.630 2442.340 21.910 ;
        RECT 2443.180 21.630 2453.840 21.910 ;
        RECT 2454.680 21.630 2465.340 21.910 ;
        RECT 2466.180 21.630 2476.840 21.910 ;
        RECT 2477.680 21.630 2488.340 21.910 ;
        RECT 2489.180 21.630 2499.840 21.910 ;
        RECT 2500.680 21.630 2511.340 21.910 ;
      LAYER met3 ;
        RECT 26.930 2833.190 2513.930 2867.915 ;
        RECT 27.330 2831.790 2513.930 2833.190 ;
        RECT 26.930 2822.990 2513.930 2831.790 ;
        RECT 26.930 2821.590 2513.530 2822.990 ;
        RECT 26.930 2734.590 2513.930 2821.590 ;
        RECT 27.330 2733.190 2513.930 2734.590 ;
        RECT 26.930 2703.310 2513.930 2733.190 ;
        RECT 26.930 2701.910 2513.530 2703.310 ;
        RECT 26.930 2635.990 2513.930 2701.910 ;
        RECT 27.330 2634.590 2513.930 2635.990 ;
        RECT 26.930 2584.310 2513.930 2634.590 ;
        RECT 26.930 2582.910 2513.530 2584.310 ;
        RECT 26.930 2536.710 2513.930 2582.910 ;
        RECT 27.330 2535.310 2513.930 2536.710 ;
        RECT 26.930 2464.630 2513.930 2535.310 ;
        RECT 26.930 2463.230 2513.530 2464.630 ;
        RECT 26.930 2438.110 2513.930 2463.230 ;
        RECT 27.330 2436.710 2513.930 2438.110 ;
        RECT 26.930 2345.630 2513.930 2436.710 ;
        RECT 26.930 2344.230 2513.530 2345.630 ;
        RECT 26.930 2339.510 2513.930 2344.230 ;
        RECT 27.330 2338.110 2513.930 2339.510 ;
        RECT 26.930 2240.910 2513.930 2338.110 ;
        RECT 27.330 2239.510 2513.930 2240.910 ;
        RECT 26.930 2225.950 2513.930 2239.510 ;
        RECT 26.930 2224.550 2513.530 2225.950 ;
        RECT 26.930 2141.630 2513.930 2224.550 ;
        RECT 27.330 2140.230 2513.930 2141.630 ;
        RECT 26.930 2106.950 2513.930 2140.230 ;
        RECT 26.930 2105.550 2513.530 2106.950 ;
        RECT 26.930 2043.030 2513.930 2105.550 ;
        RECT 27.330 2041.630 2513.930 2043.030 ;
        RECT 26.930 1987.270 2513.930 2041.630 ;
        RECT 26.930 1985.870 2513.530 1987.270 ;
        RECT 26.930 1944.430 2513.930 1985.870 ;
        RECT 27.330 1943.030 2513.930 1944.430 ;
        RECT 26.930 1868.270 2513.930 1943.030 ;
        RECT 26.930 1866.870 2513.530 1868.270 ;
        RECT 26.930 1845.150 2513.930 1866.870 ;
        RECT 27.330 1843.750 2513.930 1845.150 ;
        RECT 26.930 1748.590 2513.930 1843.750 ;
        RECT 26.930 1747.190 2513.530 1748.590 ;
        RECT 26.930 1746.550 2513.930 1747.190 ;
        RECT 27.330 1745.150 2513.930 1746.550 ;
        RECT 26.930 1647.950 2513.930 1745.150 ;
        RECT 27.330 1646.550 2513.930 1647.950 ;
        RECT 26.930 1629.590 2513.930 1646.550 ;
        RECT 26.930 1628.190 2513.530 1629.590 ;
        RECT 26.930 1549.350 2513.930 1628.190 ;
        RECT 27.330 1547.950 2513.930 1549.350 ;
        RECT 26.930 1509.910 2513.930 1547.950 ;
        RECT 26.930 1508.510 2513.530 1509.910 ;
        RECT 26.930 1450.070 2513.930 1508.510 ;
        RECT 27.330 1448.670 2513.930 1450.070 ;
        RECT 26.930 1390.230 2513.930 1448.670 ;
        RECT 26.930 1388.830 2513.530 1390.230 ;
        RECT 26.930 1351.470 2513.930 1388.830 ;
        RECT 27.330 1350.070 2513.930 1351.470 ;
        RECT 26.930 1271.230 2513.930 1350.070 ;
        RECT 26.930 1269.830 2513.530 1271.230 ;
        RECT 26.930 1252.870 2513.930 1269.830 ;
        RECT 27.330 1251.470 2513.930 1252.870 ;
        RECT 26.930 1154.270 2513.930 1251.470 ;
        RECT 27.330 1152.870 2513.930 1154.270 ;
        RECT 26.930 1151.550 2513.930 1152.870 ;
        RECT 26.930 1150.150 2513.530 1151.550 ;
        RECT 26.930 1054.990 2513.930 1150.150 ;
        RECT 27.330 1053.590 2513.930 1054.990 ;
        RECT 26.930 1032.550 2513.930 1053.590 ;
        RECT 26.930 1031.150 2513.530 1032.550 ;
        RECT 26.930 956.390 2513.930 1031.150 ;
        RECT 27.330 954.990 2513.930 956.390 ;
        RECT 26.930 912.870 2513.930 954.990 ;
        RECT 26.930 911.470 2513.530 912.870 ;
        RECT 26.930 857.790 2513.930 911.470 ;
        RECT 27.330 856.390 2513.930 857.790 ;
        RECT 26.930 793.870 2513.930 856.390 ;
        RECT 26.930 792.470 2513.530 793.870 ;
        RECT 26.930 758.510 2513.930 792.470 ;
        RECT 27.330 757.110 2513.930 758.510 ;
        RECT 26.930 674.190 2513.930 757.110 ;
        RECT 26.930 672.790 2513.530 674.190 ;
        RECT 26.930 659.910 2513.930 672.790 ;
        RECT 27.330 658.510 2513.930 659.910 ;
        RECT 26.930 561.310 2513.930 658.510 ;
        RECT 27.330 559.910 2513.930 561.310 ;
        RECT 26.930 555.190 2513.930 559.910 ;
        RECT 26.930 553.790 2513.530 555.190 ;
        RECT 26.930 462.710 2513.930 553.790 ;
        RECT 27.330 461.310 2513.930 462.710 ;
        RECT 26.930 435.510 2513.930 461.310 ;
        RECT 26.930 434.110 2513.530 435.510 ;
        RECT 26.930 363.430 2513.930 434.110 ;
        RECT 27.330 362.030 2513.930 363.430 ;
        RECT 26.930 316.510 2513.930 362.030 ;
        RECT 26.930 315.110 2513.530 316.510 ;
        RECT 26.930 264.830 2513.930 315.110 ;
        RECT 27.330 263.430 2513.930 264.830 ;
        RECT 26.930 196.830 2513.930 263.430 ;
        RECT 26.930 195.430 2513.530 196.830 ;
        RECT 26.930 166.230 2513.930 195.430 ;
        RECT 27.330 164.830 2513.930 166.230 ;
        RECT 26.930 77.830 2513.930 164.830 ;
        RECT 26.930 76.430 2513.530 77.830 ;
        RECT 26.930 67.630 2513.930 76.430 ;
        RECT 27.330 66.765 2513.930 67.630 ;
      LAYER met4 ;
        RECT 84.865 98.725 2465.235 2867.990 ;
      LAYER met5 ;
        RECT 0.000 2899.360 4.500 2899.420 ;
        RECT 0.000 2894.800 4.500 2894.860 ;
        RECT 0.000 2887.060 4.600 2893.260 ;
        RECT 2535.840 2887.060 2540.440 2893.260 ;
        RECT 0.000 2867.360 2540.440 2887.060 ;
        RECT 0.000 2844.860 2540.440 2859.660 ;
        RECT 0.000 2843.260 4.500 2843.320 ;
        RECT 0.000 2838.700 4.500 2838.760 ;
        RECT 0.000 2822.360 2540.440 2837.160 ;
        RECT 0.000 2799.860 2540.440 2814.660 ;
        RECT 0.000 2798.260 4.500 2798.320 ;
        RECT 0.000 2793.700 4.500 2793.760 ;
        RECT 0.000 2777.360 2540.440 2792.160 ;
        RECT 0.000 2754.860 2540.440 2769.660 ;
        RECT 0.000 2753.260 4.500 2753.320 ;
        RECT 0.000 2748.700 4.500 2748.760 ;
        RECT 0.000 2732.360 2540.440 2747.160 ;
        RECT 0.000 2709.860 2540.440 2724.660 ;
        RECT 0.000 2708.260 4.500 2708.320 ;
        RECT 0.000 2703.700 4.500 2703.760 ;
        RECT 0.000 2687.360 2540.440 2702.160 ;
        RECT 0.000 2664.860 2540.440 2679.660 ;
        RECT 0.000 2663.260 4.500 2663.320 ;
        RECT 0.000 2658.700 4.500 2658.760 ;
        RECT 0.000 2642.360 2540.440 2657.160 ;
        RECT 0.000 2619.860 2540.440 2634.660 ;
        RECT 0.000 2618.260 4.500 2618.320 ;
        RECT 0.000 2613.700 4.500 2613.760 ;
        RECT 0.000 2597.360 2540.440 2612.160 ;
        RECT 0.000 2574.860 2540.440 2589.660 ;
        RECT 0.000 2573.260 4.500 2573.320 ;
        RECT 0.000 2568.700 4.500 2568.760 ;
        RECT 0.000 2552.360 2540.440 2567.160 ;
        RECT 0.000 2529.860 2540.440 2544.660 ;
        RECT 0.000 2528.260 4.500 2528.320 ;
        RECT 0.000 2523.700 4.500 2523.760 ;
        RECT 0.000 2507.360 2540.440 2522.160 ;
        RECT 0.000 2484.860 2540.440 2499.660 ;
        RECT 0.000 2483.260 4.500 2483.320 ;
        RECT 0.000 2478.700 4.500 2478.760 ;
        RECT 0.000 2462.360 2540.440 2477.160 ;
        RECT 0.000 2439.860 2540.440 2454.660 ;
        RECT 0.000 2438.260 4.500 2438.320 ;
        RECT 0.000 2433.700 4.500 2433.760 ;
        RECT 0.000 2417.360 2540.440 2432.160 ;
        RECT 0.000 2394.860 2540.440 2409.660 ;
        RECT 0.000 2393.260 4.500 2393.320 ;
        RECT 0.000 2388.700 4.500 2388.760 ;
        RECT 0.000 2372.360 2540.440 2387.160 ;
        RECT 0.000 2349.860 2540.440 2364.660 ;
        RECT 0.000 2348.260 4.500 2348.320 ;
        RECT 0.000 2343.700 4.500 2343.760 ;
        RECT 0.000 2327.360 2540.440 2342.160 ;
        RECT 0.000 2304.860 2540.440 2319.660 ;
        RECT 0.000 2303.260 4.500 2303.320 ;
        RECT 0.000 2298.700 4.500 2298.760 ;
        RECT 0.000 2282.360 2540.440 2297.160 ;
        RECT 0.000 2259.860 2540.440 2274.660 ;
        RECT 0.000 2258.260 4.500 2258.320 ;
        RECT 0.000 2253.700 4.500 2253.760 ;
        RECT 0.000 2237.360 2540.440 2252.160 ;
        RECT 0.000 2214.860 2540.440 2229.660 ;
        RECT 0.000 2213.260 4.500 2213.320 ;
        RECT 0.000 2208.700 4.500 2208.760 ;
        RECT 0.000 2192.360 2540.440 2207.160 ;
        RECT 0.000 2169.860 2540.440 2184.660 ;
        RECT 0.000 2168.260 4.500 2168.320 ;
        RECT 0.000 2163.700 4.500 2163.760 ;
        RECT 0.000 2147.360 2540.440 2162.160 ;
        RECT 0.000 2124.860 2540.440 2139.660 ;
        RECT 0.000 2123.260 4.500 2123.320 ;
        RECT 0.000 2118.700 4.500 2118.760 ;
        RECT 0.000 2102.360 2540.440 2117.160 ;
        RECT 0.000 2079.860 2540.440 2094.660 ;
        RECT 0.000 2078.260 4.500 2078.320 ;
        RECT 0.000 2073.700 4.500 2073.760 ;
        RECT 0.000 2057.360 2540.440 2072.160 ;
        RECT 0.000 2034.860 2540.440 2049.660 ;
        RECT 0.000 2033.260 4.500 2033.320 ;
        RECT 0.000 2028.700 4.500 2028.760 ;
        RECT 0.000 2012.360 2540.440 2027.160 ;
        RECT 0.000 1989.860 2540.440 2004.660 ;
        RECT 0.000 1988.260 4.500 1988.320 ;
        RECT 0.000 1983.700 4.500 1983.760 ;
        RECT 0.000 1967.360 2540.440 1982.160 ;
        RECT 0.000 1944.860 2540.440 1959.660 ;
        RECT 0.000 1943.260 4.500 1943.320 ;
        RECT 0.000 1938.700 4.500 1938.760 ;
        RECT 0.000 1922.360 2540.440 1937.160 ;
        RECT 0.000 1899.860 2540.440 1914.660 ;
        RECT 0.000 1898.260 4.500 1898.320 ;
        RECT 0.000 1893.700 4.500 1893.760 ;
        RECT 0.000 1877.360 2540.440 1892.160 ;
        RECT 0.000 1854.860 2540.440 1869.660 ;
        RECT 0.000 1853.260 4.500 1853.320 ;
        RECT 0.000 1848.700 4.500 1848.760 ;
        RECT 0.000 1832.360 2540.440 1847.160 ;
        RECT 0.000 1809.860 2540.440 1824.660 ;
        RECT 0.000 1808.260 4.500 1808.320 ;
        RECT 0.000 1803.700 4.500 1803.760 ;
        RECT 0.000 1787.360 2540.440 1802.160 ;
        RECT 0.000 1764.860 2540.440 1779.660 ;
        RECT 0.000 1763.260 4.500 1763.320 ;
        RECT 0.000 1758.700 4.500 1758.760 ;
        RECT 0.000 1742.360 2540.440 1757.160 ;
        RECT 0.000 1719.860 2540.440 1734.660 ;
        RECT 0.000 1718.260 4.500 1718.320 ;
        RECT 0.000 1713.700 4.500 1713.760 ;
        RECT 0.000 1697.360 2540.440 1712.160 ;
        RECT 0.000 1674.860 2540.440 1689.660 ;
        RECT 0.000 1673.260 4.500 1673.320 ;
        RECT 0.000 1668.700 4.500 1668.760 ;
        RECT 0.000 1652.360 2540.440 1667.160 ;
        RECT 0.000 1629.860 2540.440 1644.660 ;
        RECT 0.000 1628.260 4.500 1628.320 ;
        RECT 0.000 1623.700 4.500 1623.760 ;
        RECT 0.000 1607.360 2540.440 1622.160 ;
        RECT 0.000 1584.860 2540.440 1599.660 ;
        RECT 0.000 1583.260 4.500 1583.320 ;
        RECT 0.000 1578.700 4.500 1578.760 ;
        RECT 0.000 1562.360 2540.440 1577.160 ;
        RECT 0.000 1539.860 2540.440 1554.660 ;
        RECT 0.000 1538.260 4.500 1538.320 ;
        RECT 0.000 1533.700 4.500 1533.760 ;
        RECT 0.000 1517.360 2540.440 1532.160 ;
        RECT 0.000 1494.860 2540.440 1509.660 ;
        RECT 0.000 1493.260 4.500 1493.320 ;
        RECT 0.000 1488.700 4.500 1488.760 ;
        RECT 0.000 1472.360 2540.440 1487.160 ;
        RECT 0.000 1449.860 2540.440 1464.660 ;
        RECT 0.000 1448.260 4.500 1448.320 ;
        RECT 0.000 1443.700 4.500 1443.760 ;
        RECT 0.000 1427.360 2540.440 1442.160 ;
        RECT 0.000 1404.860 2540.440 1419.660 ;
        RECT 0.000 1403.260 4.500 1403.320 ;
        RECT 0.000 1398.700 4.500 1398.760 ;
        RECT 0.000 1382.360 2540.440 1397.160 ;
        RECT 0.000 1359.860 2540.440 1374.660 ;
        RECT 0.000 1358.260 4.500 1358.320 ;
        RECT 0.000 1353.700 4.500 1353.760 ;
        RECT 0.000 1337.360 2540.440 1352.160 ;
        RECT 0.000 1314.860 2540.440 1329.660 ;
        RECT 0.000 1313.260 4.500 1313.320 ;
        RECT 0.000 1308.700 4.500 1308.760 ;
        RECT 0.000 1292.360 2540.440 1307.160 ;
        RECT 0.000 1269.860 2540.440 1284.660 ;
        RECT 0.000 1268.260 4.500 1268.320 ;
        RECT 0.000 1263.700 4.500 1263.760 ;
        RECT 0.000 1247.360 2540.440 1262.160 ;
        RECT 0.000 1224.860 2540.440 1239.660 ;
        RECT 0.000 1223.260 4.500 1223.320 ;
        RECT 0.000 1218.700 4.500 1218.760 ;
        RECT 0.000 1202.360 2540.440 1217.160 ;
        RECT 0.000 1179.860 2540.440 1194.660 ;
        RECT 0.000 1178.260 4.500 1178.320 ;
        RECT 0.000 1173.700 4.500 1173.760 ;
        RECT 0.000 1157.360 2540.440 1172.160 ;
        RECT 0.000 1134.860 2540.440 1149.660 ;
        RECT 0.000 1133.260 4.500 1133.320 ;
        RECT 0.000 1128.700 4.500 1128.760 ;
        RECT 0.000 1112.360 2540.440 1127.160 ;
        RECT 0.000 1089.860 2540.440 1104.660 ;
        RECT 0.000 1088.260 4.500 1088.320 ;
        RECT 0.000 1083.700 4.500 1083.760 ;
        RECT 0.000 1067.360 2540.440 1082.160 ;
        RECT 0.000 1044.860 2540.440 1059.660 ;
        RECT 0.000 1043.260 4.500 1043.320 ;
        RECT 0.000 1038.700 4.500 1038.760 ;
        RECT 0.000 1022.360 2540.440 1037.160 ;
        RECT 0.000 999.860 2540.440 1014.660 ;
        RECT 0.000 998.260 4.500 998.320 ;
        RECT 0.000 993.700 4.500 993.760 ;
        RECT 0.000 977.360 2540.440 992.160 ;
        RECT 0.000 954.860 2540.440 969.660 ;
        RECT 0.000 953.260 4.500 953.320 ;
        RECT 0.000 948.700 4.500 948.760 ;
        RECT 0.000 932.360 2540.440 947.160 ;
        RECT 0.000 909.860 2540.440 924.660 ;
        RECT 0.000 908.260 4.500 908.320 ;
        RECT 0.000 903.700 4.500 903.760 ;
        RECT 0.000 887.360 2540.440 902.160 ;
        RECT 0.000 864.860 2540.440 879.660 ;
        RECT 0.000 863.260 4.500 863.320 ;
        RECT 0.000 858.700 4.500 858.760 ;
        RECT 0.000 842.360 2540.440 857.160 ;
        RECT 0.000 819.860 2540.440 834.660 ;
        RECT 0.000 818.260 4.500 818.320 ;
        RECT 0.000 813.700 4.500 813.760 ;
        RECT 0.000 797.360 2540.440 812.160 ;
        RECT 0.000 774.860 2540.440 789.660 ;
        RECT 0.000 773.260 4.500 773.320 ;
        RECT 0.000 768.700 4.500 768.760 ;
        RECT 0.000 752.360 2540.440 767.160 ;
        RECT 0.000 729.860 2540.440 744.660 ;
        RECT 0.000 728.260 4.500 728.320 ;
        RECT 0.000 723.700 4.500 723.760 ;
        RECT 0.000 707.360 2540.440 722.160 ;
        RECT 0.000 684.860 2540.440 699.660 ;
        RECT 0.000 683.260 4.500 683.320 ;
        RECT 0.000 678.700 4.500 678.760 ;
        RECT 0.000 662.360 2540.440 677.160 ;
        RECT 0.000 639.860 2540.440 654.660 ;
        RECT 0.000 638.260 4.500 638.320 ;
        RECT 0.000 633.700 4.500 633.760 ;
        RECT 0.000 617.360 2540.440 632.160 ;
        RECT 0.000 594.860 2540.440 609.660 ;
        RECT 0.000 593.260 4.500 593.320 ;
        RECT 0.000 588.700 4.500 588.760 ;
        RECT 0.000 572.360 2540.440 587.160 ;
        RECT 0.000 549.860 2540.440 564.660 ;
        RECT 0.000 548.260 4.500 548.320 ;
        RECT 0.000 543.700 4.500 543.760 ;
        RECT 0.000 527.360 2540.440 542.160 ;
        RECT 0.000 504.860 2540.440 519.660 ;
        RECT 0.000 503.260 4.500 503.320 ;
        RECT 0.000 498.700 4.500 498.760 ;
        RECT 0.000 482.360 2540.440 497.160 ;
        RECT 0.000 459.860 2540.440 474.660 ;
        RECT 0.000 458.260 4.500 458.320 ;
        RECT 0.000 453.700 4.500 453.760 ;
        RECT 0.000 437.360 2540.440 452.160 ;
        RECT 0.000 414.860 2540.440 429.660 ;
        RECT 0.000 413.260 4.500 413.320 ;
        RECT 0.000 408.700 4.500 408.760 ;
        RECT 0.000 392.360 2540.440 407.160 ;
        RECT 0.000 369.860 2540.440 384.660 ;
        RECT 0.000 368.260 4.500 368.320 ;
        RECT 0.000 363.700 4.500 363.760 ;
        RECT 0.000 347.360 2540.440 362.160 ;
        RECT 0.000 324.860 2540.440 339.660 ;
        RECT 0.000 323.260 4.500 323.320 ;
        RECT 0.000 318.700 4.500 318.760 ;
        RECT 0.000 302.360 2540.440 317.160 ;
        RECT 0.000 279.860 2540.440 294.660 ;
        RECT 0.000 278.260 4.500 278.320 ;
        RECT 0.000 273.700 4.500 273.760 ;
        RECT 0.000 257.360 2540.440 272.160 ;
        RECT 0.000 234.860 2540.440 249.660 ;
        RECT 0.000 233.260 4.500 233.320 ;
        RECT 0.000 228.700 4.500 228.760 ;
        RECT 0.000 212.360 2540.440 227.160 ;
        RECT 0.000 189.860 2540.440 204.660 ;
        RECT 0.000 188.260 4.500 188.320 ;
        RECT 0.000 183.700 4.500 183.760 ;
        RECT 0.000 167.360 2540.440 182.160 ;
        RECT 0.000 144.860 2540.440 159.660 ;
        RECT 0.000 143.260 4.500 143.320 ;
        RECT 0.000 138.700 4.500 138.760 ;
        RECT 0.000 122.360 2540.440 137.160 ;
        RECT 0.000 12.360 2540.440 114.660 ;
        RECT 0.000 6.160 4.600 12.360 ;
        RECT 2535.840 6.160 2540.440 12.360 ;
        RECT 0.000 4.560 4.500 4.620 ;
        RECT 0.000 0.000 4.500 0.060 ;
  END
END fpga_core
END LIBRARY

