magic
tech sky130A
magscale 1 2
timestamp 1680088215
<< obsli1 >>
rect 1104 2159 49864 24497
<< obsm1 >>
rect 1104 2128 49864 26376
<< metal2 >>
rect 1582 26200 1638 27000
rect 2226 26200 2282 27000
rect 2870 26200 2926 27000
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26200 4858 27000
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26200 7434 27000
rect 8022 26200 8078 27000
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26200 10654 27000
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26200 12586 27000
rect 13174 26200 13230 27000
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15750 26200 15806 27000
rect 16394 26200 16450 27000
rect 17038 26200 17094 27000
rect 17682 26200 17738 27000
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26200 20958 27000
rect 21546 26200 21602 27000
rect 22190 26200 22246 27000
rect 22834 26200 22890 27000
rect 23478 26200 23534 27000
rect 24122 26200 24178 27000
rect 24766 26200 24822 27000
rect 25410 26200 25466 27000
rect 26054 26200 26110 27000
rect 26698 26200 26754 27000
rect 27342 26200 27398 27000
rect 27986 26200 28042 27000
rect 28630 26200 28686 27000
rect 29274 26200 29330 27000
rect 29918 26200 29974 27000
rect 30562 26200 30618 27000
rect 31206 26200 31262 27000
rect 31850 26200 31906 27000
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26200 33838 27000
rect 34426 26200 34482 27000
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26200 36414 27000
rect 37002 26200 37058 27000
rect 37646 26200 37702 27000
rect 38290 26200 38346 27000
rect 38934 26200 38990 27000
rect 39578 26200 39634 27000
rect 40222 26200 40278 27000
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43442 26200 43498 27000
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26200 45430 27000
rect 46018 26200 46074 27000
rect 46662 26200 46718 27000
rect 47306 26200 47362 27000
rect 47950 26200 48006 27000
rect 48594 26200 48650 27000
rect 49238 26200 49294 27000
rect 1122 0 1178 800
rect 3238 0 3294 800
rect 5354 0 5410 800
rect 7470 0 7526 800
rect 9586 0 9642 800
rect 11702 0 11758 800
rect 13818 0 13874 800
rect 15934 0 15990 800
rect 18050 0 18106 800
rect 20166 0 20222 800
rect 22282 0 22338 800
rect 24398 0 24454 800
rect 26514 0 26570 800
rect 28630 0 28686 800
rect 30746 0 30802 800
rect 32862 0 32918 800
rect 34978 0 35034 800
rect 37094 0 37150 800
rect 39210 0 39266 800
rect 41326 0 41382 800
rect 43442 0 43498 800
rect 45558 0 45614 800
rect 47674 0 47730 800
rect 49790 0 49846 800
<< obsm2 >>
rect 1122 26144 1526 26382
rect 1694 26144 2170 26382
rect 2338 26144 2814 26382
rect 2982 26144 3458 26382
rect 3626 26144 4102 26382
rect 4270 26144 4746 26382
rect 4914 26144 5390 26382
rect 5558 26144 6034 26382
rect 6202 26144 6678 26382
rect 6846 26144 7322 26382
rect 7490 26144 7966 26382
rect 8134 26144 8610 26382
rect 8778 26144 9254 26382
rect 9422 26144 9898 26382
rect 10066 26144 10542 26382
rect 10710 26144 11186 26382
rect 11354 26144 11830 26382
rect 11998 26144 12474 26382
rect 12642 26144 13118 26382
rect 13286 26144 13762 26382
rect 13930 26144 14406 26382
rect 14574 26144 15050 26382
rect 15218 26144 15694 26382
rect 15862 26144 16338 26382
rect 16506 26144 16982 26382
rect 17150 26144 17626 26382
rect 17794 26144 18270 26382
rect 18438 26144 18914 26382
rect 19082 26144 19558 26382
rect 19726 26144 20202 26382
rect 20370 26144 20846 26382
rect 21014 26144 21490 26382
rect 21658 26144 22134 26382
rect 22302 26144 22778 26382
rect 22946 26144 23422 26382
rect 23590 26144 24066 26382
rect 24234 26144 24710 26382
rect 24878 26144 25354 26382
rect 25522 26144 25998 26382
rect 26166 26144 26642 26382
rect 26810 26144 27286 26382
rect 27454 26144 27930 26382
rect 28098 26144 28574 26382
rect 28742 26144 29218 26382
rect 29386 26144 29862 26382
rect 30030 26144 30506 26382
rect 30674 26144 31150 26382
rect 31318 26144 31794 26382
rect 31962 26144 32438 26382
rect 32606 26144 33082 26382
rect 33250 26144 33726 26382
rect 33894 26144 34370 26382
rect 34538 26144 35014 26382
rect 35182 26144 35658 26382
rect 35826 26144 36302 26382
rect 36470 26144 36946 26382
rect 37114 26144 37590 26382
rect 37758 26144 38234 26382
rect 38402 26144 38878 26382
rect 39046 26144 39522 26382
rect 39690 26144 40166 26382
rect 40334 26144 42098 26382
rect 42266 26144 42742 26382
rect 42910 26144 43386 26382
rect 43554 26144 44030 26382
rect 44198 26144 44674 26382
rect 44842 26144 45318 26382
rect 45486 26144 45962 26382
rect 46130 26144 46606 26382
rect 46774 26144 47250 26382
rect 47418 26144 47894 26382
rect 48062 26144 48538 26382
rect 48706 26144 49182 26382
rect 49350 26144 49844 26382
rect 1122 856 49844 26144
rect 1234 734 3182 856
rect 3350 734 5298 856
rect 5466 734 7414 856
rect 7582 734 9530 856
rect 9698 734 11646 856
rect 11814 734 13762 856
rect 13930 734 15878 856
rect 16046 734 17994 856
rect 18162 734 20110 856
rect 20278 734 22226 856
rect 22394 734 24342 856
rect 24510 734 26458 856
rect 26626 734 28574 856
rect 28742 734 30690 856
rect 30858 734 32806 856
rect 32974 734 34922 856
rect 35090 734 37038 856
rect 37206 734 39154 856
rect 39322 734 41270 856
rect 41438 734 43386 856
rect 43554 734 45502 856
rect 45670 734 47618 856
rect 47786 734 49734 856
<< metal3 >>
rect 0 25576 800 25696
rect 50200 25440 51000 25560
rect 0 25168 800 25288
rect 50200 25032 51000 25152
rect 0 24760 800 24880
rect 50200 24624 51000 24744
rect 0 24352 800 24472
rect 50200 24216 51000 24336
rect 0 23944 800 24064
rect 50200 23808 51000 23928
rect 0 23536 800 23656
rect 50200 23400 51000 23520
rect 0 23128 800 23248
rect 50200 22992 51000 23112
rect 0 22720 800 22840
rect 50200 22584 51000 22704
rect 0 22312 800 22432
rect 50200 22176 51000 22296
rect 0 21904 800 22024
rect 50200 21768 51000 21888
rect 0 21496 800 21616
rect 50200 21360 51000 21480
rect 0 21088 800 21208
rect 50200 20952 51000 21072
rect 0 20680 800 20800
rect 50200 20544 51000 20664
rect 0 20272 800 20392
rect 50200 20136 51000 20256
rect 0 19864 800 19984
rect 50200 19728 51000 19848
rect 0 19456 800 19576
rect 50200 19320 51000 19440
rect 0 19048 800 19168
rect 50200 18912 51000 19032
rect 0 18640 800 18760
rect 50200 18504 51000 18624
rect 0 18232 800 18352
rect 50200 18096 51000 18216
rect 0 17824 800 17944
rect 50200 17688 51000 17808
rect 0 17416 800 17536
rect 50200 17280 51000 17400
rect 0 17008 800 17128
rect 50200 16872 51000 16992
rect 0 16600 800 16720
rect 50200 16464 51000 16584
rect 0 16192 800 16312
rect 50200 16056 51000 16176
rect 0 15784 800 15904
rect 50200 15648 51000 15768
rect 0 15376 800 15496
rect 50200 15240 51000 15360
rect 0 14968 800 15088
rect 50200 14832 51000 14952
rect 0 14560 800 14680
rect 50200 14424 51000 14544
rect 0 14152 800 14272
rect 50200 14016 51000 14136
rect 0 13744 800 13864
rect 50200 13608 51000 13728
rect 0 13336 800 13456
rect 50200 13200 51000 13320
rect 0 12928 800 13048
rect 50200 12792 51000 12912
rect 0 12520 800 12640
rect 50200 12384 51000 12504
rect 0 12112 800 12232
rect 50200 11976 51000 12096
rect 0 11704 800 11824
rect 50200 11568 51000 11688
rect 0 11296 800 11416
rect 50200 11160 51000 11280
rect 0 10888 800 11008
rect 50200 10752 51000 10872
rect 0 10480 800 10600
rect 50200 10344 51000 10464
rect 0 10072 800 10192
rect 50200 9936 51000 10056
rect 0 9664 800 9784
rect 50200 9528 51000 9648
rect 0 9256 800 9376
rect 50200 9120 51000 9240
rect 0 8848 800 8968
rect 50200 8712 51000 8832
rect 0 8440 800 8560
rect 50200 8304 51000 8424
rect 0 8032 800 8152
rect 50200 7896 51000 8016
rect 0 7624 800 7744
rect 50200 7488 51000 7608
rect 0 7216 800 7336
rect 50200 7080 51000 7200
rect 0 6808 800 6928
rect 50200 6672 51000 6792
rect 0 6400 800 6520
rect 50200 6264 51000 6384
rect 0 5992 800 6112
rect 50200 5856 51000 5976
rect 0 5584 800 5704
rect 50200 5448 51000 5568
rect 0 5176 800 5296
rect 50200 5040 51000 5160
rect 0 4768 800 4888
rect 50200 4632 51000 4752
rect 0 4360 800 4480
rect 50200 4224 51000 4344
rect 0 3952 800 4072
rect 50200 3816 51000 3936
rect 0 3544 800 3664
rect 50200 3408 51000 3528
rect 0 3136 800 3256
rect 50200 3000 51000 3120
rect 0 2728 800 2848
rect 50200 2592 51000 2712
rect 0 2320 800 2440
rect 50200 2184 51000 2304
rect 0 1912 800 2032
rect 50200 1776 51000 1896
rect 0 1504 800 1624
rect 50200 1368 51000 1488
<< obsm3 >>
rect 880 25640 50200 25669
rect 880 25496 50120 25640
rect 800 25368 50120 25496
rect 880 25360 50120 25368
rect 880 25232 50200 25360
rect 880 25088 50120 25232
rect 800 24960 50120 25088
rect 880 24952 50120 24960
rect 880 24824 50200 24952
rect 880 24680 50120 24824
rect 800 24552 50120 24680
rect 880 24544 50120 24552
rect 880 24416 50200 24544
rect 880 24272 50120 24416
rect 800 24144 50120 24272
rect 880 24136 50120 24144
rect 880 24008 50200 24136
rect 880 23864 50120 24008
rect 800 23736 50120 23864
rect 880 23728 50120 23736
rect 880 23600 50200 23728
rect 880 23456 50120 23600
rect 800 23328 50120 23456
rect 880 23320 50120 23328
rect 880 23192 50200 23320
rect 880 23048 50120 23192
rect 800 22920 50120 23048
rect 880 22912 50120 22920
rect 880 22784 50200 22912
rect 880 22640 50120 22784
rect 800 22512 50120 22640
rect 880 22504 50120 22512
rect 880 22376 50200 22504
rect 880 22232 50120 22376
rect 800 22104 50120 22232
rect 880 22096 50120 22104
rect 880 21968 50200 22096
rect 880 21824 50120 21968
rect 800 21696 50120 21824
rect 880 21688 50120 21696
rect 880 21560 50200 21688
rect 880 21416 50120 21560
rect 800 21288 50120 21416
rect 880 21280 50120 21288
rect 880 21152 50200 21280
rect 880 21008 50120 21152
rect 800 20880 50120 21008
rect 880 20872 50120 20880
rect 880 20744 50200 20872
rect 880 20600 50120 20744
rect 800 20472 50120 20600
rect 880 20464 50120 20472
rect 880 20336 50200 20464
rect 880 20192 50120 20336
rect 800 20064 50120 20192
rect 880 20056 50120 20064
rect 880 19928 50200 20056
rect 880 19784 50120 19928
rect 800 19656 50120 19784
rect 880 19648 50120 19656
rect 880 19520 50200 19648
rect 880 19376 50120 19520
rect 800 19248 50120 19376
rect 880 19240 50120 19248
rect 880 19112 50200 19240
rect 880 18968 50120 19112
rect 800 18840 50120 18968
rect 880 18832 50120 18840
rect 880 18704 50200 18832
rect 880 18560 50120 18704
rect 800 18432 50120 18560
rect 880 18424 50120 18432
rect 880 18296 50200 18424
rect 880 18152 50120 18296
rect 800 18024 50120 18152
rect 880 18016 50120 18024
rect 880 17888 50200 18016
rect 880 17744 50120 17888
rect 800 17616 50120 17744
rect 880 17608 50120 17616
rect 880 17480 50200 17608
rect 880 17336 50120 17480
rect 800 17208 50120 17336
rect 880 17200 50120 17208
rect 880 17072 50200 17200
rect 880 16928 50120 17072
rect 800 16800 50120 16928
rect 880 16792 50120 16800
rect 880 16664 50200 16792
rect 880 16520 50120 16664
rect 800 16392 50120 16520
rect 880 16384 50120 16392
rect 880 16256 50200 16384
rect 880 16112 50120 16256
rect 800 15984 50120 16112
rect 880 15976 50120 15984
rect 880 15848 50200 15976
rect 880 15704 50120 15848
rect 800 15576 50120 15704
rect 880 15568 50120 15576
rect 880 15440 50200 15568
rect 880 15296 50120 15440
rect 800 15168 50120 15296
rect 880 15160 50120 15168
rect 880 15032 50200 15160
rect 880 14888 50120 15032
rect 800 14760 50120 14888
rect 880 14752 50120 14760
rect 880 14624 50200 14752
rect 880 14480 50120 14624
rect 800 14352 50120 14480
rect 880 14344 50120 14352
rect 880 14216 50200 14344
rect 880 14072 50120 14216
rect 800 13944 50120 14072
rect 880 13936 50120 13944
rect 880 13808 50200 13936
rect 880 13664 50120 13808
rect 800 13536 50120 13664
rect 880 13528 50120 13536
rect 880 13400 50200 13528
rect 880 13256 50120 13400
rect 800 13128 50120 13256
rect 880 13120 50120 13128
rect 880 12992 50200 13120
rect 880 12848 50120 12992
rect 800 12720 50120 12848
rect 880 12712 50120 12720
rect 880 12584 50200 12712
rect 880 12440 50120 12584
rect 800 12312 50120 12440
rect 880 12304 50120 12312
rect 880 12176 50200 12304
rect 880 12032 50120 12176
rect 800 11904 50120 12032
rect 880 11896 50120 11904
rect 880 11768 50200 11896
rect 880 11624 50120 11768
rect 800 11496 50120 11624
rect 880 11488 50120 11496
rect 880 11360 50200 11488
rect 880 11216 50120 11360
rect 800 11088 50120 11216
rect 880 11080 50120 11088
rect 880 10952 50200 11080
rect 880 10808 50120 10952
rect 800 10680 50120 10808
rect 880 10672 50120 10680
rect 880 10544 50200 10672
rect 880 10400 50120 10544
rect 800 10272 50120 10400
rect 880 10264 50120 10272
rect 880 10136 50200 10264
rect 880 9992 50120 10136
rect 800 9864 50120 9992
rect 880 9856 50120 9864
rect 880 9728 50200 9856
rect 880 9584 50120 9728
rect 800 9456 50120 9584
rect 880 9448 50120 9456
rect 880 9320 50200 9448
rect 880 9176 50120 9320
rect 800 9048 50120 9176
rect 880 9040 50120 9048
rect 880 8912 50200 9040
rect 880 8768 50120 8912
rect 800 8640 50120 8768
rect 880 8632 50120 8640
rect 880 8504 50200 8632
rect 880 8360 50120 8504
rect 800 8232 50120 8360
rect 880 8224 50120 8232
rect 880 8096 50200 8224
rect 880 7952 50120 8096
rect 800 7824 50120 7952
rect 880 7816 50120 7824
rect 880 7688 50200 7816
rect 880 7544 50120 7688
rect 800 7416 50120 7544
rect 880 7408 50120 7416
rect 880 7280 50200 7408
rect 880 7136 50120 7280
rect 800 7008 50120 7136
rect 880 7000 50120 7008
rect 880 6872 50200 7000
rect 880 6728 50120 6872
rect 800 6600 50120 6728
rect 880 6592 50120 6600
rect 880 6464 50200 6592
rect 880 6320 50120 6464
rect 800 6192 50120 6320
rect 880 6184 50120 6192
rect 880 6056 50200 6184
rect 880 5912 50120 6056
rect 800 5784 50120 5912
rect 880 5776 50120 5784
rect 880 5648 50200 5776
rect 880 5504 50120 5648
rect 800 5376 50120 5504
rect 880 5368 50120 5376
rect 880 5240 50200 5368
rect 880 5096 50120 5240
rect 800 4968 50120 5096
rect 880 4960 50120 4968
rect 880 4832 50200 4960
rect 880 4688 50120 4832
rect 800 4560 50120 4688
rect 880 4552 50120 4560
rect 880 4424 50200 4552
rect 880 4280 50120 4424
rect 800 4152 50120 4280
rect 880 4144 50120 4152
rect 880 4016 50200 4144
rect 880 3872 50120 4016
rect 800 3744 50120 3872
rect 880 3736 50120 3744
rect 880 3608 50200 3736
rect 880 3464 50120 3608
rect 800 3336 50120 3464
rect 880 3328 50120 3336
rect 880 3200 50200 3328
rect 880 3056 50120 3200
rect 800 2928 50120 3056
rect 880 2920 50120 2928
rect 880 2792 50200 2920
rect 880 2648 50120 2792
rect 800 2520 50120 2648
rect 880 2512 50120 2520
rect 880 2384 50200 2512
rect 880 2240 50120 2384
rect 800 2112 50120 2240
rect 880 2104 50120 2112
rect 880 1976 50200 2104
rect 880 1832 50120 1976
rect 800 1704 50120 1832
rect 880 1696 50120 1704
rect 880 1568 50200 1696
rect 880 1424 50120 1568
rect 800 1395 50120 1424
<< metal4 >>
rect 2944 2128 3264 24528
rect 7944 2128 8264 24528
rect 12944 2128 13264 24528
rect 17944 2128 18264 24528
rect 22944 2128 23264 24528
rect 27944 2128 28264 24528
rect 32944 2128 33264 24528
rect 37944 2128 38264 24528
rect 42944 2128 43264 24528
rect 47944 2128 48264 24528
<< obsm4 >>
rect 14043 9011 17864 24037
rect 18344 9011 22864 24037
rect 23344 9011 27864 24037
rect 28344 9011 32864 24037
rect 33344 9011 37864 24037
rect 38344 9011 38581 24037
<< labels >>
rlabel metal4 s 7944 2128 8264 24528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17944 2128 18264 24528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27944 2128 28264 24528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37944 2128 38264 24528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47944 2128 48264 24528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2944 2128 3264 24528 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12944 2128 13264 24528 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 22944 2128 23264 24528 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 32944 2128 33264 24528 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 42944 2128 43264 24528 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 9586 0 9642 800 6 ccff_head
port 3 nsew signal input
rlabel metal2 s 49238 26200 49294 27000 6 ccff_head_1
port 4 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 ccff_tail
port 5 nsew signal output
rlabel metal2 s 1582 26200 1638 27000 6 ccff_tail_0
port 6 nsew signal output
rlabel metal3 s 0 1504 800 1624 6 chanx_left_in[0]
port 7 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 chanx_left_in[10]
port 8 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 chanx_left_in[11]
port 9 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 chanx_left_in[12]
port 10 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 chanx_left_in[13]
port 11 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 chanx_left_in[14]
port 12 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[15]
port 13 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[16]
port 14 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 chanx_left_in[17]
port 15 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 chanx_left_in[18]
port 16 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[19]
port 17 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 chanx_left_in[1]
port 18 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[20]
port 19 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[21]
port 20 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 chanx_left_in[22]
port 21 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[23]
port 22 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[24]
port 23 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 chanx_left_in[25]
port 24 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 chanx_left_in[26]
port 25 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 chanx_left_in[27]
port 26 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 chanx_left_in[28]
port 27 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 chanx_left_in[29]
port 28 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 chanx_left_in[2]
port 29 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 chanx_left_in[3]
port 30 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 chanx_left_in[4]
port 31 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 chanx_left_in[5]
port 32 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 chanx_left_in[6]
port 33 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[7]
port 34 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[8]
port 35 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[9]
port 36 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[0]
port 37 nsew signal output
rlabel metal3 s 0 17824 800 17944 6 chanx_left_out[10]
port 38 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 chanx_left_out[11]
port 39 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 chanx_left_out[12]
port 40 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 chanx_left_out[13]
port 41 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 chanx_left_out[14]
port 42 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 chanx_left_out[15]
port 43 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[16]
port 44 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[17]
port 45 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 chanx_left_out[18]
port 46 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 chanx_left_out[19]
port 47 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[1]
port 48 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 chanx_left_out[20]
port 49 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 chanx_left_out[21]
port 50 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 chanx_left_out[22]
port 51 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 chanx_left_out[23]
port 52 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 chanx_left_out[24]
port 53 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 chanx_left_out[25]
port 54 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 chanx_left_out[26]
port 55 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 chanx_left_out[27]
port 56 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 chanx_left_out[28]
port 57 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 chanx_left_out[29]
port 58 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[2]
port 59 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[3]
port 60 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 chanx_left_out[4]
port 61 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 chanx_left_out[5]
port 62 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 chanx_left_out[6]
port 63 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 chanx_left_out[7]
port 64 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[8]
port 65 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[9]
port 66 nsew signal output
rlabel metal3 s 50200 13608 51000 13728 6 chanx_right_in_0[0]
port 67 nsew signal input
rlabel metal3 s 50200 17688 51000 17808 6 chanx_right_in_0[10]
port 68 nsew signal input
rlabel metal3 s 50200 18096 51000 18216 6 chanx_right_in_0[11]
port 69 nsew signal input
rlabel metal3 s 50200 18504 51000 18624 6 chanx_right_in_0[12]
port 70 nsew signal input
rlabel metal3 s 50200 18912 51000 19032 6 chanx_right_in_0[13]
port 71 nsew signal input
rlabel metal3 s 50200 19320 51000 19440 6 chanx_right_in_0[14]
port 72 nsew signal input
rlabel metal3 s 50200 19728 51000 19848 6 chanx_right_in_0[15]
port 73 nsew signal input
rlabel metal3 s 50200 20136 51000 20256 6 chanx_right_in_0[16]
port 74 nsew signal input
rlabel metal3 s 50200 20544 51000 20664 6 chanx_right_in_0[17]
port 75 nsew signal input
rlabel metal3 s 50200 20952 51000 21072 6 chanx_right_in_0[18]
port 76 nsew signal input
rlabel metal3 s 50200 21360 51000 21480 6 chanx_right_in_0[19]
port 77 nsew signal input
rlabel metal3 s 50200 14016 51000 14136 6 chanx_right_in_0[1]
port 78 nsew signal input
rlabel metal3 s 50200 21768 51000 21888 6 chanx_right_in_0[20]
port 79 nsew signal input
rlabel metal3 s 50200 22176 51000 22296 6 chanx_right_in_0[21]
port 80 nsew signal input
rlabel metal3 s 50200 22584 51000 22704 6 chanx_right_in_0[22]
port 81 nsew signal input
rlabel metal3 s 50200 22992 51000 23112 6 chanx_right_in_0[23]
port 82 nsew signal input
rlabel metal3 s 50200 23400 51000 23520 6 chanx_right_in_0[24]
port 83 nsew signal input
rlabel metal3 s 50200 23808 51000 23928 6 chanx_right_in_0[25]
port 84 nsew signal input
rlabel metal3 s 50200 24216 51000 24336 6 chanx_right_in_0[26]
port 85 nsew signal input
rlabel metal3 s 50200 24624 51000 24744 6 chanx_right_in_0[27]
port 86 nsew signal input
rlabel metal3 s 50200 25032 51000 25152 6 chanx_right_in_0[28]
port 87 nsew signal input
rlabel metal3 s 50200 25440 51000 25560 6 chanx_right_in_0[29]
port 88 nsew signal input
rlabel metal3 s 50200 14424 51000 14544 6 chanx_right_in_0[2]
port 89 nsew signal input
rlabel metal3 s 50200 14832 51000 14952 6 chanx_right_in_0[3]
port 90 nsew signal input
rlabel metal3 s 50200 15240 51000 15360 6 chanx_right_in_0[4]
port 91 nsew signal input
rlabel metal3 s 50200 15648 51000 15768 6 chanx_right_in_0[5]
port 92 nsew signal input
rlabel metal3 s 50200 16056 51000 16176 6 chanx_right_in_0[6]
port 93 nsew signal input
rlabel metal3 s 50200 16464 51000 16584 6 chanx_right_in_0[7]
port 94 nsew signal input
rlabel metal3 s 50200 16872 51000 16992 6 chanx_right_in_0[8]
port 95 nsew signal input
rlabel metal3 s 50200 17280 51000 17400 6 chanx_right_in_0[9]
port 96 nsew signal input
rlabel metal3 s 50200 1368 51000 1488 6 chanx_right_out_0[0]
port 97 nsew signal output
rlabel metal3 s 50200 5448 51000 5568 6 chanx_right_out_0[10]
port 98 nsew signal output
rlabel metal3 s 50200 5856 51000 5976 6 chanx_right_out_0[11]
port 99 nsew signal output
rlabel metal3 s 50200 6264 51000 6384 6 chanx_right_out_0[12]
port 100 nsew signal output
rlabel metal3 s 50200 6672 51000 6792 6 chanx_right_out_0[13]
port 101 nsew signal output
rlabel metal3 s 50200 7080 51000 7200 6 chanx_right_out_0[14]
port 102 nsew signal output
rlabel metal3 s 50200 7488 51000 7608 6 chanx_right_out_0[15]
port 103 nsew signal output
rlabel metal3 s 50200 7896 51000 8016 6 chanx_right_out_0[16]
port 104 nsew signal output
rlabel metal3 s 50200 8304 51000 8424 6 chanx_right_out_0[17]
port 105 nsew signal output
rlabel metal3 s 50200 8712 51000 8832 6 chanx_right_out_0[18]
port 106 nsew signal output
rlabel metal3 s 50200 9120 51000 9240 6 chanx_right_out_0[19]
port 107 nsew signal output
rlabel metal3 s 50200 1776 51000 1896 6 chanx_right_out_0[1]
port 108 nsew signal output
rlabel metal3 s 50200 9528 51000 9648 6 chanx_right_out_0[20]
port 109 nsew signal output
rlabel metal3 s 50200 9936 51000 10056 6 chanx_right_out_0[21]
port 110 nsew signal output
rlabel metal3 s 50200 10344 51000 10464 6 chanx_right_out_0[22]
port 111 nsew signal output
rlabel metal3 s 50200 10752 51000 10872 6 chanx_right_out_0[23]
port 112 nsew signal output
rlabel metal3 s 50200 11160 51000 11280 6 chanx_right_out_0[24]
port 113 nsew signal output
rlabel metal3 s 50200 11568 51000 11688 6 chanx_right_out_0[25]
port 114 nsew signal output
rlabel metal3 s 50200 11976 51000 12096 6 chanx_right_out_0[26]
port 115 nsew signal output
rlabel metal3 s 50200 12384 51000 12504 6 chanx_right_out_0[27]
port 116 nsew signal output
rlabel metal3 s 50200 12792 51000 12912 6 chanx_right_out_0[28]
port 117 nsew signal output
rlabel metal3 s 50200 13200 51000 13320 6 chanx_right_out_0[29]
port 118 nsew signal output
rlabel metal3 s 50200 2184 51000 2304 6 chanx_right_out_0[2]
port 119 nsew signal output
rlabel metal3 s 50200 2592 51000 2712 6 chanx_right_out_0[3]
port 120 nsew signal output
rlabel metal3 s 50200 3000 51000 3120 6 chanx_right_out_0[4]
port 121 nsew signal output
rlabel metal3 s 50200 3408 51000 3528 6 chanx_right_out_0[5]
port 122 nsew signal output
rlabel metal3 s 50200 3816 51000 3936 6 chanx_right_out_0[6]
port 123 nsew signal output
rlabel metal3 s 50200 4224 51000 4344 6 chanx_right_out_0[7]
port 124 nsew signal output
rlabel metal3 s 50200 4632 51000 4752 6 chanx_right_out_0[8]
port 125 nsew signal output
rlabel metal3 s 50200 5040 51000 5160 6 chanx_right_out_0[9]
port 126 nsew signal output
rlabel metal2 s 21546 26200 21602 27000 6 chany_top_in[0]
port 127 nsew signal input
rlabel metal2 s 27986 26200 28042 27000 6 chany_top_in[10]
port 128 nsew signal input
rlabel metal2 s 28630 26200 28686 27000 6 chany_top_in[11]
port 129 nsew signal input
rlabel metal2 s 29274 26200 29330 27000 6 chany_top_in[12]
port 130 nsew signal input
rlabel metal2 s 29918 26200 29974 27000 6 chany_top_in[13]
port 131 nsew signal input
rlabel metal2 s 30562 26200 30618 27000 6 chany_top_in[14]
port 132 nsew signal input
rlabel metal2 s 31206 26200 31262 27000 6 chany_top_in[15]
port 133 nsew signal input
rlabel metal2 s 31850 26200 31906 27000 6 chany_top_in[16]
port 134 nsew signal input
rlabel metal2 s 32494 26200 32550 27000 6 chany_top_in[17]
port 135 nsew signal input
rlabel metal2 s 33138 26200 33194 27000 6 chany_top_in[18]
port 136 nsew signal input
rlabel metal2 s 33782 26200 33838 27000 6 chany_top_in[19]
port 137 nsew signal input
rlabel metal2 s 22190 26200 22246 27000 6 chany_top_in[1]
port 138 nsew signal input
rlabel metal2 s 34426 26200 34482 27000 6 chany_top_in[20]
port 139 nsew signal input
rlabel metal2 s 35070 26200 35126 27000 6 chany_top_in[21]
port 140 nsew signal input
rlabel metal2 s 35714 26200 35770 27000 6 chany_top_in[22]
port 141 nsew signal input
rlabel metal2 s 36358 26200 36414 27000 6 chany_top_in[23]
port 142 nsew signal input
rlabel metal2 s 37002 26200 37058 27000 6 chany_top_in[24]
port 143 nsew signal input
rlabel metal2 s 37646 26200 37702 27000 6 chany_top_in[25]
port 144 nsew signal input
rlabel metal2 s 38290 26200 38346 27000 6 chany_top_in[26]
port 145 nsew signal input
rlabel metal2 s 38934 26200 38990 27000 6 chany_top_in[27]
port 146 nsew signal input
rlabel metal2 s 39578 26200 39634 27000 6 chany_top_in[28]
port 147 nsew signal input
rlabel metal2 s 40222 26200 40278 27000 6 chany_top_in[29]
port 148 nsew signal input
rlabel metal2 s 22834 26200 22890 27000 6 chany_top_in[2]
port 149 nsew signal input
rlabel metal2 s 23478 26200 23534 27000 6 chany_top_in[3]
port 150 nsew signal input
rlabel metal2 s 24122 26200 24178 27000 6 chany_top_in[4]
port 151 nsew signal input
rlabel metal2 s 24766 26200 24822 27000 6 chany_top_in[5]
port 152 nsew signal input
rlabel metal2 s 25410 26200 25466 27000 6 chany_top_in[6]
port 153 nsew signal input
rlabel metal2 s 26054 26200 26110 27000 6 chany_top_in[7]
port 154 nsew signal input
rlabel metal2 s 26698 26200 26754 27000 6 chany_top_in[8]
port 155 nsew signal input
rlabel metal2 s 27342 26200 27398 27000 6 chany_top_in[9]
port 156 nsew signal input
rlabel metal2 s 2226 26200 2282 27000 6 chany_top_out[0]
port 157 nsew signal output
rlabel metal2 s 8666 26200 8722 27000 6 chany_top_out[10]
port 158 nsew signal output
rlabel metal2 s 9310 26200 9366 27000 6 chany_top_out[11]
port 159 nsew signal output
rlabel metal2 s 9954 26200 10010 27000 6 chany_top_out[12]
port 160 nsew signal output
rlabel metal2 s 10598 26200 10654 27000 6 chany_top_out[13]
port 161 nsew signal output
rlabel metal2 s 11242 26200 11298 27000 6 chany_top_out[14]
port 162 nsew signal output
rlabel metal2 s 11886 26200 11942 27000 6 chany_top_out[15]
port 163 nsew signal output
rlabel metal2 s 12530 26200 12586 27000 6 chany_top_out[16]
port 164 nsew signal output
rlabel metal2 s 13174 26200 13230 27000 6 chany_top_out[17]
port 165 nsew signal output
rlabel metal2 s 13818 26200 13874 27000 6 chany_top_out[18]
port 166 nsew signal output
rlabel metal2 s 14462 26200 14518 27000 6 chany_top_out[19]
port 167 nsew signal output
rlabel metal2 s 2870 26200 2926 27000 6 chany_top_out[1]
port 168 nsew signal output
rlabel metal2 s 15106 26200 15162 27000 6 chany_top_out[20]
port 169 nsew signal output
rlabel metal2 s 15750 26200 15806 27000 6 chany_top_out[21]
port 170 nsew signal output
rlabel metal2 s 16394 26200 16450 27000 6 chany_top_out[22]
port 171 nsew signal output
rlabel metal2 s 17038 26200 17094 27000 6 chany_top_out[23]
port 172 nsew signal output
rlabel metal2 s 17682 26200 17738 27000 6 chany_top_out[24]
port 173 nsew signal output
rlabel metal2 s 18326 26200 18382 27000 6 chany_top_out[25]
port 174 nsew signal output
rlabel metal2 s 18970 26200 19026 27000 6 chany_top_out[26]
port 175 nsew signal output
rlabel metal2 s 19614 26200 19670 27000 6 chany_top_out[27]
port 176 nsew signal output
rlabel metal2 s 20258 26200 20314 27000 6 chany_top_out[28]
port 177 nsew signal output
rlabel metal2 s 20902 26200 20958 27000 6 chany_top_out[29]
port 178 nsew signal output
rlabel metal2 s 3514 26200 3570 27000 6 chany_top_out[2]
port 179 nsew signal output
rlabel metal2 s 4158 26200 4214 27000 6 chany_top_out[3]
port 180 nsew signal output
rlabel metal2 s 4802 26200 4858 27000 6 chany_top_out[4]
port 181 nsew signal output
rlabel metal2 s 5446 26200 5502 27000 6 chany_top_out[5]
port 182 nsew signal output
rlabel metal2 s 6090 26200 6146 27000 6 chany_top_out[6]
port 183 nsew signal output
rlabel metal2 s 6734 26200 6790 27000 6 chany_top_out[7]
port 184 nsew signal output
rlabel metal2 s 7378 26200 7434 27000 6 chany_top_out[8]
port 185 nsew signal output
rlabel metal2 s 8022 26200 8078 27000 6 chany_top_out[9]
port 186 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 gfpga_pad_io_soc_dir[0]
port 187 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 gfpga_pad_io_soc_dir[1]
port 188 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 gfpga_pad_io_soc_dir[2]
port 189 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 gfpga_pad_io_soc_dir[3]
port 190 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 gfpga_pad_io_soc_in[0]
port 191 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 gfpga_pad_io_soc_in[1]
port 192 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 gfpga_pad_io_soc_in[2]
port 193 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 gfpga_pad_io_soc_in[3]
port 194 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 gfpga_pad_io_soc_out[0]
port 195 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 gfpga_pad_io_soc_out[1]
port 196 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 gfpga_pad_io_soc_out[2]
port 197 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 gfpga_pad_io_soc_out[3]
port 198 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 isol_n
port 199 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 prog_clk
port 200 nsew signal input
rlabel metal2 s 42154 26200 42210 27000 6 prog_reset_top_in
port 201 nsew signal input
rlabel metal2 s 42798 26200 42854 27000 6 reset_top_in
port 202 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 203 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 204 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 205 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 206 nsew signal input
rlabel metal2 s 43442 26200 43498 27000 6 test_enable_top_in
port 207 nsew signal input
rlabel metal2 s 45374 26200 45430 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 208 nsew signal input
rlabel metal2 s 46018 26200 46074 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 209 nsew signal input
rlabel metal2 s 46662 26200 46718 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 210 nsew signal input
rlabel metal2 s 47306 26200 47362 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 211 nsew signal input
rlabel metal2 s 47950 26200 48006 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 212 nsew signal input
rlabel metal2 s 48594 26200 48650 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 213 nsew signal input
rlabel metal2 s 44086 26200 44142 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 214 nsew signal input
rlabel metal2 s 44730 26200 44786 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 215 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 top_width_0_height_0_subtile_0__pin_inpad_0_
port 216 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 top_width_0_height_0_subtile_1__pin_inpad_0_
port 217 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 top_width_0_height_0_subtile_2__pin_inpad_0_
port 218 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 top_width_0_height_0_subtile_3__pin_inpad_0_
port 219 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 51000 27000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2876800
string GDS_FILE /home/hosni/OpenFPGA/clear/openlane/bottom_tile/runs/23_03_29_04_08/results/signoff/bottom_tile.magic.gds
string GDS_START 165170
<< end >>

