magic
tech sky130A
magscale 1 2
timestamp 1656945641
<< obsli1 >>
rect 1104 2159 21896 20689
<< obsm1 >>
rect 382 2128 22526 20720
<< metal2 >>
rect 386 22200 442 23000
rect 938 22200 994 23000
rect 1490 22200 1546 23000
rect 2042 22200 2098 23000
rect 2594 22200 2650 23000
rect 3146 22200 3202 23000
rect 3698 22200 3754 23000
rect 4250 22200 4306 23000
rect 4802 22200 4858 23000
rect 5354 22200 5410 23000
rect 5906 22200 5962 23000
rect 6458 22200 6514 23000
rect 7010 22200 7066 23000
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10874 22200 10930 23000
rect 11426 22200 11482 23000
rect 11978 22200 12034 23000
rect 12530 22200 12586 23000
rect 13082 22200 13138 23000
rect 13634 22200 13690 23000
rect 14186 22200 14242 23000
rect 14738 22200 14794 23000
rect 15290 22200 15346 23000
rect 15842 22200 15898 23000
rect 16394 22200 16450 23000
rect 16946 22200 17002 23000
rect 17498 22200 17554 23000
rect 18050 22200 18106 23000
rect 18602 22200 18658 23000
rect 19154 22200 19210 23000
rect 19706 22200 19762 23000
rect 20258 22200 20314 23000
rect 20810 22200 20866 23000
rect 21362 22200 21418 23000
rect 21914 22200 21970 23000
rect 22466 22200 22522 23000
<< obsm2 >>
rect 498 22144 882 22250
rect 1050 22144 1434 22250
rect 1602 22144 1986 22250
rect 2154 22144 2538 22250
rect 2706 22144 3090 22250
rect 3258 22144 3642 22250
rect 3810 22144 4194 22250
rect 4362 22144 4746 22250
rect 4914 22144 5298 22250
rect 5466 22144 5850 22250
rect 6018 22144 6402 22250
rect 6570 22144 6954 22250
rect 7122 22144 7506 22250
rect 7674 22144 8058 22250
rect 8226 22144 8610 22250
rect 8778 22144 9162 22250
rect 9330 22144 9714 22250
rect 9882 22144 10266 22250
rect 10434 22144 10818 22250
rect 10986 22144 11370 22250
rect 11538 22144 11922 22250
rect 12090 22144 12474 22250
rect 12642 22144 13026 22250
rect 13194 22144 13578 22250
rect 13746 22144 14130 22250
rect 14298 22144 14682 22250
rect 14850 22144 15234 22250
rect 15402 22144 15786 22250
rect 15954 22144 16338 22250
rect 16506 22144 16890 22250
rect 17058 22144 17442 22250
rect 17610 22144 17994 22250
rect 18162 22144 18546 22250
rect 18714 22144 19098 22250
rect 19266 22144 19650 22250
rect 19818 22144 20202 22250
rect 20370 22144 20754 22250
rect 20922 22144 21306 22250
rect 21474 22144 21858 22250
rect 22026 22144 22410 22250
rect 388 1391 22520 22144
<< metal3 >>
rect 22200 21360 23000 21480
rect 22200 20952 23000 21072
rect 22200 20544 23000 20664
rect 22200 20136 23000 20256
rect 22200 19728 23000 19848
rect 22200 19320 23000 19440
rect 22200 18912 23000 19032
rect 22200 18504 23000 18624
rect 22200 18096 23000 18216
rect 22200 17688 23000 17808
rect 0 17144 800 17264
rect 22200 17280 23000 17400
rect 22200 16872 23000 16992
rect 22200 16464 23000 16584
rect 22200 16056 23000 16176
rect 22200 15648 23000 15768
rect 22200 15240 23000 15360
rect 22200 14832 23000 14952
rect 22200 14424 23000 14544
rect 22200 14016 23000 14136
rect 22200 13608 23000 13728
rect 22200 13200 23000 13320
rect 22200 12792 23000 12912
rect 22200 12384 23000 12504
rect 22200 11976 23000 12096
rect 22200 11568 23000 11688
rect 22200 11160 23000 11280
rect 22200 10752 23000 10872
rect 22200 10344 23000 10464
rect 22200 9936 23000 10056
rect 22200 9528 23000 9648
rect 22200 9120 23000 9240
rect 22200 8712 23000 8832
rect 22200 8304 23000 8424
rect 22200 7896 23000 8016
rect 22200 7488 23000 7608
rect 22200 7080 23000 7200
rect 22200 6672 23000 6792
rect 22200 6264 23000 6384
rect 0 5720 800 5840
rect 22200 5856 23000 5976
rect 22200 5448 23000 5568
rect 22200 5040 23000 5160
rect 22200 4632 23000 4752
rect 22200 4224 23000 4344
rect 22200 3816 23000 3936
rect 22200 3408 23000 3528
rect 22200 3000 23000 3120
rect 22200 2592 23000 2712
rect 22200 2184 23000 2304
rect 22200 1776 23000 1896
rect 22200 1368 23000 1488
<< obsm3 >>
rect 800 21280 22120 21453
rect 800 21152 22202 21280
rect 800 20872 22120 21152
rect 800 20744 22202 20872
rect 800 20464 22120 20744
rect 800 20336 22202 20464
rect 800 20056 22120 20336
rect 800 19928 22202 20056
rect 800 19648 22120 19928
rect 800 19520 22202 19648
rect 800 19240 22120 19520
rect 800 19112 22202 19240
rect 800 18832 22120 19112
rect 800 18704 22202 18832
rect 800 18424 22120 18704
rect 800 18296 22202 18424
rect 800 18016 22120 18296
rect 800 17888 22202 18016
rect 800 17608 22120 17888
rect 800 17480 22202 17608
rect 800 17344 22120 17480
rect 880 17200 22120 17344
rect 880 17072 22202 17200
rect 880 17064 22120 17072
rect 800 16792 22120 17064
rect 800 16664 22202 16792
rect 800 16384 22120 16664
rect 800 16256 22202 16384
rect 800 15976 22120 16256
rect 800 15848 22202 15976
rect 800 15568 22120 15848
rect 800 15440 22202 15568
rect 800 15160 22120 15440
rect 800 15032 22202 15160
rect 800 14752 22120 15032
rect 800 14624 22202 14752
rect 800 14344 22120 14624
rect 800 14216 22202 14344
rect 800 13936 22120 14216
rect 800 13808 22202 13936
rect 800 13528 22120 13808
rect 800 13400 22202 13528
rect 800 13120 22120 13400
rect 800 12992 22202 13120
rect 800 12712 22120 12992
rect 800 12584 22202 12712
rect 800 12304 22120 12584
rect 800 12176 22202 12304
rect 800 11896 22120 12176
rect 800 11768 22202 11896
rect 800 11488 22120 11768
rect 800 11360 22202 11488
rect 800 11080 22120 11360
rect 800 10952 22202 11080
rect 800 10672 22120 10952
rect 800 10544 22202 10672
rect 800 10264 22120 10544
rect 800 10136 22202 10264
rect 800 9856 22120 10136
rect 800 9728 22202 9856
rect 800 9448 22120 9728
rect 800 9320 22202 9448
rect 800 9040 22120 9320
rect 800 8912 22202 9040
rect 800 8632 22120 8912
rect 800 8504 22202 8632
rect 800 8224 22120 8504
rect 800 8096 22202 8224
rect 800 7816 22120 8096
rect 800 7688 22202 7816
rect 800 7408 22120 7688
rect 800 7280 22202 7408
rect 800 7000 22120 7280
rect 800 6872 22202 7000
rect 800 6592 22120 6872
rect 800 6464 22202 6592
rect 800 6184 22120 6464
rect 800 6056 22202 6184
rect 800 5920 22120 6056
rect 880 5776 22120 5920
rect 880 5648 22202 5776
rect 880 5640 22120 5648
rect 800 5368 22120 5640
rect 800 5240 22202 5368
rect 800 4960 22120 5240
rect 800 4832 22202 4960
rect 800 4552 22120 4832
rect 800 4424 22202 4552
rect 800 4144 22120 4424
rect 800 4016 22202 4144
rect 800 3736 22120 4016
rect 800 3608 22202 3736
rect 800 3328 22120 3608
rect 800 3200 22202 3328
rect 800 2920 22120 3200
rect 800 2792 22202 2920
rect 800 2512 22120 2792
rect 800 2384 22202 2512
rect 800 2104 22120 2384
rect 800 1976 22202 2104
rect 800 1696 22120 1976
rect 800 1568 22202 1696
rect 800 1395 22120 1568
<< metal4 >>
rect 3543 2128 3863 20720
rect 6142 2128 6462 20720
rect 8741 2128 9061 20720
rect 11340 2128 11660 20720
rect 13939 2128 14259 20720
rect 16538 2128 16858 20720
rect 19137 2128 19457 20720
rect 21736 2128 22056 20720
<< obsm4 >>
rect 19563 13227 19629 18053
<< labels >>
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 21736 2128 22056 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 5720 800 5840 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 ccff_tail
port 4 nsew signal output
rlabel metal3 s 22200 5040 23000 5160 6 chanx_right_in[0]
port 5 nsew signal input
rlabel metal3 s 22200 9120 23000 9240 6 chanx_right_in[10]
port 6 nsew signal input
rlabel metal3 s 22200 9528 23000 9648 6 chanx_right_in[11]
port 7 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[12]
port 8 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[13]
port 9 nsew signal input
rlabel metal3 s 22200 10752 23000 10872 6 chanx_right_in[14]
port 10 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[15]
port 11 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[16]
port 12 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_in[17]
port 13 nsew signal input
rlabel metal3 s 22200 12384 23000 12504 6 chanx_right_in[18]
port 14 nsew signal input
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_in[19]
port 15 nsew signal input
rlabel metal3 s 22200 5448 23000 5568 6 chanx_right_in[1]
port 16 nsew signal input
rlabel metal3 s 22200 5856 23000 5976 6 chanx_right_in[2]
port 17 nsew signal input
rlabel metal3 s 22200 6264 23000 6384 6 chanx_right_in[3]
port 18 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[4]
port 19 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[5]
port 20 nsew signal input
rlabel metal3 s 22200 7488 23000 7608 6 chanx_right_in[6]
port 21 nsew signal input
rlabel metal3 s 22200 7896 23000 8016 6 chanx_right_in[7]
port 22 nsew signal input
rlabel metal3 s 22200 8304 23000 8424 6 chanx_right_in[8]
port 23 nsew signal input
rlabel metal3 s 22200 8712 23000 8832 6 chanx_right_in[9]
port 24 nsew signal input
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_out[0]
port 25 nsew signal output
rlabel metal3 s 22200 17280 23000 17400 6 chanx_right_out[10]
port 26 nsew signal output
rlabel metal3 s 22200 17688 23000 17808 6 chanx_right_out[11]
port 27 nsew signal output
rlabel metal3 s 22200 18096 23000 18216 6 chanx_right_out[12]
port 28 nsew signal output
rlabel metal3 s 22200 18504 23000 18624 6 chanx_right_out[13]
port 29 nsew signal output
rlabel metal3 s 22200 18912 23000 19032 6 chanx_right_out[14]
port 30 nsew signal output
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[15]
port 31 nsew signal output
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[16]
port 32 nsew signal output
rlabel metal3 s 22200 20136 23000 20256 6 chanx_right_out[17]
port 33 nsew signal output
rlabel metal3 s 22200 20544 23000 20664 6 chanx_right_out[18]
port 34 nsew signal output
rlabel metal3 s 22200 20952 23000 21072 6 chanx_right_out[19]
port 35 nsew signal output
rlabel metal3 s 22200 13608 23000 13728 6 chanx_right_out[1]
port 36 nsew signal output
rlabel metal3 s 22200 14016 23000 14136 6 chanx_right_out[2]
port 37 nsew signal output
rlabel metal3 s 22200 14424 23000 14544 6 chanx_right_out[3]
port 38 nsew signal output
rlabel metal3 s 22200 14832 23000 14952 6 chanx_right_out[4]
port 39 nsew signal output
rlabel metal3 s 22200 15240 23000 15360 6 chanx_right_out[5]
port 40 nsew signal output
rlabel metal3 s 22200 15648 23000 15768 6 chanx_right_out[6]
port 41 nsew signal output
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[7]
port 42 nsew signal output
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[8]
port 43 nsew signal output
rlabel metal3 s 22200 16872 23000 16992 6 chanx_right_out[9]
port 44 nsew signal output
rlabel metal2 s 938 22200 994 23000 6 chany_top_in[0]
port 45 nsew signal input
rlabel metal2 s 6458 22200 6514 23000 6 chany_top_in[10]
port 46 nsew signal input
rlabel metal2 s 7010 22200 7066 23000 6 chany_top_in[11]
port 47 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[12]
port 48 nsew signal input
rlabel metal2 s 8114 22200 8170 23000 6 chany_top_in[13]
port 49 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[14]
port 50 nsew signal input
rlabel metal2 s 9218 22200 9274 23000 6 chany_top_in[15]
port 51 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[16]
port 52 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[17]
port 53 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_in[18]
port 54 nsew signal input
rlabel metal2 s 11426 22200 11482 23000 6 chany_top_in[19]
port 55 nsew signal input
rlabel metal2 s 1490 22200 1546 23000 6 chany_top_in[1]
port 56 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 chany_top_in[2]
port 57 nsew signal input
rlabel metal2 s 2594 22200 2650 23000 6 chany_top_in[3]
port 58 nsew signal input
rlabel metal2 s 3146 22200 3202 23000 6 chany_top_in[4]
port 59 nsew signal input
rlabel metal2 s 3698 22200 3754 23000 6 chany_top_in[5]
port 60 nsew signal input
rlabel metal2 s 4250 22200 4306 23000 6 chany_top_in[6]
port 61 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[7]
port 62 nsew signal input
rlabel metal2 s 5354 22200 5410 23000 6 chany_top_in[8]
port 63 nsew signal input
rlabel metal2 s 5906 22200 5962 23000 6 chany_top_in[9]
port 64 nsew signal input
rlabel metal2 s 11978 22200 12034 23000 6 chany_top_out[0]
port 65 nsew signal output
rlabel metal2 s 17498 22200 17554 23000 6 chany_top_out[10]
port 66 nsew signal output
rlabel metal2 s 18050 22200 18106 23000 6 chany_top_out[11]
port 67 nsew signal output
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[12]
port 68 nsew signal output
rlabel metal2 s 19154 22200 19210 23000 6 chany_top_out[13]
port 69 nsew signal output
rlabel metal2 s 19706 22200 19762 23000 6 chany_top_out[14]
port 70 nsew signal output
rlabel metal2 s 20258 22200 20314 23000 6 chany_top_out[15]
port 71 nsew signal output
rlabel metal2 s 20810 22200 20866 23000 6 chany_top_out[16]
port 72 nsew signal output
rlabel metal2 s 21362 22200 21418 23000 6 chany_top_out[17]
port 73 nsew signal output
rlabel metal2 s 21914 22200 21970 23000 6 chany_top_out[18]
port 74 nsew signal output
rlabel metal2 s 22466 22200 22522 23000 6 chany_top_out[19]
port 75 nsew signal output
rlabel metal2 s 12530 22200 12586 23000 6 chany_top_out[1]
port 76 nsew signal output
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[2]
port 77 nsew signal output
rlabel metal2 s 13634 22200 13690 23000 6 chany_top_out[3]
port 78 nsew signal output
rlabel metal2 s 14186 22200 14242 23000 6 chany_top_out[4]
port 79 nsew signal output
rlabel metal2 s 14738 22200 14794 23000 6 chany_top_out[5]
port 80 nsew signal output
rlabel metal2 s 15290 22200 15346 23000 6 chany_top_out[6]
port 81 nsew signal output
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[7]
port 82 nsew signal output
rlabel metal2 s 16394 22200 16450 23000 6 chany_top_out[8]
port 83 nsew signal output
rlabel metal2 s 16946 22200 17002 23000 6 chany_top_out[9]
port 84 nsew signal output
rlabel metal3 s 22200 21360 23000 21480 6 prog_clk_0_E_in
port 85 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_11_
port 86 nsew signal input
rlabel metal3 s 22200 3816 23000 3936 6 right_bottom_grid_pin_13_
port 87 nsew signal input
rlabel metal3 s 22200 4224 23000 4344 6 right_bottom_grid_pin_15_
port 88 nsew signal input
rlabel metal3 s 22200 4632 23000 4752 6 right_bottom_grid_pin_17_
port 89 nsew signal input
rlabel metal3 s 22200 1368 23000 1488 6 right_bottom_grid_pin_1_
port 90 nsew signal input
rlabel metal3 s 22200 1776 23000 1896 6 right_bottom_grid_pin_3_
port 91 nsew signal input
rlabel metal3 s 22200 2184 23000 2304 6 right_bottom_grid_pin_5_
port 92 nsew signal input
rlabel metal3 s 22200 2592 23000 2712 6 right_bottom_grid_pin_7_
port 93 nsew signal input
rlabel metal3 s 22200 3000 23000 3120 6 right_bottom_grid_pin_9_
port 94 nsew signal input
rlabel metal2 s 386 22200 442 23000 6 top_left_grid_pin_1_
port 95 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 813060
string GDS_FILE /home/marwan/clear_signoff_final/openlane/sb_0__0_/runs/sb_0__0_/results/signoff/sb_0__0_.magic.gds
string GDS_START 65026
<< end >>

