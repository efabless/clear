magic
tech sky130A
magscale 1 2
timestamp 1656942943
<< viali >>
rect 4353 14025 4387 14059
rect 4537 13889 4571 13923
rect 4905 13889 4939 13923
rect 5089 13821 5123 13855
rect 4169 12937 4203 12971
rect 5917 12937 5951 12971
rect 14473 12937 14507 12971
rect 4598 12869 4632 12903
rect 6101 12801 6135 12835
rect 14289 12801 14323 12835
rect 4353 12733 4387 12767
rect 5733 12597 5767 12631
rect 6469 12597 6503 12631
rect 14197 12597 14231 12631
rect 4629 12393 4663 12427
rect 7481 12393 7515 12427
rect 9413 12393 9447 12427
rect 5181 12325 5215 12359
rect 4813 12189 4847 12223
rect 5365 12189 5399 12223
rect 7665 12189 7699 12223
rect 9597 12189 9631 12223
rect 5549 12121 5583 12155
rect 4997 12053 5031 12087
rect 7757 12053 7791 12087
rect 7941 12053 7975 12087
rect 9781 12053 9815 12087
rect 7297 11849 7331 11883
rect 7665 11849 7699 11883
rect 8769 11849 8803 11883
rect 9045 11781 9079 11815
rect 7113 11713 7147 11747
rect 7481 11713 7515 11747
rect 7849 11713 7883 11747
rect 8309 11713 8343 11747
rect 8953 11713 8987 11747
rect 8585 11645 8619 11679
rect 8125 11509 8159 11543
rect 6469 11305 6503 11339
rect 6929 11305 6963 11339
rect 8769 11305 8803 11339
rect 7205 11237 7239 11271
rect 8953 11237 8987 11271
rect 7757 11169 7791 11203
rect 8125 11169 8159 11203
rect 9505 11169 9539 11203
rect 9873 11169 9907 11203
rect 6745 11101 6779 11135
rect 7113 11101 7147 11135
rect 7573 11101 7607 11135
rect 8401 11101 8435 11135
rect 9321 11101 9355 11135
rect 9413 11101 9447 11135
rect 7665 11033 7699 11067
rect 6009 10965 6043 10999
rect 6285 10965 6319 10999
rect 8309 10965 8343 10999
rect 5365 10761 5399 10795
rect 6009 10761 6043 10795
rect 7297 10761 7331 10795
rect 9137 10761 9171 10795
rect 10241 10761 10275 10795
rect 11621 10761 11655 10795
rect 5181 10693 5215 10727
rect 12265 10693 12299 10727
rect 3468 10625 3502 10659
rect 5825 10625 5859 10659
rect 6193 10625 6227 10659
rect 6837 10625 6871 10659
rect 8024 10625 8058 10659
rect 9505 10625 9539 10659
rect 9873 10625 9907 10659
rect 11161 10625 11195 10659
rect 7021 10557 7055 10591
rect 7205 10557 7239 10591
rect 7757 10557 7791 10591
rect 10057 10557 10091 10591
rect 11897 10557 11931 10591
rect 5641 10489 5675 10523
rect 9321 10489 9355 10523
rect 10425 10489 10459 10523
rect 3571 10421 3605 10455
rect 6377 10421 6411 10455
rect 6653 10421 6687 10455
rect 7665 10421 7699 10455
rect 9689 10421 9723 10455
rect 10609 10421 10643 10455
rect 9045 10217 9079 10251
rect 12265 10217 12299 10251
rect 13001 10217 13035 10251
rect 13553 10217 13587 10251
rect 5089 10149 5123 10183
rect 8585 10149 8619 10183
rect 11529 10149 11563 10183
rect 13737 10149 13771 10183
rect 5733 10081 5767 10115
rect 8677 10081 8711 10115
rect 9597 10081 9631 10115
rect 10333 10081 10367 10115
rect 10425 10081 10459 10115
rect 4997 10013 5031 10047
rect 5457 10013 5491 10047
rect 7205 10013 7239 10047
rect 9413 10013 9447 10047
rect 10241 10013 10275 10047
rect 10977 10013 11011 10047
rect 11345 10013 11379 10047
rect 11713 10013 11747 10047
rect 12081 10013 12115 10047
rect 12449 10013 12483 10047
rect 12817 10013 12851 10047
rect 13185 10013 13219 10047
rect 6009 9945 6043 9979
rect 6101 9945 6135 9979
rect 7021 9945 7055 9979
rect 7472 9945 7506 9979
rect 4813 9877 4847 9911
rect 5549 9877 5583 9911
rect 9505 9877 9539 9911
rect 9873 9877 9907 9911
rect 10793 9877 10827 9911
rect 11161 9877 11195 9911
rect 11897 9877 11931 9911
rect 12633 9877 12667 9911
rect 13369 9877 13403 9911
rect 6653 9673 6687 9707
rect 1593 9605 1627 9639
rect 8064 9605 8098 9639
rect 8861 9605 8895 9639
rect 11253 9605 11287 9639
rect 5457 9537 5491 9571
rect 5825 9537 5859 9571
rect 6193 9537 6227 9571
rect 6469 9537 6503 9571
rect 6837 9537 6871 9571
rect 8769 9537 8803 9571
rect 9505 9537 9539 9571
rect 9873 9537 9907 9571
rect 10333 9537 10367 9571
rect 10701 9537 10735 9571
rect 11069 9537 11103 9571
rect 12265 9537 12299 9571
rect 12633 9537 12667 9571
rect 1501 9469 1535 9503
rect 1777 9469 1811 9503
rect 8302 9469 8336 9503
rect 9045 9469 9079 9503
rect 6009 9401 6043 9435
rect 8401 9401 8435 9435
rect 9321 9401 9355 9435
rect 10885 9401 10919 9435
rect 12081 9401 12115 9435
rect 12449 9401 12483 9435
rect 12817 9401 12851 9435
rect 5273 9333 5307 9367
rect 5641 9333 5675 9367
rect 6929 9333 6963 9367
rect 9689 9333 9723 9367
rect 10149 9333 10183 9367
rect 10517 9333 10551 9367
rect 11621 9333 11655 9367
rect 11805 9333 11839 9367
rect 13001 9333 13035 9367
rect 6009 9129 6043 9163
rect 8217 9129 8251 9163
rect 9413 9129 9447 9163
rect 10149 9129 10183 9163
rect 6837 8993 6871 9027
rect 9689 8993 9723 9027
rect 6377 8925 6411 8959
rect 7104 8925 7138 8959
rect 8677 8925 8711 8959
rect 9229 8925 9263 8959
rect 9873 8857 9907 8891
rect 1501 8789 1535 8823
rect 5641 8789 5675 8823
rect 8493 8789 8527 8823
rect 9045 8789 9079 8823
rect 10057 8789 10091 8823
rect 7113 8585 7147 8619
rect 7481 8585 7515 8619
rect 8033 8585 8067 8619
rect 8493 8585 8527 8619
rect 8953 8585 8987 8619
rect 11713 8517 11747 8551
rect 7573 8449 7607 8483
rect 8401 8449 8435 8483
rect 12541 8449 12575 8483
rect 7665 8381 7699 8415
rect 8677 8381 8711 8415
rect 12725 8313 12759 8347
rect 9137 8245 9171 8279
rect 5733 7497 5767 7531
rect 7849 7497 7883 7531
rect 9597 7497 9631 7531
rect 4997 7429 5031 7463
rect 5457 7429 5491 7463
rect 3525 7361 3559 7395
rect 4813 7361 4847 7395
rect 5365 7361 5399 7395
rect 5917 7361 5951 7395
rect 7665 7361 7699 7395
rect 9505 7361 9539 7395
rect 3249 7293 3283 7327
rect 6101 7293 6135 7327
rect 9321 7225 9355 7259
rect 4629 7157 4663 7191
rect 5181 7157 5215 7191
rect 7481 7157 7515 7191
<< metal1 >>
rect 4154 17892 4160 17944
rect 4212 17932 4218 17944
rect 4338 17932 4344 17944
rect 4212 17904 4344 17932
rect 4212 17892 4218 17904
rect 4338 17892 4344 17904
rect 4396 17892 4402 17944
rect 1104 17434 16008 17456
rect 1104 17382 4698 17434
rect 4750 17382 4762 17434
rect 4814 17382 4826 17434
rect 4878 17382 4890 17434
rect 4942 17382 4954 17434
rect 5006 17382 8446 17434
rect 8498 17382 8510 17434
rect 8562 17382 8574 17434
rect 8626 17382 8638 17434
rect 8690 17382 8702 17434
rect 8754 17382 12194 17434
rect 12246 17382 12258 17434
rect 12310 17382 12322 17434
rect 12374 17382 12386 17434
rect 12438 17382 12450 17434
rect 12502 17382 16008 17434
rect 1104 17360 16008 17382
rect 1104 16890 16008 16912
rect 1104 16838 2824 16890
rect 2876 16838 2888 16890
rect 2940 16838 2952 16890
rect 3004 16838 3016 16890
rect 3068 16838 3080 16890
rect 3132 16838 6572 16890
rect 6624 16838 6636 16890
rect 6688 16838 6700 16890
rect 6752 16838 6764 16890
rect 6816 16838 6828 16890
rect 6880 16838 10320 16890
rect 10372 16838 10384 16890
rect 10436 16838 10448 16890
rect 10500 16838 10512 16890
rect 10564 16838 10576 16890
rect 10628 16838 14068 16890
rect 14120 16838 14132 16890
rect 14184 16838 14196 16890
rect 14248 16838 14260 16890
rect 14312 16838 14324 16890
rect 14376 16838 16008 16890
rect 1104 16816 16008 16838
rect 5718 16532 5724 16584
rect 5776 16572 5782 16584
rect 6086 16572 6092 16584
rect 5776 16544 6092 16572
rect 5776 16532 5782 16544
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 1104 16346 16008 16368
rect 1104 16294 4698 16346
rect 4750 16294 4762 16346
rect 4814 16294 4826 16346
rect 4878 16294 4890 16346
rect 4942 16294 4954 16346
rect 5006 16294 8446 16346
rect 8498 16294 8510 16346
rect 8562 16294 8574 16346
rect 8626 16294 8638 16346
rect 8690 16294 8702 16346
rect 8754 16294 12194 16346
rect 12246 16294 12258 16346
rect 12310 16294 12322 16346
rect 12374 16294 12386 16346
rect 12438 16294 12450 16346
rect 12502 16294 16008 16346
rect 1104 16272 16008 16294
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 6454 16096 6460 16108
rect 5776 16068 6460 16096
rect 5776 16056 5782 16068
rect 6454 16056 6460 16068
rect 6512 16056 6518 16108
rect 3786 15988 3792 16040
rect 3844 16028 3850 16040
rect 5350 16028 5356 16040
rect 3844 16000 5356 16028
rect 3844 15988 3850 16000
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 6454 15920 6460 15972
rect 6512 15960 6518 15972
rect 11514 15960 11520 15972
rect 6512 15932 11520 15960
rect 6512 15920 6518 15932
rect 11514 15920 11520 15932
rect 11572 15920 11578 15972
rect 7190 15852 7196 15904
rect 7248 15892 7254 15904
rect 10778 15892 10784 15904
rect 7248 15864 10784 15892
rect 7248 15852 7254 15864
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 1104 15802 16008 15824
rect 1104 15750 2824 15802
rect 2876 15750 2888 15802
rect 2940 15750 2952 15802
rect 3004 15750 3016 15802
rect 3068 15750 3080 15802
rect 3132 15750 6572 15802
rect 6624 15750 6636 15802
rect 6688 15750 6700 15802
rect 6752 15750 6764 15802
rect 6816 15750 6828 15802
rect 6880 15750 10320 15802
rect 10372 15750 10384 15802
rect 10436 15750 10448 15802
rect 10500 15750 10512 15802
rect 10564 15750 10576 15802
rect 10628 15750 14068 15802
rect 14120 15750 14132 15802
rect 14184 15750 14196 15802
rect 14248 15750 14260 15802
rect 14312 15750 14324 15802
rect 14376 15750 16008 15802
rect 1104 15728 16008 15750
rect 7098 15648 7104 15700
rect 7156 15688 7162 15700
rect 9674 15688 9680 15700
rect 7156 15660 9680 15688
rect 7156 15648 7162 15660
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 11146 15648 11152 15700
rect 11204 15688 11210 15700
rect 14826 15688 14832 15700
rect 11204 15660 14832 15688
rect 11204 15648 11210 15660
rect 14826 15648 14832 15660
rect 14884 15648 14890 15700
rect 4338 15580 4344 15632
rect 4396 15620 4402 15632
rect 7650 15620 7656 15632
rect 4396 15592 7656 15620
rect 4396 15580 4402 15592
rect 7650 15580 7656 15592
rect 7708 15580 7714 15632
rect 8202 15580 8208 15632
rect 8260 15620 8266 15632
rect 11974 15620 11980 15632
rect 8260 15592 11980 15620
rect 8260 15580 8266 15592
rect 11974 15580 11980 15592
rect 12032 15580 12038 15632
rect 3418 15512 3424 15564
rect 3476 15552 3482 15564
rect 5810 15552 5816 15564
rect 3476 15524 5816 15552
rect 3476 15512 3482 15524
rect 5810 15512 5816 15524
rect 5868 15512 5874 15564
rect 8846 15512 8852 15564
rect 8904 15552 8910 15564
rect 12618 15552 12624 15564
rect 8904 15524 12624 15552
rect 8904 15512 8910 15524
rect 12618 15512 12624 15524
rect 12676 15512 12682 15564
rect 2314 15444 2320 15496
rect 2372 15484 2378 15496
rect 3970 15484 3976 15496
rect 2372 15456 3976 15484
rect 2372 15444 2378 15456
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 7466 15444 7472 15496
rect 7524 15484 7530 15496
rect 9398 15484 9404 15496
rect 7524 15456 9404 15484
rect 7524 15444 7530 15456
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 10134 15444 10140 15496
rect 10192 15484 10198 15496
rect 12066 15484 12072 15496
rect 10192 15456 12072 15484
rect 10192 15444 10198 15456
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 3142 15376 3148 15428
rect 3200 15416 3206 15428
rect 5902 15416 5908 15428
rect 3200 15388 5908 15416
rect 3200 15376 3206 15388
rect 5902 15376 5908 15388
rect 5960 15376 5966 15428
rect 7834 15376 7840 15428
rect 7892 15416 7898 15428
rect 10778 15416 10784 15428
rect 7892 15388 10784 15416
rect 7892 15376 7898 15388
rect 10778 15376 10784 15388
rect 10836 15376 10842 15428
rect 11054 15376 11060 15428
rect 11112 15416 11118 15428
rect 12986 15416 12992 15428
rect 11112 15388 12992 15416
rect 11112 15376 11118 15388
rect 12986 15376 12992 15388
rect 13044 15376 13050 15428
rect 13814 15376 13820 15428
rect 13872 15416 13878 15428
rect 15562 15416 15568 15428
rect 13872 15388 15568 15416
rect 13872 15376 13878 15388
rect 15562 15376 15568 15388
rect 15620 15376 15626 15428
rect 1578 15308 1584 15360
rect 1636 15348 1642 15360
rect 4062 15348 4068 15360
rect 1636 15320 4068 15348
rect 1636 15308 1642 15320
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 5258 15308 5264 15360
rect 5316 15348 5322 15360
rect 7466 15348 7472 15360
rect 5316 15320 7472 15348
rect 5316 15308 5322 15320
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 9030 15308 9036 15360
rect 9088 15348 9094 15360
rect 10226 15348 10232 15360
rect 9088 15320 10232 15348
rect 9088 15308 9094 15320
rect 10226 15308 10232 15320
rect 10284 15308 10290 15360
rect 10686 15308 10692 15360
rect 10744 15348 10750 15360
rect 13354 15348 13360 15360
rect 10744 15320 13360 15348
rect 10744 15308 10750 15320
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 14458 15308 14464 15360
rect 14516 15348 14522 15360
rect 15930 15348 15936 15360
rect 14516 15320 15936 15348
rect 14516 15308 14522 15320
rect 15930 15308 15936 15320
rect 15988 15308 15994 15360
rect 1104 15258 16008 15280
rect 1104 15206 4698 15258
rect 4750 15206 4762 15258
rect 4814 15206 4826 15258
rect 4878 15206 4890 15258
rect 4942 15206 4954 15258
rect 5006 15206 8446 15258
rect 8498 15206 8510 15258
rect 8562 15206 8574 15258
rect 8626 15206 8638 15258
rect 8690 15206 8702 15258
rect 8754 15206 12194 15258
rect 12246 15206 12258 15258
rect 12310 15206 12322 15258
rect 12374 15206 12386 15258
rect 12438 15206 12450 15258
rect 12502 15206 16008 15258
rect 1104 15184 16008 15206
rect 1104 14714 16008 14736
rect 1104 14662 2824 14714
rect 2876 14662 2888 14714
rect 2940 14662 2952 14714
rect 3004 14662 3016 14714
rect 3068 14662 3080 14714
rect 3132 14662 6572 14714
rect 6624 14662 6636 14714
rect 6688 14662 6700 14714
rect 6752 14662 6764 14714
rect 6816 14662 6828 14714
rect 6880 14662 10320 14714
rect 10372 14662 10384 14714
rect 10436 14662 10448 14714
rect 10500 14662 10512 14714
rect 10564 14662 10576 14714
rect 10628 14662 14068 14714
rect 14120 14662 14132 14714
rect 14184 14662 14196 14714
rect 14248 14662 14260 14714
rect 14312 14662 14324 14714
rect 14376 14662 16008 14714
rect 1104 14640 16008 14662
rect 1104 14170 16008 14192
rect 1104 14118 4698 14170
rect 4750 14118 4762 14170
rect 4814 14118 4826 14170
rect 4878 14118 4890 14170
rect 4942 14118 4954 14170
rect 5006 14118 8446 14170
rect 8498 14118 8510 14170
rect 8562 14118 8574 14170
rect 8626 14118 8638 14170
rect 8690 14118 8702 14170
rect 8754 14118 12194 14170
rect 12246 14118 12258 14170
rect 12310 14118 12322 14170
rect 12374 14118 12386 14170
rect 12438 14118 12450 14170
rect 12502 14118 16008 14170
rect 1104 14096 16008 14118
rect 1210 14016 1216 14068
rect 1268 14056 1274 14068
rect 4341 14059 4399 14065
rect 4341 14056 4353 14059
rect 1268 14028 4353 14056
rect 1268 14016 1274 14028
rect 4341 14025 4353 14028
rect 4387 14056 4399 14059
rect 4387 14028 4568 14056
rect 4387 14025 4399 14028
rect 4341 14019 4399 14025
rect 4540 13929 4568 14028
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13889 4583 13923
rect 4525 13883 4583 13889
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13920 4951 13923
rect 9582 13920 9588 13932
rect 4939 13892 9588 13920
rect 4939 13889 4951 13892
rect 4893 13883 4951 13889
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 3510 13812 3516 13864
rect 3568 13852 3574 13864
rect 5077 13855 5135 13861
rect 5077 13852 5089 13855
rect 3568 13824 5089 13852
rect 3568 13812 3574 13824
rect 5077 13821 5089 13824
rect 5123 13821 5135 13855
rect 5077 13815 5135 13821
rect 1104 13626 16008 13648
rect 1104 13574 2824 13626
rect 2876 13574 2888 13626
rect 2940 13574 2952 13626
rect 3004 13574 3016 13626
rect 3068 13574 3080 13626
rect 3132 13574 6572 13626
rect 6624 13574 6636 13626
rect 6688 13574 6700 13626
rect 6752 13574 6764 13626
rect 6816 13574 6828 13626
rect 6880 13574 10320 13626
rect 10372 13574 10384 13626
rect 10436 13574 10448 13626
rect 10500 13574 10512 13626
rect 10564 13574 10576 13626
rect 10628 13574 14068 13626
rect 14120 13574 14132 13626
rect 14184 13574 14196 13626
rect 14248 13574 14260 13626
rect 14312 13574 14324 13626
rect 14376 13574 16008 13626
rect 1104 13552 16008 13574
rect 1104 13082 16008 13104
rect 1104 13030 4698 13082
rect 4750 13030 4762 13082
rect 4814 13030 4826 13082
rect 4878 13030 4890 13082
rect 4942 13030 4954 13082
rect 5006 13030 8446 13082
rect 8498 13030 8510 13082
rect 8562 13030 8574 13082
rect 8626 13030 8638 13082
rect 8690 13030 8702 13082
rect 8754 13030 12194 13082
rect 12246 13030 12258 13082
rect 12310 13030 12322 13082
rect 12374 13030 12386 13082
rect 12438 13030 12450 13082
rect 12502 13030 16008 13082
rect 1104 13008 16008 13030
rect 4154 12968 4160 12980
rect 4115 12940 4160 12968
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 5902 12968 5908 12980
rect 5863 12940 5908 12968
rect 5902 12928 5908 12940
rect 5960 12928 5966 12980
rect 13722 12928 13728 12980
rect 13780 12968 13786 12980
rect 14461 12971 14519 12977
rect 14461 12968 14473 12971
rect 13780 12940 14473 12968
rect 13780 12928 13786 12940
rect 14461 12937 14473 12940
rect 14507 12937 14519 12971
rect 14461 12931 14519 12937
rect 4172 12900 4200 12928
rect 4586 12903 4644 12909
rect 4586 12900 4598 12903
rect 4172 12872 4598 12900
rect 4586 12869 4598 12872
rect 4632 12869 4644 12903
rect 4586 12863 4644 12869
rect 6089 12835 6147 12841
rect 6089 12801 6101 12835
rect 6135 12832 6147 12835
rect 14277 12835 14335 12841
rect 6135 12804 6500 12832
rect 6135 12801 6147 12804
rect 6089 12795 6147 12801
rect 4338 12764 4344 12776
rect 4299 12736 4344 12764
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 5721 12631 5779 12637
rect 5721 12597 5733 12631
rect 5767 12628 5779 12631
rect 6362 12628 6368 12640
rect 5767 12600 6368 12628
rect 5767 12597 5779 12600
rect 5721 12591 5779 12597
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 6472 12637 6500 12804
rect 14277 12801 14289 12835
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 6457 12631 6515 12637
rect 6457 12597 6469 12631
rect 6503 12628 6515 12631
rect 8202 12628 8208 12640
rect 6503 12600 8208 12628
rect 6503 12597 6515 12600
rect 6457 12591 6515 12597
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 9582 12588 9588 12640
rect 9640 12628 9646 12640
rect 12434 12628 12440 12640
rect 9640 12600 12440 12628
rect 9640 12588 9646 12600
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 14185 12631 14243 12637
rect 14185 12597 14197 12631
rect 14231 12628 14243 12631
rect 14292 12628 14320 12795
rect 14642 12628 14648 12640
rect 14231 12600 14648 12628
rect 14231 12597 14243 12600
rect 14185 12591 14243 12597
rect 14642 12588 14648 12600
rect 14700 12588 14706 12640
rect 1104 12538 16008 12560
rect 1104 12486 2824 12538
rect 2876 12486 2888 12538
rect 2940 12486 2952 12538
rect 3004 12486 3016 12538
rect 3068 12486 3080 12538
rect 3132 12486 6572 12538
rect 6624 12486 6636 12538
rect 6688 12486 6700 12538
rect 6752 12486 6764 12538
rect 6816 12486 6828 12538
rect 6880 12486 10320 12538
rect 10372 12486 10384 12538
rect 10436 12486 10448 12538
rect 10500 12486 10512 12538
rect 10564 12486 10576 12538
rect 10628 12486 14068 12538
rect 14120 12486 14132 12538
rect 14184 12486 14196 12538
rect 14248 12486 14260 12538
rect 14312 12486 14324 12538
rect 14376 12486 16008 12538
rect 1104 12464 16008 12486
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 4617 12427 4675 12433
rect 4617 12424 4629 12427
rect 4120 12396 4629 12424
rect 4120 12384 4126 12396
rect 4617 12393 4629 12396
rect 4663 12393 4675 12427
rect 7466 12424 7472 12436
rect 7427 12396 7472 12424
rect 4617 12387 4675 12393
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8938 12424 8944 12436
rect 8352 12396 8944 12424
rect 8352 12384 8358 12396
rect 8938 12384 8944 12396
rect 8996 12384 9002 12436
rect 9398 12424 9404 12436
rect 9359 12396 9404 12424
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 3970 12316 3976 12368
rect 4028 12356 4034 12368
rect 5169 12359 5227 12365
rect 5169 12356 5181 12359
rect 4028 12328 5181 12356
rect 4028 12316 4034 12328
rect 5169 12325 5181 12328
rect 5215 12325 5227 12359
rect 5169 12319 5227 12325
rect 7190 12316 7196 12368
rect 7248 12356 7254 12368
rect 10962 12356 10968 12368
rect 7248 12328 10968 12356
rect 7248 12316 7254 12328
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 9766 12248 9772 12300
rect 9824 12288 9830 12300
rect 9950 12288 9956 12300
rect 9824 12260 9956 12288
rect 9824 12248 9830 12260
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12220 4859 12223
rect 5353 12223 5411 12229
rect 4847 12192 5028 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 5000 12093 5028 12192
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 7653 12223 7711 12229
rect 5399 12192 5580 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 5552 12161 5580 12192
rect 7653 12189 7665 12223
rect 7699 12220 7711 12223
rect 7742 12220 7748 12232
rect 7699 12192 7748 12220
rect 7699 12189 7711 12192
rect 7653 12183 7711 12189
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12220 9643 12223
rect 9631 12192 9812 12220
rect 9631 12189 9643 12192
rect 9585 12183 9643 12189
rect 5537 12155 5595 12161
rect 5537 12121 5549 12155
rect 5583 12152 5595 12155
rect 9122 12152 9128 12164
rect 5583 12124 9128 12152
rect 5583 12121 5595 12124
rect 5537 12115 5595 12121
rect 9122 12112 9128 12124
rect 9180 12112 9186 12164
rect 9784 12096 9812 12192
rect 4985 12087 5043 12093
rect 4985 12053 4997 12087
rect 5031 12084 5043 12087
rect 5902 12084 5908 12096
rect 5031 12056 5908 12084
rect 5031 12053 5043 12056
rect 4985 12047 5043 12053
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 7742 12084 7748 12096
rect 7703 12056 7748 12084
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 7926 12084 7932 12096
rect 7887 12056 7932 12084
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 9766 12084 9772 12096
rect 9727 12056 9772 12084
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 1104 11994 16008 12016
rect 1104 11942 4698 11994
rect 4750 11942 4762 11994
rect 4814 11942 4826 11994
rect 4878 11942 4890 11994
rect 4942 11942 4954 11994
rect 5006 11942 8446 11994
rect 8498 11942 8510 11994
rect 8562 11942 8574 11994
rect 8626 11942 8638 11994
rect 8690 11942 8702 11994
rect 8754 11942 12194 11994
rect 12246 11942 12258 11994
rect 12310 11942 12322 11994
rect 12374 11942 12386 11994
rect 12438 11942 12450 11994
rect 12502 11942 16008 11994
rect 1104 11920 16008 11942
rect 5350 11840 5356 11892
rect 5408 11880 5414 11892
rect 7285 11883 7343 11889
rect 7285 11880 7297 11883
rect 5408 11852 7297 11880
rect 5408 11840 5414 11852
rect 7285 11849 7297 11852
rect 7331 11849 7343 11883
rect 7650 11880 7656 11892
rect 7611 11852 7656 11880
rect 7285 11843 7343 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 8757 11883 8815 11889
rect 8757 11849 8769 11883
rect 8803 11880 8815 11883
rect 11882 11880 11888 11892
rect 8803 11852 11888 11880
rect 8803 11849 8815 11852
rect 8757 11843 8815 11849
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11744 7159 11747
rect 7469 11747 7527 11753
rect 7469 11744 7481 11747
rect 7147 11716 7481 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 7469 11713 7481 11716
rect 7515 11744 7527 11747
rect 7558 11744 7564 11756
rect 7515 11716 7564 11744
rect 7515 11713 7527 11716
rect 7469 11707 7527 11713
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 7837 11747 7895 11753
rect 7837 11713 7849 11747
rect 7883 11744 7895 11747
rect 7926 11744 7932 11756
rect 7883 11716 7932 11744
rect 7883 11713 7895 11716
rect 7837 11707 7895 11713
rect 7852 11608 7880 11707
rect 7926 11704 7932 11716
rect 7984 11704 7990 11756
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11744 8355 11747
rect 8772 11744 8800 11843
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 9033 11815 9091 11821
rect 9033 11781 9045 11815
rect 9079 11812 9091 11815
rect 9950 11812 9956 11824
rect 9079 11784 9956 11812
rect 9079 11781 9091 11784
rect 9033 11775 9091 11781
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 8343 11716 8800 11744
rect 8941 11747 8999 11753
rect 8343 11713 8355 11716
rect 8297 11707 8355 11713
rect 8941 11713 8953 11747
rect 8987 11744 8999 11747
rect 9122 11744 9128 11756
rect 8987 11716 9128 11744
rect 8987 11713 8999 11716
rect 8941 11707 8999 11713
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 9306 11676 9312 11688
rect 8619 11648 9312 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 11238 11608 11244 11620
rect 7852 11580 11244 11608
rect 11238 11568 11244 11580
rect 11296 11568 11302 11620
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 6178 11540 6184 11552
rect 5776 11512 6184 11540
rect 5776 11500 5782 11512
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 8110 11540 8116 11552
rect 8071 11512 8116 11540
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 1104 11450 16008 11472
rect 1104 11398 2824 11450
rect 2876 11398 2888 11450
rect 2940 11398 2952 11450
rect 3004 11398 3016 11450
rect 3068 11398 3080 11450
rect 3132 11398 6572 11450
rect 6624 11398 6636 11450
rect 6688 11398 6700 11450
rect 6752 11398 6764 11450
rect 6816 11398 6828 11450
rect 6880 11398 10320 11450
rect 10372 11398 10384 11450
rect 10436 11398 10448 11450
rect 10500 11398 10512 11450
rect 10564 11398 10576 11450
rect 10628 11398 14068 11450
rect 14120 11398 14132 11450
rect 14184 11398 14196 11450
rect 14248 11398 14260 11450
rect 14312 11398 14324 11450
rect 14376 11398 16008 11450
rect 1104 11376 16008 11398
rect 6454 11336 6460 11348
rect 6415 11308 6460 11336
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 6917 11339 6975 11345
rect 6917 11305 6929 11339
rect 6963 11336 6975 11339
rect 7006 11336 7012 11348
rect 6963 11308 7012 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 8757 11339 8815 11345
rect 8757 11305 8769 11339
rect 8803 11336 8815 11339
rect 10226 11336 10232 11348
rect 8803 11308 10232 11336
rect 8803 11305 8815 11308
rect 8757 11299 8815 11305
rect 10226 11296 10232 11308
rect 10284 11296 10290 11348
rect 5534 11228 5540 11280
rect 5592 11268 5598 11280
rect 7193 11271 7251 11277
rect 7193 11268 7205 11271
rect 5592 11240 7205 11268
rect 5592 11228 5598 11240
rect 7193 11237 7205 11240
rect 7239 11237 7251 11271
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 7193 11231 7251 11237
rect 7576 11240 8953 11268
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 6779 11104 7113 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 7101 11101 7113 11104
rect 7147 11132 7159 11135
rect 7190 11132 7196 11144
rect 7147 11104 7196 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7576 11141 7604 11240
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 9950 11268 9956 11280
rect 8941 11231 8999 11237
rect 9048 11240 9956 11268
rect 7650 11160 7656 11212
rect 7708 11200 7714 11212
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 7708 11172 7757 11200
rect 7708 11160 7714 11172
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 8113 11203 8171 11209
rect 8113 11200 8125 11203
rect 8076 11172 8125 11200
rect 8076 11160 8082 11172
rect 8113 11169 8125 11172
rect 8159 11169 8171 11203
rect 9048 11200 9076 11240
rect 9950 11228 9956 11240
rect 10008 11228 10014 11280
rect 9490 11200 9496 11212
rect 8113 11163 8171 11169
rect 8404 11172 9076 11200
rect 9451 11172 9496 11200
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 7834 11092 7840 11144
rect 7892 11132 7898 11144
rect 8404 11141 8432 11172
rect 9490 11160 9496 11172
rect 9548 11160 9554 11212
rect 9861 11203 9919 11209
rect 9861 11169 9873 11203
rect 9907 11200 9919 11203
rect 11146 11200 11152 11212
rect 9907 11172 11152 11200
rect 9907 11169 9919 11172
rect 9861 11163 9919 11169
rect 8389 11135 8447 11141
rect 8389 11132 8401 11135
rect 7892 11104 8401 11132
rect 7892 11092 7898 11104
rect 8389 11101 8401 11104
rect 8435 11101 8447 11135
rect 9306 11132 9312 11144
rect 9267 11104 9312 11132
rect 8389 11095 8447 11101
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 9876 11132 9904 11163
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 9456 11104 9904 11132
rect 9456 11092 9462 11104
rect 7653 11067 7711 11073
rect 7653 11033 7665 11067
rect 7699 11064 7711 11067
rect 9030 11064 9036 11076
rect 7699 11036 9036 11064
rect 7699 11033 7711 11036
rect 7653 11027 7711 11033
rect 9030 11024 9036 11036
rect 9088 11024 9094 11076
rect 9122 11024 9128 11076
rect 9180 11024 9186 11076
rect 5997 10999 6055 11005
rect 5997 10965 6009 10999
rect 6043 10996 6055 10999
rect 6086 10996 6092 11008
rect 6043 10968 6092 10996
rect 6043 10965 6055 10968
rect 5997 10959 6055 10965
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 6270 10996 6276 11008
rect 6231 10968 6276 10996
rect 6270 10956 6276 10968
rect 6328 10956 6334 11008
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 8018 10996 8024 11008
rect 7524 10968 8024 10996
rect 7524 10956 7530 10968
rect 8018 10956 8024 10968
rect 8076 10956 8082 11008
rect 8297 10999 8355 11005
rect 8297 10965 8309 10999
rect 8343 10996 8355 10999
rect 9140 10996 9168 11024
rect 8343 10968 9168 10996
rect 8343 10965 8355 10968
rect 8297 10959 8355 10965
rect 1104 10906 16008 10928
rect 1104 10854 4698 10906
rect 4750 10854 4762 10906
rect 4814 10854 4826 10906
rect 4878 10854 4890 10906
rect 4942 10854 4954 10906
rect 5006 10854 8446 10906
rect 8498 10854 8510 10906
rect 8562 10854 8574 10906
rect 8626 10854 8638 10906
rect 8690 10854 8702 10906
rect 8754 10854 12194 10906
rect 12246 10854 12258 10906
rect 12310 10854 12322 10906
rect 12374 10854 12386 10906
rect 12438 10854 12450 10906
rect 12502 10854 16008 10906
rect 1104 10832 16008 10854
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 5350 10792 5356 10804
rect 4212 10764 5356 10792
rect 4212 10752 4218 10764
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 5997 10795 6055 10801
rect 5997 10792 6009 10795
rect 5868 10764 6009 10792
rect 5868 10752 5874 10764
rect 5997 10761 6009 10764
rect 6043 10761 6055 10795
rect 7282 10792 7288 10804
rect 7195 10764 7288 10792
rect 5997 10755 6055 10761
rect 7282 10752 7288 10764
rect 7340 10792 7346 10804
rect 8294 10792 8300 10804
rect 7340 10764 8300 10792
rect 7340 10752 7346 10764
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 9582 10792 9588 10804
rect 9171 10764 9588 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 10229 10795 10287 10801
rect 10229 10761 10241 10795
rect 10275 10792 10287 10795
rect 10686 10792 10692 10804
rect 10275 10764 10692 10792
rect 10275 10761 10287 10764
rect 10229 10755 10287 10761
rect 4982 10684 4988 10736
rect 5040 10724 5046 10736
rect 5169 10727 5227 10733
rect 5169 10724 5181 10727
rect 5040 10696 5181 10724
rect 5040 10684 5046 10696
rect 5169 10693 5181 10696
rect 5215 10724 5227 10727
rect 9214 10724 9220 10736
rect 5215 10696 9220 10724
rect 5215 10693 5227 10696
rect 5169 10687 5227 10693
rect 9214 10684 9220 10696
rect 9272 10684 9278 10736
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 3510 10665 3516 10668
rect 3456 10659 3516 10665
rect 3456 10656 3468 10659
rect 3292 10628 3468 10656
rect 3292 10616 3298 10628
rect 3456 10625 3468 10628
rect 3502 10625 3516 10659
rect 3456 10619 3516 10625
rect 3510 10616 3516 10619
rect 3568 10656 3574 10668
rect 5813 10659 5871 10665
rect 3568 10628 3604 10656
rect 3568 10616 3574 10628
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 6086 10656 6092 10668
rect 5859 10628 6092 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 6086 10616 6092 10628
rect 6144 10616 6150 10668
rect 6181 10659 6239 10665
rect 6181 10625 6193 10659
rect 6227 10656 6239 10659
rect 6270 10656 6276 10668
rect 6227 10628 6276 10656
rect 6227 10625 6239 10628
rect 6181 10619 6239 10625
rect 6270 10616 6276 10628
rect 6328 10616 6334 10668
rect 6454 10616 6460 10668
rect 6512 10656 6518 10668
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6512 10628 6837 10656
rect 6512 10616 6518 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 7466 10656 7472 10668
rect 6825 10619 6883 10625
rect 7024 10628 7472 10656
rect 6362 10548 6368 10600
rect 6420 10588 6426 10600
rect 7024 10597 7052 10628
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 8018 10665 8024 10668
rect 8012 10656 8024 10665
rect 7979 10628 8024 10656
rect 8012 10619 8024 10628
rect 8018 10616 8024 10619
rect 8076 10616 8082 10668
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9306 10656 9312 10668
rect 9088 10628 9312 10656
rect 9088 10616 9094 10628
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10656 9919 10659
rect 10244 10656 10272 10755
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11609 10795 11667 10801
rect 11609 10792 11621 10795
rect 11388 10764 11621 10792
rect 11388 10752 11394 10764
rect 11609 10761 11621 10764
rect 11655 10792 11667 10795
rect 13906 10792 13912 10804
rect 11655 10764 13912 10792
rect 11655 10761 11667 10764
rect 11609 10755 11667 10761
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 12066 10684 12072 10736
rect 12124 10724 12130 10736
rect 12253 10727 12311 10733
rect 12253 10724 12265 10727
rect 12124 10696 12265 10724
rect 12124 10684 12130 10696
rect 12253 10693 12265 10696
rect 12299 10724 12311 10727
rect 15102 10724 15108 10736
rect 12299 10696 15108 10724
rect 12299 10693 12311 10696
rect 12253 10687 12311 10693
rect 15102 10684 15108 10696
rect 15160 10684 15166 10736
rect 9907 10628 10272 10656
rect 9907 10625 9919 10628
rect 9861 10619 9919 10625
rect 7009 10591 7067 10597
rect 7009 10588 7021 10591
rect 6420 10560 7021 10588
rect 6420 10548 6426 10560
rect 7009 10557 7021 10560
rect 7055 10557 7067 10591
rect 7193 10591 7251 10597
rect 7193 10588 7205 10591
rect 7009 10551 7067 10557
rect 7116 10560 7205 10588
rect 5629 10523 5687 10529
rect 5629 10520 5641 10523
rect 2746 10492 5641 10520
rect 2746 10464 2774 10492
rect 5629 10489 5641 10492
rect 5675 10489 5687 10523
rect 5629 10483 5687 10489
rect 5902 10480 5908 10532
rect 5960 10520 5966 10532
rect 7116 10520 7144 10560
rect 7193 10557 7205 10560
rect 7239 10588 7251 10591
rect 7374 10588 7380 10600
rect 7239 10560 7380 10588
rect 7239 10557 7251 10560
rect 7193 10551 7251 10557
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10557 7803 10591
rect 9508 10588 9536 10619
rect 10962 10616 10968 10668
rect 11020 10656 11026 10668
rect 11149 10659 11207 10665
rect 11149 10656 11161 10659
rect 11020 10628 11161 10656
rect 11020 10616 11026 10628
rect 11149 10625 11161 10628
rect 11195 10656 11207 10659
rect 13630 10656 13636 10668
rect 11195 10628 13636 10656
rect 11195 10625 11207 10628
rect 11149 10619 11207 10625
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9508 10560 10057 10588
rect 7745 10551 7803 10557
rect 10045 10557 10057 10560
rect 10091 10588 10103 10591
rect 11054 10588 11060 10600
rect 10091 10560 11060 10588
rect 10091 10557 10103 10560
rect 10045 10551 10103 10557
rect 7760 10520 7788 10551
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 11756 10560 11897 10588
rect 11756 10548 11762 10560
rect 11885 10557 11897 10560
rect 11931 10588 11943 10591
rect 14550 10588 14556 10600
rect 11931 10560 14556 10588
rect 11931 10557 11943 10560
rect 11885 10551 11943 10557
rect 14550 10548 14556 10560
rect 14608 10548 14614 10600
rect 5960 10492 7144 10520
rect 7208 10492 7788 10520
rect 5960 10480 5966 10492
rect 2682 10412 2688 10464
rect 2740 10424 2774 10464
rect 3559 10455 3617 10461
rect 2740 10412 2746 10424
rect 3559 10421 3571 10455
rect 3605 10452 3617 10455
rect 5258 10452 5264 10464
rect 3605 10424 5264 10452
rect 3605 10421 3617 10424
rect 3559 10415 3617 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 6380 10461 6408 10492
rect 7208 10464 7236 10492
rect 8754 10480 8760 10532
rect 8812 10520 8818 10532
rect 9309 10523 9367 10529
rect 9309 10520 9321 10523
rect 8812 10492 9321 10520
rect 8812 10480 8818 10492
rect 9309 10489 9321 10492
rect 9355 10489 9367 10523
rect 9309 10483 9367 10489
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 10413 10523 10471 10529
rect 10413 10520 10425 10523
rect 9824 10492 10425 10520
rect 9824 10480 9830 10492
rect 10413 10489 10425 10492
rect 10459 10520 10471 10523
rect 10686 10520 10692 10532
rect 10459 10492 10692 10520
rect 10459 10489 10471 10492
rect 10413 10483 10471 10489
rect 10686 10480 10692 10492
rect 10744 10480 10750 10532
rect 12526 10520 12532 10532
rect 12406 10492 12532 10520
rect 6365 10455 6423 10461
rect 6365 10421 6377 10455
rect 6411 10421 6423 10455
rect 6365 10415 6423 10421
rect 6454 10412 6460 10464
rect 6512 10452 6518 10464
rect 6641 10455 6699 10461
rect 6641 10452 6653 10455
rect 6512 10424 6653 10452
rect 6512 10412 6518 10424
rect 6641 10421 6653 10424
rect 6687 10421 6699 10455
rect 6641 10415 6699 10421
rect 7190 10412 7196 10464
rect 7248 10412 7254 10464
rect 7653 10455 7711 10461
rect 7653 10421 7665 10455
rect 7699 10452 7711 10455
rect 8846 10452 8852 10464
rect 7699 10424 8852 10452
rect 7699 10421 7711 10424
rect 7653 10415 7711 10421
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 9950 10452 9956 10464
rect 9723 10424 9956 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10042 10412 10048 10464
rect 10100 10452 10106 10464
rect 10597 10455 10655 10461
rect 10597 10452 10609 10455
rect 10100 10424 10609 10452
rect 10100 10412 10106 10424
rect 10597 10421 10609 10424
rect 10643 10452 10655 10455
rect 12406 10452 12434 10492
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 10643 10424 12434 10452
rect 10643 10421 10655 10424
rect 10597 10415 10655 10421
rect 1104 10362 16008 10384
rect 1104 10310 2824 10362
rect 2876 10310 2888 10362
rect 2940 10310 2952 10362
rect 3004 10310 3016 10362
rect 3068 10310 3080 10362
rect 3132 10310 6572 10362
rect 6624 10310 6636 10362
rect 6688 10310 6700 10362
rect 6752 10310 6764 10362
rect 6816 10310 6828 10362
rect 6880 10310 10320 10362
rect 10372 10310 10384 10362
rect 10436 10310 10448 10362
rect 10500 10310 10512 10362
rect 10564 10310 10576 10362
rect 10628 10310 14068 10362
rect 14120 10310 14132 10362
rect 14184 10310 14196 10362
rect 14248 10310 14260 10362
rect 14312 10310 14324 10362
rect 14376 10310 16008 10362
rect 1104 10288 16008 10310
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 8754 10248 8760 10260
rect 5868 10220 8760 10248
rect 5868 10208 5874 10220
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 9033 10251 9091 10257
rect 9033 10217 9045 10251
rect 9079 10248 9091 10251
rect 9306 10248 9312 10260
rect 9079 10220 9312 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 10042 10248 10048 10260
rect 9640 10220 10048 10248
rect 9640 10208 9646 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10778 10208 10784 10260
rect 10836 10248 10842 10260
rect 12253 10251 12311 10257
rect 12253 10248 12265 10251
rect 10836 10220 12265 10248
rect 10836 10208 10842 10220
rect 12253 10217 12265 10220
rect 12299 10217 12311 10251
rect 12989 10251 13047 10257
rect 12989 10248 13001 10251
rect 12253 10211 12311 10217
rect 12406 10220 13001 10248
rect 3510 10140 3516 10192
rect 3568 10180 3574 10192
rect 5077 10183 5135 10189
rect 5077 10180 5089 10183
rect 3568 10152 5089 10180
rect 3568 10140 3574 10152
rect 5077 10149 5089 10152
rect 5123 10149 5135 10183
rect 5077 10143 5135 10149
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 8573 10183 8631 10189
rect 8573 10180 8585 10183
rect 8444 10152 8585 10180
rect 8444 10140 8450 10152
rect 8573 10149 8585 10152
rect 8619 10149 8631 10183
rect 8573 10143 8631 10149
rect 9324 10152 10364 10180
rect 5350 10072 5356 10124
rect 5408 10112 5414 10124
rect 5721 10115 5779 10121
rect 5408 10084 5672 10112
rect 5408 10072 5414 10084
rect 4982 10044 4988 10056
rect 4943 10016 4988 10044
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5534 10044 5540 10056
rect 5491 10016 5540 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 5644 10044 5672 10084
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 5767 10084 7328 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 7190 10044 7196 10056
rect 5644 10016 5856 10044
rect 7151 10016 7196 10044
rect 5258 9936 5264 9988
rect 5316 9976 5322 9988
rect 5828 9976 5856 10016
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7300 10044 7328 10084
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 8665 10115 8723 10121
rect 8665 10112 8677 10115
rect 8352 10084 8677 10112
rect 8352 10072 8358 10084
rect 8665 10081 8677 10084
rect 8711 10081 8723 10115
rect 8665 10075 8723 10081
rect 8018 10044 8024 10056
rect 7300 10016 8024 10044
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 8754 10044 8760 10056
rect 8128 10016 8760 10044
rect 5997 9979 6055 9985
rect 5997 9976 6009 9979
rect 5316 9948 5764 9976
rect 5828 9948 6009 9976
rect 5316 9936 5322 9948
rect 3786 9868 3792 9920
rect 3844 9908 3850 9920
rect 4801 9911 4859 9917
rect 4801 9908 4813 9911
rect 3844 9880 4813 9908
rect 3844 9868 3850 9880
rect 4801 9877 4813 9880
rect 4847 9877 4859 9911
rect 4801 9871 4859 9877
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 5736 9908 5764 9948
rect 5997 9945 6009 9948
rect 6043 9945 6055 9979
rect 5997 9939 6055 9945
rect 6089 9979 6147 9985
rect 6089 9945 6101 9979
rect 6135 9945 6147 9979
rect 6089 9939 6147 9945
rect 6104 9908 6132 9939
rect 6362 9936 6368 9988
rect 6420 9976 6426 9988
rect 6822 9976 6828 9988
rect 6420 9948 6828 9976
rect 6420 9936 6426 9948
rect 6822 9936 6828 9948
rect 6880 9976 6886 9988
rect 7466 9985 7472 9988
rect 7009 9979 7067 9985
rect 7009 9976 7021 9979
rect 6880 9948 7021 9976
rect 6880 9936 6886 9948
rect 7009 9945 7021 9948
rect 7055 9945 7067 9979
rect 7460 9976 7472 9985
rect 7427 9948 7472 9976
rect 7009 9939 7067 9945
rect 7460 9939 7472 9948
rect 7524 9976 7530 9988
rect 8128 9976 8156 10016
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 8846 10004 8852 10056
rect 8904 10044 8910 10056
rect 9324 10044 9352 10152
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 10336 10121 10364 10152
rect 10870 10140 10876 10192
rect 10928 10180 10934 10192
rect 11517 10183 11575 10189
rect 11517 10180 11529 10183
rect 10928 10152 11529 10180
rect 10928 10140 10934 10152
rect 11517 10149 11529 10152
rect 11563 10149 11575 10183
rect 11517 10143 11575 10149
rect 9585 10115 9643 10121
rect 9585 10112 9597 10115
rect 9548 10084 9597 10112
rect 9548 10072 9554 10084
rect 9585 10081 9597 10084
rect 9631 10112 9643 10115
rect 10321 10115 10379 10121
rect 9631 10084 10088 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 8904 10016 9352 10044
rect 9401 10047 9459 10053
rect 8904 10004 8910 10016
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 7524 9948 8156 9976
rect 9416 9976 9444 10007
rect 10060 9976 10088 10084
rect 10321 10081 10333 10115
rect 10367 10081 10379 10115
rect 10321 10075 10379 10081
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10081 10471 10115
rect 12406 10112 12434 10220
rect 12989 10217 13001 10220
rect 13035 10217 13047 10251
rect 12989 10211 13047 10217
rect 13541 10251 13599 10257
rect 13541 10217 13553 10251
rect 13587 10248 13599 10251
rect 13814 10248 13820 10260
rect 13587 10220 13820 10248
rect 13587 10217 13599 10220
rect 13541 10211 13599 10217
rect 13556 10112 13584 10211
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 13725 10183 13783 10189
rect 13725 10149 13737 10183
rect 13771 10180 13783 10183
rect 14458 10180 14464 10192
rect 13771 10152 14464 10180
rect 13771 10149 13783 10152
rect 13725 10143 13783 10149
rect 10413 10075 10471 10081
rect 11072 10084 12434 10112
rect 12820 10084 13584 10112
rect 10226 10044 10232 10056
rect 10187 10016 10232 10044
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 10428 10044 10456 10075
rect 10962 10044 10968 10056
rect 10336 10016 10456 10044
rect 10923 10016 10968 10044
rect 10336 9976 10364 10016
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11072 9976 11100 10084
rect 11330 10044 11336 10056
rect 11291 10016 11336 10044
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 11698 10044 11704 10056
rect 11659 10016 11704 10044
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 12066 10044 12072 10056
rect 12027 10016 12072 10044
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 12820 10053 12848 10084
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10044 13231 10047
rect 13740 10044 13768 10143
rect 14458 10140 14464 10152
rect 14516 10140 14522 10192
rect 13219 10016 13768 10044
rect 13219 10013 13231 10016
rect 13173 10007 13231 10013
rect 9416 9948 9996 9976
rect 10060 9948 10364 9976
rect 10980 9948 11100 9976
rect 12452 9976 12480 10007
rect 12452 9948 13400 9976
rect 7466 9936 7472 9939
rect 7524 9936 7530 9948
rect 5592 9880 5637 9908
rect 5736 9880 6132 9908
rect 5592 9868 5598 9880
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 9493 9911 9551 9917
rect 9493 9908 9505 9911
rect 7984 9880 9505 9908
rect 7984 9868 7990 9880
rect 9493 9877 9505 9880
rect 9539 9908 9551 9911
rect 9582 9908 9588 9920
rect 9539 9880 9588 9908
rect 9539 9877 9551 9880
rect 9493 9871 9551 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 9858 9908 9864 9920
rect 9819 9880 9864 9908
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 9968 9908 9996 9948
rect 10980 9920 11008 9948
rect 13372 9920 13400 9948
rect 10594 9908 10600 9920
rect 9968 9880 10600 9908
rect 10594 9868 10600 9880
rect 10652 9868 10658 9920
rect 10778 9908 10784 9920
rect 10739 9880 10784 9908
rect 10778 9868 10784 9880
rect 10836 9868 10842 9920
rect 10962 9868 10968 9920
rect 11020 9868 11026 9920
rect 11146 9908 11152 9920
rect 11107 9880 11152 9908
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 11882 9908 11888 9920
rect 11843 9880 11888 9908
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 12621 9911 12679 9917
rect 12621 9908 12633 9911
rect 12584 9880 12633 9908
rect 12584 9868 12590 9880
rect 12621 9877 12633 9880
rect 12667 9877 12679 9911
rect 13354 9908 13360 9920
rect 13315 9880 13360 9908
rect 12621 9871 12679 9877
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 1104 9818 16008 9840
rect 1104 9766 4698 9818
rect 4750 9766 4762 9818
rect 4814 9766 4826 9818
rect 4878 9766 4890 9818
rect 4942 9766 4954 9818
rect 5006 9766 8446 9818
rect 8498 9766 8510 9818
rect 8562 9766 8574 9818
rect 8626 9766 8638 9818
rect 8690 9766 8702 9818
rect 8754 9766 12194 9818
rect 12246 9766 12258 9818
rect 12310 9766 12322 9818
rect 12374 9766 12386 9818
rect 12438 9766 12450 9818
rect 12502 9766 16008 9818
rect 1104 9744 16008 9766
rect 6641 9707 6699 9713
rect 6641 9704 6653 9707
rect 5276 9676 6653 9704
rect 1581 9639 1639 9645
rect 1581 9605 1593 9639
rect 1627 9636 1639 9639
rect 3234 9636 3240 9648
rect 1627 9608 3240 9636
rect 1627 9605 1639 9608
rect 1581 9599 1639 9605
rect 3234 9596 3240 9608
rect 3292 9596 3298 9648
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 5276 9636 5304 9676
rect 6641 9673 6653 9676
rect 6687 9673 6699 9707
rect 6641 9667 6699 9673
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 7248 9676 8340 9704
rect 7248 9664 7254 9676
rect 6914 9636 6920 9648
rect 4304 9608 5304 9636
rect 6196 9608 6920 9636
rect 4304 9596 4310 9608
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 5718 9568 5724 9580
rect 5491 9540 5724 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6196 9577 6224 9608
rect 6914 9596 6920 9608
rect 6972 9636 6978 9648
rect 7098 9636 7104 9648
rect 6972 9608 7104 9636
rect 6972 9596 6978 9608
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 7742 9596 7748 9648
rect 7800 9636 7806 9648
rect 8052 9639 8110 9645
rect 8052 9636 8064 9639
rect 7800 9608 8064 9636
rect 7800 9596 7806 9608
rect 8052 9605 8064 9608
rect 8098 9605 8110 9639
rect 8052 9599 8110 9605
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9537 5871 9571
rect 5813 9531 5871 9537
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 6457 9571 6515 9577
rect 6457 9537 6469 9571
rect 6503 9568 6515 9571
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6503 9540 6837 9568
rect 6503 9537 6515 9540
rect 6457 9531 6515 9537
rect 6825 9537 6837 9540
rect 6871 9568 6883 9571
rect 7466 9568 7472 9580
rect 6871 9540 7472 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 1486 9500 1492 9512
rect 1447 9472 1492 9500
rect 1486 9460 1492 9472
rect 1544 9460 1550 9512
rect 1762 9500 1768 9512
rect 1723 9472 1768 9500
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 5828 9500 5856 9531
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 8312 9512 8340 9676
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 8938 9704 8944 9716
rect 8444 9676 8944 9704
rect 8444 9664 8450 9676
rect 8938 9664 8944 9676
rect 8996 9704 9002 9716
rect 9490 9704 9496 9716
rect 8996 9676 9496 9704
rect 8996 9664 9002 9676
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 8404 9636 8432 9664
rect 8570 9636 8576 9648
rect 8404 9608 8576 9636
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 8662 9596 8668 9648
rect 8720 9636 8726 9648
rect 8849 9639 8907 9645
rect 8849 9636 8861 9639
rect 8720 9608 8861 9636
rect 8720 9596 8726 9608
rect 8849 9605 8861 9608
rect 8895 9636 8907 9639
rect 10226 9636 10232 9648
rect 8895 9608 10232 9636
rect 8895 9605 8907 9608
rect 8849 9599 8907 9605
rect 10226 9596 10232 9608
rect 10284 9596 10290 9648
rect 11241 9639 11299 9645
rect 11241 9636 11253 9639
rect 10336 9608 11253 9636
rect 8754 9568 8760 9580
rect 8715 9540 8760 9568
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 9490 9568 9496 9580
rect 9451 9540 9496 9568
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 9766 9568 9772 9580
rect 9600 9540 9772 9568
rect 8294 9509 8300 9512
rect 8290 9500 8300 9509
rect 5408 9472 5856 9500
rect 8255 9472 8300 9500
rect 5408 9460 5414 9472
rect 8290 9463 8300 9472
rect 8294 9460 8300 9463
rect 8352 9460 8358 9512
rect 8570 9460 8576 9512
rect 8628 9500 8634 9512
rect 9030 9500 9036 9512
rect 8628 9472 8708 9500
rect 8991 9472 9036 9500
rect 8628 9460 8634 9472
rect 3418 9392 3424 9444
rect 3476 9432 3482 9444
rect 5997 9435 6055 9441
rect 3476 9404 5764 9432
rect 3476 9392 3482 9404
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 5261 9367 5319 9373
rect 5261 9364 5273 9367
rect 1728 9336 5273 9364
rect 1728 9324 1734 9336
rect 5261 9333 5273 9336
rect 5307 9333 5319 9367
rect 5626 9364 5632 9376
rect 5587 9336 5632 9364
rect 5261 9327 5319 9333
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 5736 9364 5764 9404
rect 5997 9401 6009 9435
rect 6043 9401 6055 9435
rect 5997 9395 6055 9401
rect 6012 9364 6040 9395
rect 8386 9392 8392 9444
rect 8444 9432 8450 9444
rect 8680 9432 8708 9472
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9398 9460 9404 9512
rect 9456 9500 9462 9512
rect 9600 9500 9628 9540
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 10042 9568 10048 9580
rect 9907 9540 10048 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 10336 9577 10364 9608
rect 11241 9605 11253 9608
rect 11287 9636 11299 9639
rect 13538 9636 13544 9648
rect 11287 9608 13544 9636
rect 11287 9605 11299 9608
rect 11241 9599 11299 9605
rect 13538 9596 13544 9608
rect 13596 9596 13602 9648
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9537 10379 9571
rect 10321 9531 10379 9537
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9568 11115 9571
rect 11790 9568 11796 9580
rect 11103 9540 11796 9568
rect 11103 9537 11115 9540
rect 11057 9531 11115 9537
rect 9456 9472 9628 9500
rect 9456 9460 9462 9472
rect 9674 9460 9680 9512
rect 9732 9460 9738 9512
rect 10704 9500 10732 9531
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9568 12311 9571
rect 12621 9571 12679 9577
rect 12299 9540 12434 9568
rect 12299 9537 12311 9540
rect 12253 9531 12311 9537
rect 12406 9500 12434 9540
rect 12621 9537 12633 9571
rect 12667 9568 12679 9571
rect 12986 9568 12992 9580
rect 12667 9540 12992 9568
rect 12667 9537 12679 9540
rect 12621 9531 12679 9537
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 10704 9472 11652 9500
rect 12406 9472 12848 9500
rect 9309 9435 9367 9441
rect 9309 9432 9321 9435
rect 8444 9404 8489 9432
rect 8680 9404 9321 9432
rect 8444 9392 8450 9404
rect 9309 9401 9321 9404
rect 9355 9401 9367 9435
rect 9692 9432 9720 9460
rect 10873 9435 10931 9441
rect 10873 9432 10885 9435
rect 9692 9404 10885 9432
rect 9309 9395 9367 9401
rect 10873 9401 10885 9404
rect 10919 9401 10931 9435
rect 10873 9395 10931 9401
rect 11624 9376 11652 9472
rect 11974 9392 11980 9444
rect 12032 9432 12038 9444
rect 12069 9435 12127 9441
rect 12069 9432 12081 9435
rect 12032 9404 12081 9432
rect 12032 9392 12038 9404
rect 12069 9401 12081 9404
rect 12115 9401 12127 9435
rect 12069 9395 12127 9401
rect 12437 9435 12495 9441
rect 12437 9401 12449 9435
rect 12483 9432 12495 9435
rect 12618 9432 12624 9444
rect 12483 9404 12624 9432
rect 12483 9401 12495 9404
rect 12437 9395 12495 9401
rect 12618 9392 12624 9404
rect 12676 9392 12682 9444
rect 12820 9441 12848 9472
rect 12805 9435 12863 9441
rect 12805 9401 12817 9435
rect 12851 9432 12863 9435
rect 15102 9432 15108 9444
rect 12851 9404 15108 9432
rect 12851 9401 12863 9404
rect 12805 9395 12863 9401
rect 15102 9392 15108 9404
rect 15160 9392 15166 9444
rect 5736 9336 6040 9364
rect 6917 9367 6975 9373
rect 6917 9333 6929 9367
rect 6963 9364 6975 9367
rect 7098 9364 7104 9376
rect 6963 9336 7104 9364
rect 6963 9333 6975 9336
rect 6917 9327 6975 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 9122 9324 9128 9376
rect 9180 9364 9186 9376
rect 9582 9364 9588 9376
rect 9180 9336 9588 9364
rect 9180 9324 9186 9336
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 9766 9364 9772 9376
rect 9723 9336 9772 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 10137 9367 10195 9373
rect 10137 9333 10149 9367
rect 10183 9364 10195 9367
rect 10318 9364 10324 9376
rect 10183 9336 10324 9364
rect 10183 9333 10195 9336
rect 10137 9327 10195 9333
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10502 9364 10508 9376
rect 10463 9336 10508 9364
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 11606 9364 11612 9376
rect 11567 9336 11612 9364
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 11790 9364 11796 9376
rect 11751 9336 11796 9364
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 12986 9364 12992 9376
rect 12947 9336 12992 9364
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 1104 9274 16008 9296
rect 1104 9222 2824 9274
rect 2876 9222 2888 9274
rect 2940 9222 2952 9274
rect 3004 9222 3016 9274
rect 3068 9222 3080 9274
rect 3132 9222 6572 9274
rect 6624 9222 6636 9274
rect 6688 9222 6700 9274
rect 6752 9222 6764 9274
rect 6816 9222 6828 9274
rect 6880 9222 10320 9274
rect 10372 9222 10384 9274
rect 10436 9222 10448 9274
rect 10500 9222 10512 9274
rect 10564 9222 10576 9274
rect 10628 9222 14068 9274
rect 14120 9222 14132 9274
rect 14184 9222 14196 9274
rect 14248 9222 14260 9274
rect 14312 9222 14324 9274
rect 14376 9222 16008 9274
rect 1104 9200 16008 9222
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 5994 9160 6000 9172
rect 5408 9132 6000 9160
rect 5408 9120 5414 9132
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 7190 9160 7196 9172
rect 6840 9132 7196 9160
rect 4338 9052 4344 9104
rect 4396 9092 4402 9104
rect 6840 9092 6868 9132
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 8018 9120 8024 9172
rect 8076 9160 8082 9172
rect 8205 9163 8263 9169
rect 8205 9160 8217 9163
rect 8076 9132 8217 9160
rect 8076 9120 8082 9132
rect 8205 9129 8217 9132
rect 8251 9129 8263 9163
rect 8205 9123 8263 9129
rect 8754 9120 8760 9172
rect 8812 9160 8818 9172
rect 9122 9160 9128 9172
rect 8812 9132 9128 9160
rect 8812 9120 8818 9132
rect 9122 9120 9128 9132
rect 9180 9160 9186 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 9180 9132 9413 9160
rect 9180 9120 9186 9132
rect 9401 9129 9413 9132
rect 9447 9129 9459 9163
rect 10134 9160 10140 9172
rect 10095 9132 10140 9160
rect 9401 9123 9459 9129
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 4396 9064 6868 9092
rect 4396 9052 4402 9064
rect 6840 9033 6868 9064
rect 7834 9052 7840 9104
rect 7892 9092 7898 9104
rect 11882 9092 11888 9104
rect 7892 9064 11888 9092
rect 7892 9052 7898 9064
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 9024 6883 9027
rect 9306 9024 9312 9036
rect 6871 8996 6905 9024
rect 7852 8996 9312 9024
rect 6871 8993 6883 8996
rect 6825 8987 6883 8993
rect 6365 8959 6423 8965
rect 6365 8925 6377 8959
rect 6411 8956 6423 8959
rect 6914 8956 6920 8968
rect 6411 8928 6920 8956
rect 6411 8925 6423 8928
rect 6365 8919 6423 8925
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 7098 8965 7104 8968
rect 7092 8956 7104 8965
rect 7059 8928 7104 8956
rect 7092 8919 7104 8928
rect 7098 8916 7104 8919
rect 7156 8916 7162 8968
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 7852 8956 7880 8996
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 9548 8996 9689 9024
rect 9548 8984 9554 8996
rect 9677 8993 9689 8996
rect 9723 9024 9735 9027
rect 12802 9024 12808 9036
rect 9723 8996 12808 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 7524 8928 7880 8956
rect 7524 8916 7530 8928
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 8386 8956 8392 8968
rect 8260 8928 8392 8956
rect 8260 8916 8266 8928
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 8665 8959 8723 8965
rect 8665 8925 8677 8959
rect 8711 8925 8723 8959
rect 8665 8919 8723 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 10134 8956 10140 8968
rect 9263 8928 10140 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 4614 8848 4620 8900
rect 4672 8888 4678 8900
rect 4672 8860 5856 8888
rect 4672 8848 4678 8860
rect 1486 8820 1492 8832
rect 1399 8792 1492 8820
rect 1486 8780 1492 8792
rect 1544 8820 1550 8832
rect 3142 8820 3148 8832
rect 1544 8792 3148 8820
rect 1544 8780 1550 8792
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 5629 8823 5687 8829
rect 5629 8789 5641 8823
rect 5675 8820 5687 8823
rect 5718 8820 5724 8832
rect 5675 8792 5724 8820
rect 5675 8789 5687 8792
rect 5629 8783 5687 8789
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 5828 8820 5856 8860
rect 5902 8848 5908 8900
rect 5960 8888 5966 8900
rect 8570 8888 8576 8900
rect 5960 8860 8576 8888
rect 5960 8848 5966 8860
rect 8570 8848 8576 8860
rect 8628 8848 8634 8900
rect 8680 8888 8708 8919
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 9674 8888 9680 8900
rect 8680 8860 9680 8888
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 9861 8891 9919 8897
rect 9861 8857 9873 8891
rect 9907 8888 9919 8891
rect 10226 8888 10232 8900
rect 9907 8860 10232 8888
rect 9907 8857 9919 8860
rect 9861 8851 9919 8857
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 8481 8823 8539 8829
rect 8481 8820 8493 8823
rect 5828 8792 8493 8820
rect 8481 8789 8493 8792
rect 8527 8789 8539 8823
rect 9030 8820 9036 8832
rect 8991 8792 9036 8820
rect 8481 8783 8539 8789
rect 9030 8780 9036 8792
rect 9088 8780 9094 8832
rect 10042 8820 10048 8832
rect 10003 8792 10048 8820
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 1104 8730 16008 8752
rect 1104 8678 4698 8730
rect 4750 8678 4762 8730
rect 4814 8678 4826 8730
rect 4878 8678 4890 8730
rect 4942 8678 4954 8730
rect 5006 8678 8446 8730
rect 8498 8678 8510 8730
rect 8562 8678 8574 8730
rect 8626 8678 8638 8730
rect 8690 8678 8702 8730
rect 8754 8678 12194 8730
rect 12246 8678 12258 8730
rect 12310 8678 12322 8730
rect 12374 8678 12386 8730
rect 12438 8678 12450 8730
rect 12502 8678 16008 8730
rect 1104 8656 16008 8678
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 7101 8619 7159 8625
rect 7101 8616 7113 8619
rect 5592 8588 7113 8616
rect 5592 8576 5598 8588
rect 7101 8585 7113 8588
rect 7147 8585 7159 8619
rect 7101 8579 7159 8585
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7515 8588 8033 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 8202 8576 8208 8628
rect 8260 8616 8266 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 8260 8588 8493 8616
rect 8260 8576 8266 8588
rect 8481 8585 8493 8588
rect 8527 8585 8539 8619
rect 8481 8579 8539 8585
rect 8941 8619 8999 8625
rect 8941 8585 8953 8619
rect 8987 8616 8999 8619
rect 9674 8616 9680 8628
rect 8987 8588 9680 8616
rect 8987 8585 8999 8588
rect 8941 8579 8999 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 11701 8551 11759 8557
rect 11701 8548 11713 8551
rect 8352 8520 11713 8548
rect 8352 8508 8358 8520
rect 11701 8517 11713 8520
rect 11747 8517 11759 8551
rect 11701 8511 11759 8517
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8480 7619 8483
rect 7607 8452 8340 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 7098 8372 7104 8424
rect 7156 8412 7162 8424
rect 7650 8412 7656 8424
rect 7156 8384 7656 8412
rect 7156 8372 7162 8384
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 8312 8412 8340 8452
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 9858 8480 9864 8492
rect 8444 8452 8489 8480
rect 8588 8452 9864 8480
rect 8444 8440 8450 8452
rect 8588 8412 8616 8452
rect 9858 8440 9864 8452
rect 9916 8440 9922 8492
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 12575 8452 12756 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 8312 8384 8616 8412
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8412 8723 8415
rect 8846 8412 8852 8424
rect 8711 8384 8852 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 8846 8372 8852 8384
rect 8904 8372 8910 8424
rect 12728 8356 12756 8452
rect 12710 8344 12716 8356
rect 12671 8316 12716 8344
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 8386 8236 8392 8288
rect 8444 8276 8450 8288
rect 9125 8279 9183 8285
rect 9125 8276 9137 8279
rect 8444 8248 9137 8276
rect 8444 8236 8450 8248
rect 9125 8245 9137 8248
rect 9171 8276 9183 8279
rect 9490 8276 9496 8288
rect 9171 8248 9496 8276
rect 9171 8245 9183 8248
rect 9125 8239 9183 8245
rect 9490 8236 9496 8248
rect 9548 8236 9554 8288
rect 1104 8186 16008 8208
rect 1104 8134 2824 8186
rect 2876 8134 2888 8186
rect 2940 8134 2952 8186
rect 3004 8134 3016 8186
rect 3068 8134 3080 8186
rect 3132 8134 6572 8186
rect 6624 8134 6636 8186
rect 6688 8134 6700 8186
rect 6752 8134 6764 8186
rect 6816 8134 6828 8186
rect 6880 8134 10320 8186
rect 10372 8134 10384 8186
rect 10436 8134 10448 8186
rect 10500 8134 10512 8186
rect 10564 8134 10576 8186
rect 10628 8134 14068 8186
rect 14120 8134 14132 8186
rect 14184 8134 14196 8186
rect 14248 8134 14260 8186
rect 14312 8134 14324 8186
rect 14376 8134 16008 8186
rect 1104 8112 16008 8134
rect 5074 7896 5080 7948
rect 5132 7936 5138 7948
rect 7282 7936 7288 7948
rect 5132 7908 7288 7936
rect 5132 7896 5138 7908
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 1104 7642 16008 7664
rect 1104 7590 4698 7642
rect 4750 7590 4762 7642
rect 4814 7590 4826 7642
rect 4878 7590 4890 7642
rect 4942 7590 4954 7642
rect 5006 7590 8446 7642
rect 8498 7590 8510 7642
rect 8562 7590 8574 7642
rect 8626 7590 8638 7642
rect 8690 7590 8702 7642
rect 8754 7590 12194 7642
rect 12246 7590 12258 7642
rect 12310 7590 12322 7642
rect 12374 7590 12386 7642
rect 12438 7590 12450 7642
rect 12502 7590 16008 7642
rect 1104 7568 16008 7590
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 3384 7500 5733 7528
rect 3384 7488 3390 7500
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 7742 7528 7748 7540
rect 5721 7491 5779 7497
rect 5920 7500 7748 7528
rect 4985 7463 5043 7469
rect 4985 7460 4997 7463
rect 4816 7432 4997 7460
rect 3510 7392 3516 7404
rect 3471 7364 3516 7392
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 4816 7401 4844 7432
rect 4985 7429 4997 7432
rect 5031 7460 5043 7463
rect 5074 7460 5080 7472
rect 5031 7432 5080 7460
rect 5031 7429 5043 7432
rect 4985 7423 5043 7429
rect 5074 7420 5080 7432
rect 5132 7420 5138 7472
rect 5445 7463 5503 7469
rect 5445 7460 5457 7463
rect 5368 7432 5457 7460
rect 5368 7401 5396 7432
rect 5445 7429 5457 7432
rect 5491 7460 5503 7463
rect 5920 7460 5948 7500
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 7837 7531 7895 7537
rect 7837 7497 7849 7531
rect 7883 7528 7895 7531
rect 7926 7528 7932 7540
rect 7883 7500 7932 7528
rect 7883 7497 7895 7500
rect 7837 7491 7895 7497
rect 5491 7432 5948 7460
rect 5491 7429 5503 7432
rect 5445 7423 5503 7429
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7392 7711 7395
rect 7852 7392 7880 7491
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 9398 7488 9404 7540
rect 9456 7528 9462 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 9456 7500 9597 7528
rect 9456 7488 9462 7500
rect 9508 7401 9536 7500
rect 9585 7497 9597 7500
rect 9631 7497 9643 7531
rect 9585 7491 9643 7497
rect 7699 7364 7880 7392
rect 9493 7395 9551 7401
rect 7699 7361 7711 7364
rect 7653 7355 7711 7361
rect 9493 7361 9505 7395
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 3234 7324 3240 7336
rect 3195 7296 3240 7324
rect 3234 7284 3240 7296
rect 3292 7284 3298 7336
rect 5920 7324 5948 7355
rect 6089 7327 6147 7333
rect 6089 7324 6101 7327
rect 5920 7296 6101 7324
rect 6089 7293 6101 7296
rect 6135 7324 6147 7327
rect 9122 7324 9128 7336
rect 6135 7296 9128 7324
rect 6135 7293 6147 7296
rect 6089 7287 6147 7293
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 5074 7216 5080 7268
rect 5132 7256 5138 7268
rect 5132 7228 6132 7256
rect 5132 7216 5138 7228
rect 4614 7188 4620 7200
rect 4575 7160 4620 7188
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 5166 7188 5172 7200
rect 5127 7160 5172 7188
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 6104 7188 6132 7228
rect 7282 7216 7288 7268
rect 7340 7256 7346 7268
rect 9309 7259 9367 7265
rect 9309 7256 9321 7259
rect 7340 7228 9321 7256
rect 7340 7216 7346 7228
rect 9309 7225 9321 7228
rect 9355 7225 9367 7259
rect 9309 7219 9367 7225
rect 7469 7191 7527 7197
rect 7469 7188 7481 7191
rect 6104 7160 7481 7188
rect 7469 7157 7481 7160
rect 7515 7157 7527 7191
rect 7469 7151 7527 7157
rect 1104 7098 16008 7120
rect 1104 7046 2824 7098
rect 2876 7046 2888 7098
rect 2940 7046 2952 7098
rect 3004 7046 3016 7098
rect 3068 7046 3080 7098
rect 3132 7046 6572 7098
rect 6624 7046 6636 7098
rect 6688 7046 6700 7098
rect 6752 7046 6764 7098
rect 6816 7046 6828 7098
rect 6880 7046 10320 7098
rect 10372 7046 10384 7098
rect 10436 7046 10448 7098
rect 10500 7046 10512 7098
rect 10564 7046 10576 7098
rect 10628 7046 14068 7098
rect 14120 7046 14132 7098
rect 14184 7046 14196 7098
rect 14248 7046 14260 7098
rect 14312 7046 14324 7098
rect 14376 7046 16008 7098
rect 1104 7024 16008 7046
rect 1104 6554 16008 6576
rect 1104 6502 4698 6554
rect 4750 6502 4762 6554
rect 4814 6502 4826 6554
rect 4878 6502 4890 6554
rect 4942 6502 4954 6554
rect 5006 6502 8446 6554
rect 8498 6502 8510 6554
rect 8562 6502 8574 6554
rect 8626 6502 8638 6554
rect 8690 6502 8702 6554
rect 8754 6502 12194 6554
rect 12246 6502 12258 6554
rect 12310 6502 12322 6554
rect 12374 6502 12386 6554
rect 12438 6502 12450 6554
rect 12502 6502 16008 6554
rect 1104 6480 16008 6502
rect 1104 6010 16008 6032
rect 1104 5958 2824 6010
rect 2876 5958 2888 6010
rect 2940 5958 2952 6010
rect 3004 5958 3016 6010
rect 3068 5958 3080 6010
rect 3132 5958 6572 6010
rect 6624 5958 6636 6010
rect 6688 5958 6700 6010
rect 6752 5958 6764 6010
rect 6816 5958 6828 6010
rect 6880 5958 10320 6010
rect 10372 5958 10384 6010
rect 10436 5958 10448 6010
rect 10500 5958 10512 6010
rect 10564 5958 10576 6010
rect 10628 5958 14068 6010
rect 14120 5958 14132 6010
rect 14184 5958 14196 6010
rect 14248 5958 14260 6010
rect 14312 5958 14324 6010
rect 14376 5958 16008 6010
rect 1104 5936 16008 5958
rect 1104 5466 16008 5488
rect 1104 5414 4698 5466
rect 4750 5414 4762 5466
rect 4814 5414 4826 5466
rect 4878 5414 4890 5466
rect 4942 5414 4954 5466
rect 5006 5414 8446 5466
rect 8498 5414 8510 5466
rect 8562 5414 8574 5466
rect 8626 5414 8638 5466
rect 8690 5414 8702 5466
rect 8754 5414 12194 5466
rect 12246 5414 12258 5466
rect 12310 5414 12322 5466
rect 12374 5414 12386 5466
rect 12438 5414 12450 5466
rect 12502 5414 16008 5466
rect 1104 5392 16008 5414
rect 1104 4922 16008 4944
rect 1104 4870 2824 4922
rect 2876 4870 2888 4922
rect 2940 4870 2952 4922
rect 3004 4870 3016 4922
rect 3068 4870 3080 4922
rect 3132 4870 6572 4922
rect 6624 4870 6636 4922
rect 6688 4870 6700 4922
rect 6752 4870 6764 4922
rect 6816 4870 6828 4922
rect 6880 4870 10320 4922
rect 10372 4870 10384 4922
rect 10436 4870 10448 4922
rect 10500 4870 10512 4922
rect 10564 4870 10576 4922
rect 10628 4870 14068 4922
rect 14120 4870 14132 4922
rect 14184 4870 14196 4922
rect 14248 4870 14260 4922
rect 14312 4870 14324 4922
rect 14376 4870 16008 4922
rect 1104 4848 16008 4870
rect 1104 4378 16008 4400
rect 1104 4326 4698 4378
rect 4750 4326 4762 4378
rect 4814 4326 4826 4378
rect 4878 4326 4890 4378
rect 4942 4326 4954 4378
rect 5006 4326 8446 4378
rect 8498 4326 8510 4378
rect 8562 4326 8574 4378
rect 8626 4326 8638 4378
rect 8690 4326 8702 4378
rect 8754 4326 12194 4378
rect 12246 4326 12258 4378
rect 12310 4326 12322 4378
rect 12374 4326 12386 4378
rect 12438 4326 12450 4378
rect 12502 4326 16008 4378
rect 1104 4304 16008 4326
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 6454 4128 6460 4140
rect 4028 4100 6460 4128
rect 4028 4088 4034 4100
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 8846 4128 8852 4140
rect 7432 4100 8852 4128
rect 7432 4088 7438 4100
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 9674 4088 9680 4140
rect 9732 4128 9738 4140
rect 12066 4128 12072 4140
rect 9732 4100 12072 4128
rect 9732 4088 9738 4100
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 15746 4128 15752 4140
rect 13044 4100 15752 4128
rect 13044 4088 13050 4100
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 5718 4020 5724 4072
rect 5776 4060 5782 4072
rect 9122 4060 9128 4072
rect 5776 4032 9128 4060
rect 5776 4020 5782 4032
rect 9122 4020 9128 4032
rect 9180 4020 9186 4072
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 11698 4060 11704 4072
rect 9364 4032 11704 4060
rect 9364 4020 9370 4032
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 13354 4020 13360 4072
rect 13412 4060 13418 4072
rect 15010 4060 15016 4072
rect 13412 4032 15016 4060
rect 13412 4020 13418 4032
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 3602 3952 3608 4004
rect 3660 3992 3666 4004
rect 7006 3992 7012 4004
rect 3660 3964 7012 3992
rect 3660 3952 3666 3964
rect 7006 3952 7012 3964
rect 7064 3952 7070 4004
rect 8294 3952 8300 4004
rect 8352 3992 8358 4004
rect 10962 3992 10968 4004
rect 8352 3964 10968 3992
rect 8352 3952 8358 3964
rect 10962 3952 10968 3964
rect 11020 3952 11026 4004
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 8110 3924 8116 3936
rect 4396 3896 8116 3924
rect 4396 3884 4402 3896
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 1104 3834 16008 3856
rect 1104 3782 2824 3834
rect 2876 3782 2888 3834
rect 2940 3782 2952 3834
rect 3004 3782 3016 3834
rect 3068 3782 3080 3834
rect 3132 3782 6572 3834
rect 6624 3782 6636 3834
rect 6688 3782 6700 3834
rect 6752 3782 6764 3834
rect 6816 3782 6828 3834
rect 6880 3782 10320 3834
rect 10372 3782 10384 3834
rect 10436 3782 10448 3834
rect 10500 3782 10512 3834
rect 10564 3782 10576 3834
rect 10628 3782 14068 3834
rect 14120 3782 14132 3834
rect 14184 3782 14196 3834
rect 14248 3782 14260 3834
rect 14312 3782 14324 3834
rect 14376 3782 16008 3834
rect 1104 3760 16008 3782
rect 1394 3680 1400 3732
rect 1452 3720 1458 3732
rect 4614 3720 4620 3732
rect 1452 3692 4620 3720
rect 1452 3680 1458 3692
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 6086 3680 6092 3732
rect 6144 3720 6150 3732
rect 9858 3720 9864 3732
rect 6144 3692 9864 3720
rect 6144 3680 6150 3692
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 11790 3680 11796 3732
rect 11848 3720 11854 3732
rect 13906 3720 13912 3732
rect 11848 3692 13912 3720
rect 11848 3680 11854 3692
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 10686 3612 10692 3664
rect 10744 3652 10750 3664
rect 14642 3652 14648 3664
rect 10744 3624 14648 3652
rect 10744 3612 10750 3624
rect 14642 3612 14648 3624
rect 14700 3612 14706 3664
rect 4614 3544 4620 3596
rect 4672 3584 4678 3596
rect 9030 3584 9036 3596
rect 4672 3556 9036 3584
rect 4672 3544 4678 3556
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 12526 3584 12532 3596
rect 9548 3556 12532 3584
rect 9548 3544 9554 3556
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 2130 3476 2136 3528
rect 2188 3516 2194 3528
rect 5166 3516 5172 3528
rect 2188 3488 5172 3516
rect 2188 3476 2194 3488
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 7558 3476 7564 3528
rect 7616 3516 7622 3528
rect 10962 3516 10968 3528
rect 7616 3488 10968 3516
rect 7616 3476 7622 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 1762 3408 1768 3460
rect 1820 3448 1826 3460
rect 3786 3448 3792 3460
rect 1820 3420 3792 3448
rect 1820 3408 1826 3420
rect 3786 3408 3792 3420
rect 3844 3408 3850 3460
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 10870 3448 10876 3460
rect 6972 3420 10876 3448
rect 6972 3408 6978 3420
rect 10870 3408 10876 3420
rect 10928 3408 10934 3460
rect 11606 3408 11612 3460
rect 11664 3448 11670 3460
rect 13814 3448 13820 3460
rect 11664 3420 13820 3448
rect 11664 3408 11670 3420
rect 13814 3408 13820 3420
rect 13872 3408 13878 3460
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 13170 3380 13176 3392
rect 10100 3352 13176 3380
rect 10100 3340 10106 3352
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 1104 3290 16008 3312
rect 1104 3238 4698 3290
rect 4750 3238 4762 3290
rect 4814 3238 4826 3290
rect 4878 3238 4890 3290
rect 4942 3238 4954 3290
rect 5006 3238 8446 3290
rect 8498 3238 8510 3290
rect 8562 3238 8574 3290
rect 8626 3238 8638 3290
rect 8690 3238 8702 3290
rect 8754 3238 12194 3290
rect 12246 3238 12258 3290
rect 12310 3238 12322 3290
rect 12374 3238 12386 3290
rect 12438 3238 12450 3290
rect 12502 3238 16008 3290
rect 1104 3216 16008 3238
rect 6270 3136 6276 3188
rect 6328 3176 6334 3188
rect 10686 3176 10692 3188
rect 6328 3148 10692 3176
rect 6328 3136 6334 3148
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 2498 3068 2504 3120
rect 2556 3108 2562 3120
rect 5626 3108 5632 3120
rect 2556 3080 5632 3108
rect 2556 3068 2562 3080
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 6178 3068 6184 3120
rect 6236 3108 6242 3120
rect 10778 3108 10784 3120
rect 6236 3080 10784 3108
rect 6236 3068 6242 3080
rect 10778 3068 10784 3080
rect 10836 3068 10842 3120
rect 5810 2796 5816 2848
rect 5868 2836 5874 2848
rect 9950 2836 9956 2848
rect 5868 2808 9956 2836
rect 5868 2796 5874 2808
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 1104 2746 16008 2768
rect 1104 2694 2824 2746
rect 2876 2694 2888 2746
rect 2940 2694 2952 2746
rect 3004 2694 3016 2746
rect 3068 2694 3080 2746
rect 3132 2694 6572 2746
rect 6624 2694 6636 2746
rect 6688 2694 6700 2746
rect 6752 2694 6764 2746
rect 6816 2694 6828 2746
rect 6880 2694 10320 2746
rect 10372 2694 10384 2746
rect 10436 2694 10448 2746
rect 10500 2694 10512 2746
rect 10564 2694 10576 2746
rect 10628 2694 14068 2746
rect 14120 2694 14132 2746
rect 14184 2694 14196 2746
rect 14248 2694 14260 2746
rect 14312 2694 14324 2746
rect 14376 2694 16008 2746
rect 1104 2672 16008 2694
rect 2866 2592 2872 2644
rect 2924 2632 2930 2644
rect 3326 2632 3332 2644
rect 2924 2604 3332 2632
rect 2924 2592 2930 2604
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 6362 2592 6368 2644
rect 6420 2632 6426 2644
rect 12434 2632 12440 2644
rect 6420 2604 12440 2632
rect 6420 2592 6426 2604
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 1104 2202 16008 2224
rect 1104 2150 4698 2202
rect 4750 2150 4762 2202
rect 4814 2150 4826 2202
rect 4878 2150 4890 2202
rect 4942 2150 4954 2202
rect 5006 2150 8446 2202
rect 8498 2150 8510 2202
rect 8562 2150 8574 2202
rect 8626 2150 8638 2202
rect 8690 2150 8702 2202
rect 8754 2150 12194 2202
rect 12246 2150 12258 2202
rect 12310 2150 12322 2202
rect 12374 2150 12386 2202
rect 12438 2150 12450 2202
rect 12502 2150 16008 2202
rect 1104 2128 16008 2150
<< via1 >>
rect 4160 17892 4212 17944
rect 4344 17892 4396 17944
rect 4698 17382 4750 17434
rect 4762 17382 4814 17434
rect 4826 17382 4878 17434
rect 4890 17382 4942 17434
rect 4954 17382 5006 17434
rect 8446 17382 8498 17434
rect 8510 17382 8562 17434
rect 8574 17382 8626 17434
rect 8638 17382 8690 17434
rect 8702 17382 8754 17434
rect 12194 17382 12246 17434
rect 12258 17382 12310 17434
rect 12322 17382 12374 17434
rect 12386 17382 12438 17434
rect 12450 17382 12502 17434
rect 2824 16838 2876 16890
rect 2888 16838 2940 16890
rect 2952 16838 3004 16890
rect 3016 16838 3068 16890
rect 3080 16838 3132 16890
rect 6572 16838 6624 16890
rect 6636 16838 6688 16890
rect 6700 16838 6752 16890
rect 6764 16838 6816 16890
rect 6828 16838 6880 16890
rect 10320 16838 10372 16890
rect 10384 16838 10436 16890
rect 10448 16838 10500 16890
rect 10512 16838 10564 16890
rect 10576 16838 10628 16890
rect 14068 16838 14120 16890
rect 14132 16838 14184 16890
rect 14196 16838 14248 16890
rect 14260 16838 14312 16890
rect 14324 16838 14376 16890
rect 5724 16532 5776 16584
rect 6092 16532 6144 16584
rect 4698 16294 4750 16346
rect 4762 16294 4814 16346
rect 4826 16294 4878 16346
rect 4890 16294 4942 16346
rect 4954 16294 5006 16346
rect 8446 16294 8498 16346
rect 8510 16294 8562 16346
rect 8574 16294 8626 16346
rect 8638 16294 8690 16346
rect 8702 16294 8754 16346
rect 12194 16294 12246 16346
rect 12258 16294 12310 16346
rect 12322 16294 12374 16346
rect 12386 16294 12438 16346
rect 12450 16294 12502 16346
rect 5724 16056 5776 16108
rect 6460 16056 6512 16108
rect 3792 15988 3844 16040
rect 5356 15988 5408 16040
rect 6460 15920 6512 15972
rect 11520 15920 11572 15972
rect 7196 15852 7248 15904
rect 10784 15852 10836 15904
rect 2824 15750 2876 15802
rect 2888 15750 2940 15802
rect 2952 15750 3004 15802
rect 3016 15750 3068 15802
rect 3080 15750 3132 15802
rect 6572 15750 6624 15802
rect 6636 15750 6688 15802
rect 6700 15750 6752 15802
rect 6764 15750 6816 15802
rect 6828 15750 6880 15802
rect 10320 15750 10372 15802
rect 10384 15750 10436 15802
rect 10448 15750 10500 15802
rect 10512 15750 10564 15802
rect 10576 15750 10628 15802
rect 14068 15750 14120 15802
rect 14132 15750 14184 15802
rect 14196 15750 14248 15802
rect 14260 15750 14312 15802
rect 14324 15750 14376 15802
rect 7104 15648 7156 15700
rect 9680 15648 9732 15700
rect 11152 15648 11204 15700
rect 14832 15648 14884 15700
rect 4344 15580 4396 15632
rect 7656 15580 7708 15632
rect 8208 15580 8260 15632
rect 11980 15580 12032 15632
rect 3424 15512 3476 15564
rect 5816 15512 5868 15564
rect 8852 15512 8904 15564
rect 12624 15512 12676 15564
rect 2320 15444 2372 15496
rect 3976 15444 4028 15496
rect 7472 15444 7524 15496
rect 9404 15444 9456 15496
rect 10140 15444 10192 15496
rect 12072 15444 12124 15496
rect 3148 15376 3200 15428
rect 5908 15376 5960 15428
rect 7840 15376 7892 15428
rect 10784 15376 10836 15428
rect 11060 15376 11112 15428
rect 12992 15376 13044 15428
rect 13820 15376 13872 15428
rect 15568 15376 15620 15428
rect 1584 15308 1636 15360
rect 4068 15308 4120 15360
rect 5264 15308 5316 15360
rect 7472 15308 7524 15360
rect 9036 15308 9088 15360
rect 10232 15308 10284 15360
rect 10692 15308 10744 15360
rect 13360 15308 13412 15360
rect 14464 15308 14516 15360
rect 15936 15308 15988 15360
rect 4698 15206 4750 15258
rect 4762 15206 4814 15258
rect 4826 15206 4878 15258
rect 4890 15206 4942 15258
rect 4954 15206 5006 15258
rect 8446 15206 8498 15258
rect 8510 15206 8562 15258
rect 8574 15206 8626 15258
rect 8638 15206 8690 15258
rect 8702 15206 8754 15258
rect 12194 15206 12246 15258
rect 12258 15206 12310 15258
rect 12322 15206 12374 15258
rect 12386 15206 12438 15258
rect 12450 15206 12502 15258
rect 2824 14662 2876 14714
rect 2888 14662 2940 14714
rect 2952 14662 3004 14714
rect 3016 14662 3068 14714
rect 3080 14662 3132 14714
rect 6572 14662 6624 14714
rect 6636 14662 6688 14714
rect 6700 14662 6752 14714
rect 6764 14662 6816 14714
rect 6828 14662 6880 14714
rect 10320 14662 10372 14714
rect 10384 14662 10436 14714
rect 10448 14662 10500 14714
rect 10512 14662 10564 14714
rect 10576 14662 10628 14714
rect 14068 14662 14120 14714
rect 14132 14662 14184 14714
rect 14196 14662 14248 14714
rect 14260 14662 14312 14714
rect 14324 14662 14376 14714
rect 4698 14118 4750 14170
rect 4762 14118 4814 14170
rect 4826 14118 4878 14170
rect 4890 14118 4942 14170
rect 4954 14118 5006 14170
rect 8446 14118 8498 14170
rect 8510 14118 8562 14170
rect 8574 14118 8626 14170
rect 8638 14118 8690 14170
rect 8702 14118 8754 14170
rect 12194 14118 12246 14170
rect 12258 14118 12310 14170
rect 12322 14118 12374 14170
rect 12386 14118 12438 14170
rect 12450 14118 12502 14170
rect 1216 14016 1268 14068
rect 9588 13880 9640 13932
rect 3516 13812 3568 13864
rect 2824 13574 2876 13626
rect 2888 13574 2940 13626
rect 2952 13574 3004 13626
rect 3016 13574 3068 13626
rect 3080 13574 3132 13626
rect 6572 13574 6624 13626
rect 6636 13574 6688 13626
rect 6700 13574 6752 13626
rect 6764 13574 6816 13626
rect 6828 13574 6880 13626
rect 10320 13574 10372 13626
rect 10384 13574 10436 13626
rect 10448 13574 10500 13626
rect 10512 13574 10564 13626
rect 10576 13574 10628 13626
rect 14068 13574 14120 13626
rect 14132 13574 14184 13626
rect 14196 13574 14248 13626
rect 14260 13574 14312 13626
rect 14324 13574 14376 13626
rect 4698 13030 4750 13082
rect 4762 13030 4814 13082
rect 4826 13030 4878 13082
rect 4890 13030 4942 13082
rect 4954 13030 5006 13082
rect 8446 13030 8498 13082
rect 8510 13030 8562 13082
rect 8574 13030 8626 13082
rect 8638 13030 8690 13082
rect 8702 13030 8754 13082
rect 12194 13030 12246 13082
rect 12258 13030 12310 13082
rect 12322 13030 12374 13082
rect 12386 13030 12438 13082
rect 12450 13030 12502 13082
rect 4160 12971 4212 12980
rect 4160 12937 4169 12971
rect 4169 12937 4203 12971
rect 4203 12937 4212 12971
rect 4160 12928 4212 12937
rect 5908 12971 5960 12980
rect 5908 12937 5917 12971
rect 5917 12937 5951 12971
rect 5951 12937 5960 12971
rect 5908 12928 5960 12937
rect 13728 12928 13780 12980
rect 4344 12767 4396 12776
rect 4344 12733 4353 12767
rect 4353 12733 4387 12767
rect 4387 12733 4396 12767
rect 4344 12724 4396 12733
rect 6368 12588 6420 12640
rect 8208 12588 8260 12640
rect 9588 12588 9640 12640
rect 12440 12588 12492 12640
rect 14648 12588 14700 12640
rect 2824 12486 2876 12538
rect 2888 12486 2940 12538
rect 2952 12486 3004 12538
rect 3016 12486 3068 12538
rect 3080 12486 3132 12538
rect 6572 12486 6624 12538
rect 6636 12486 6688 12538
rect 6700 12486 6752 12538
rect 6764 12486 6816 12538
rect 6828 12486 6880 12538
rect 10320 12486 10372 12538
rect 10384 12486 10436 12538
rect 10448 12486 10500 12538
rect 10512 12486 10564 12538
rect 10576 12486 10628 12538
rect 14068 12486 14120 12538
rect 14132 12486 14184 12538
rect 14196 12486 14248 12538
rect 14260 12486 14312 12538
rect 14324 12486 14376 12538
rect 4068 12384 4120 12436
rect 7472 12427 7524 12436
rect 7472 12393 7481 12427
rect 7481 12393 7515 12427
rect 7515 12393 7524 12427
rect 7472 12384 7524 12393
rect 8300 12384 8352 12436
rect 8944 12384 8996 12436
rect 9404 12427 9456 12436
rect 9404 12393 9413 12427
rect 9413 12393 9447 12427
rect 9447 12393 9456 12427
rect 9404 12384 9456 12393
rect 3976 12316 4028 12368
rect 7196 12316 7248 12368
rect 10968 12316 11020 12368
rect 9772 12248 9824 12300
rect 9956 12248 10008 12300
rect 7748 12180 7800 12232
rect 9128 12112 9180 12164
rect 5908 12044 5960 12096
rect 7748 12087 7800 12096
rect 7748 12053 7757 12087
rect 7757 12053 7791 12087
rect 7791 12053 7800 12087
rect 7748 12044 7800 12053
rect 7932 12087 7984 12096
rect 7932 12053 7941 12087
rect 7941 12053 7975 12087
rect 7975 12053 7984 12087
rect 7932 12044 7984 12053
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 4698 11942 4750 11994
rect 4762 11942 4814 11994
rect 4826 11942 4878 11994
rect 4890 11942 4942 11994
rect 4954 11942 5006 11994
rect 8446 11942 8498 11994
rect 8510 11942 8562 11994
rect 8574 11942 8626 11994
rect 8638 11942 8690 11994
rect 8702 11942 8754 11994
rect 12194 11942 12246 11994
rect 12258 11942 12310 11994
rect 12322 11942 12374 11994
rect 12386 11942 12438 11994
rect 12450 11942 12502 11994
rect 5356 11840 5408 11892
rect 7656 11883 7708 11892
rect 7656 11849 7665 11883
rect 7665 11849 7699 11883
rect 7699 11849 7708 11883
rect 7656 11840 7708 11849
rect 7564 11704 7616 11756
rect 7932 11704 7984 11756
rect 11888 11840 11940 11892
rect 9956 11772 10008 11824
rect 9128 11704 9180 11756
rect 9312 11636 9364 11688
rect 11244 11568 11296 11620
rect 5724 11500 5776 11552
rect 6184 11500 6236 11552
rect 8116 11543 8168 11552
rect 8116 11509 8125 11543
rect 8125 11509 8159 11543
rect 8159 11509 8168 11543
rect 8116 11500 8168 11509
rect 2824 11398 2876 11450
rect 2888 11398 2940 11450
rect 2952 11398 3004 11450
rect 3016 11398 3068 11450
rect 3080 11398 3132 11450
rect 6572 11398 6624 11450
rect 6636 11398 6688 11450
rect 6700 11398 6752 11450
rect 6764 11398 6816 11450
rect 6828 11398 6880 11450
rect 10320 11398 10372 11450
rect 10384 11398 10436 11450
rect 10448 11398 10500 11450
rect 10512 11398 10564 11450
rect 10576 11398 10628 11450
rect 14068 11398 14120 11450
rect 14132 11398 14184 11450
rect 14196 11398 14248 11450
rect 14260 11398 14312 11450
rect 14324 11398 14376 11450
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 7012 11296 7064 11348
rect 10232 11296 10284 11348
rect 5540 11228 5592 11280
rect 7196 11092 7248 11144
rect 7656 11160 7708 11212
rect 8024 11160 8076 11212
rect 9956 11228 10008 11280
rect 9496 11203 9548 11212
rect 7840 11092 7892 11144
rect 9496 11169 9505 11203
rect 9505 11169 9539 11203
rect 9539 11169 9548 11203
rect 9496 11160 9548 11169
rect 9312 11135 9364 11144
rect 9312 11101 9321 11135
rect 9321 11101 9355 11135
rect 9355 11101 9364 11135
rect 9312 11092 9364 11101
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 11152 11160 11204 11212
rect 9404 11092 9456 11101
rect 9036 11024 9088 11076
rect 9128 11024 9180 11076
rect 6092 10956 6144 11008
rect 6276 10999 6328 11008
rect 6276 10965 6285 10999
rect 6285 10965 6319 10999
rect 6319 10965 6328 10999
rect 6276 10956 6328 10965
rect 7472 10956 7524 11008
rect 8024 10956 8076 11008
rect 4698 10854 4750 10906
rect 4762 10854 4814 10906
rect 4826 10854 4878 10906
rect 4890 10854 4942 10906
rect 4954 10854 5006 10906
rect 8446 10854 8498 10906
rect 8510 10854 8562 10906
rect 8574 10854 8626 10906
rect 8638 10854 8690 10906
rect 8702 10854 8754 10906
rect 12194 10854 12246 10906
rect 12258 10854 12310 10906
rect 12322 10854 12374 10906
rect 12386 10854 12438 10906
rect 12450 10854 12502 10906
rect 4160 10752 4212 10804
rect 5356 10795 5408 10804
rect 5356 10761 5365 10795
rect 5365 10761 5399 10795
rect 5399 10761 5408 10795
rect 5356 10752 5408 10761
rect 5816 10752 5868 10804
rect 7288 10795 7340 10804
rect 7288 10761 7297 10795
rect 7297 10761 7331 10795
rect 7331 10761 7340 10795
rect 7288 10752 7340 10761
rect 8300 10752 8352 10804
rect 9588 10752 9640 10804
rect 4988 10684 5040 10736
rect 9220 10684 9272 10736
rect 3240 10616 3292 10668
rect 3516 10616 3568 10668
rect 6092 10616 6144 10668
rect 6276 10616 6328 10668
rect 6460 10616 6512 10668
rect 6368 10548 6420 10600
rect 7472 10616 7524 10668
rect 8024 10659 8076 10668
rect 8024 10625 8058 10659
rect 8058 10625 8076 10659
rect 8024 10616 8076 10625
rect 9036 10616 9088 10668
rect 9312 10616 9364 10668
rect 10692 10752 10744 10804
rect 11336 10752 11388 10804
rect 13912 10752 13964 10804
rect 12072 10684 12124 10736
rect 15108 10684 15160 10736
rect 5908 10480 5960 10532
rect 7380 10548 7432 10600
rect 10968 10616 11020 10668
rect 13636 10616 13688 10668
rect 11060 10548 11112 10600
rect 11704 10548 11756 10600
rect 14556 10548 14608 10600
rect 2688 10412 2740 10464
rect 5264 10412 5316 10464
rect 8760 10480 8812 10532
rect 9772 10480 9824 10532
rect 10692 10480 10744 10532
rect 6460 10412 6512 10464
rect 7196 10412 7248 10464
rect 8852 10412 8904 10464
rect 9956 10412 10008 10464
rect 10048 10412 10100 10464
rect 12532 10480 12584 10532
rect 2824 10310 2876 10362
rect 2888 10310 2940 10362
rect 2952 10310 3004 10362
rect 3016 10310 3068 10362
rect 3080 10310 3132 10362
rect 6572 10310 6624 10362
rect 6636 10310 6688 10362
rect 6700 10310 6752 10362
rect 6764 10310 6816 10362
rect 6828 10310 6880 10362
rect 10320 10310 10372 10362
rect 10384 10310 10436 10362
rect 10448 10310 10500 10362
rect 10512 10310 10564 10362
rect 10576 10310 10628 10362
rect 14068 10310 14120 10362
rect 14132 10310 14184 10362
rect 14196 10310 14248 10362
rect 14260 10310 14312 10362
rect 14324 10310 14376 10362
rect 5816 10208 5868 10260
rect 8760 10208 8812 10260
rect 9312 10208 9364 10260
rect 9588 10208 9640 10260
rect 10048 10208 10100 10260
rect 10784 10208 10836 10260
rect 3516 10140 3568 10192
rect 8392 10140 8444 10192
rect 5356 10072 5408 10124
rect 4988 10047 5040 10056
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 5540 10004 5592 10056
rect 7196 10047 7248 10056
rect 5264 9936 5316 9988
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 8300 10072 8352 10124
rect 8024 10004 8076 10056
rect 3792 9868 3844 9920
rect 5540 9911 5592 9920
rect 5540 9877 5549 9911
rect 5549 9877 5583 9911
rect 5583 9877 5592 9911
rect 6368 9936 6420 9988
rect 6828 9936 6880 9988
rect 7472 9979 7524 9988
rect 7472 9945 7506 9979
rect 7506 9945 7524 9979
rect 8760 10004 8812 10056
rect 8852 10004 8904 10056
rect 9496 10072 9548 10124
rect 10876 10140 10928 10192
rect 13820 10208 13872 10260
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 10968 10047 11020 10056
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 12072 10047 12124 10056
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 14464 10140 14516 10192
rect 7472 9936 7524 9945
rect 5540 9868 5592 9877
rect 7932 9868 7984 9920
rect 9588 9868 9640 9920
rect 9864 9911 9916 9920
rect 9864 9877 9873 9911
rect 9873 9877 9907 9911
rect 9907 9877 9916 9911
rect 9864 9868 9916 9877
rect 10600 9868 10652 9920
rect 10784 9911 10836 9920
rect 10784 9877 10793 9911
rect 10793 9877 10827 9911
rect 10827 9877 10836 9911
rect 10784 9868 10836 9877
rect 10968 9868 11020 9920
rect 11152 9911 11204 9920
rect 11152 9877 11161 9911
rect 11161 9877 11195 9911
rect 11195 9877 11204 9911
rect 11152 9868 11204 9877
rect 11888 9911 11940 9920
rect 11888 9877 11897 9911
rect 11897 9877 11931 9911
rect 11931 9877 11940 9911
rect 11888 9868 11940 9877
rect 12532 9868 12584 9920
rect 13360 9911 13412 9920
rect 13360 9877 13369 9911
rect 13369 9877 13403 9911
rect 13403 9877 13412 9911
rect 13360 9868 13412 9877
rect 4698 9766 4750 9818
rect 4762 9766 4814 9818
rect 4826 9766 4878 9818
rect 4890 9766 4942 9818
rect 4954 9766 5006 9818
rect 8446 9766 8498 9818
rect 8510 9766 8562 9818
rect 8574 9766 8626 9818
rect 8638 9766 8690 9818
rect 8702 9766 8754 9818
rect 12194 9766 12246 9818
rect 12258 9766 12310 9818
rect 12322 9766 12374 9818
rect 12386 9766 12438 9818
rect 12450 9766 12502 9818
rect 3240 9596 3292 9648
rect 4252 9596 4304 9648
rect 7196 9664 7248 9716
rect 5724 9528 5776 9580
rect 6920 9596 6972 9648
rect 7104 9596 7156 9648
rect 7748 9596 7800 9648
rect 1492 9503 1544 9512
rect 1492 9469 1501 9503
rect 1501 9469 1535 9503
rect 1535 9469 1544 9503
rect 1492 9460 1544 9469
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 5356 9460 5408 9512
rect 7472 9528 7524 9580
rect 8392 9664 8444 9716
rect 8944 9664 8996 9716
rect 9496 9664 9548 9716
rect 8576 9596 8628 9648
rect 8668 9596 8720 9648
rect 10232 9596 10284 9648
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 9496 9571 9548 9580
rect 9496 9537 9505 9571
rect 9505 9537 9539 9571
rect 9539 9537 9548 9571
rect 9496 9528 9548 9537
rect 8300 9503 8352 9512
rect 8300 9469 8302 9503
rect 8302 9469 8336 9503
rect 8336 9469 8352 9503
rect 8300 9460 8352 9469
rect 8576 9460 8628 9512
rect 9036 9503 9088 9512
rect 3424 9392 3476 9444
rect 1676 9324 1728 9376
rect 5632 9367 5684 9376
rect 5632 9333 5641 9367
rect 5641 9333 5675 9367
rect 5675 9333 5684 9367
rect 5632 9324 5684 9333
rect 8392 9435 8444 9444
rect 8392 9401 8401 9435
rect 8401 9401 8435 9435
rect 8435 9401 8444 9435
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 9404 9460 9456 9512
rect 9772 9528 9824 9580
rect 10048 9528 10100 9580
rect 13544 9596 13596 9648
rect 9680 9460 9732 9512
rect 11796 9528 11848 9580
rect 12992 9528 13044 9580
rect 8392 9392 8444 9401
rect 11980 9392 12032 9444
rect 12624 9392 12676 9444
rect 15108 9392 15160 9444
rect 7104 9324 7156 9376
rect 9128 9324 9180 9376
rect 9588 9324 9640 9376
rect 9772 9324 9824 9376
rect 10324 9324 10376 9376
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 11612 9367 11664 9376
rect 11612 9333 11621 9367
rect 11621 9333 11655 9367
rect 11655 9333 11664 9367
rect 11612 9324 11664 9333
rect 11796 9367 11848 9376
rect 11796 9333 11805 9367
rect 11805 9333 11839 9367
rect 11839 9333 11848 9367
rect 11796 9324 11848 9333
rect 12992 9367 13044 9376
rect 12992 9333 13001 9367
rect 13001 9333 13035 9367
rect 13035 9333 13044 9367
rect 12992 9324 13044 9333
rect 2824 9222 2876 9274
rect 2888 9222 2940 9274
rect 2952 9222 3004 9274
rect 3016 9222 3068 9274
rect 3080 9222 3132 9274
rect 6572 9222 6624 9274
rect 6636 9222 6688 9274
rect 6700 9222 6752 9274
rect 6764 9222 6816 9274
rect 6828 9222 6880 9274
rect 10320 9222 10372 9274
rect 10384 9222 10436 9274
rect 10448 9222 10500 9274
rect 10512 9222 10564 9274
rect 10576 9222 10628 9274
rect 14068 9222 14120 9274
rect 14132 9222 14184 9274
rect 14196 9222 14248 9274
rect 14260 9222 14312 9274
rect 14324 9222 14376 9274
rect 5356 9120 5408 9172
rect 6000 9163 6052 9172
rect 6000 9129 6009 9163
rect 6009 9129 6043 9163
rect 6043 9129 6052 9163
rect 6000 9120 6052 9129
rect 4344 9052 4396 9104
rect 7196 9120 7248 9172
rect 8024 9120 8076 9172
rect 8760 9120 8812 9172
rect 9128 9120 9180 9172
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 7840 9052 7892 9104
rect 11888 9052 11940 9104
rect 6920 8916 6972 8968
rect 7104 8959 7156 8968
rect 7104 8925 7138 8959
rect 7138 8925 7156 8959
rect 7104 8916 7156 8925
rect 7472 8916 7524 8968
rect 9312 8984 9364 9036
rect 9496 8984 9548 9036
rect 12808 8984 12860 9036
rect 8208 8916 8260 8968
rect 8392 8916 8444 8968
rect 4620 8848 4672 8900
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 3148 8780 3200 8832
rect 5724 8780 5776 8832
rect 5908 8848 5960 8900
rect 8576 8848 8628 8900
rect 10140 8916 10192 8968
rect 9680 8848 9732 8900
rect 10232 8848 10284 8900
rect 9036 8823 9088 8832
rect 9036 8789 9045 8823
rect 9045 8789 9079 8823
rect 9079 8789 9088 8823
rect 9036 8780 9088 8789
rect 10048 8823 10100 8832
rect 10048 8789 10057 8823
rect 10057 8789 10091 8823
rect 10091 8789 10100 8823
rect 10048 8780 10100 8789
rect 4698 8678 4750 8730
rect 4762 8678 4814 8730
rect 4826 8678 4878 8730
rect 4890 8678 4942 8730
rect 4954 8678 5006 8730
rect 8446 8678 8498 8730
rect 8510 8678 8562 8730
rect 8574 8678 8626 8730
rect 8638 8678 8690 8730
rect 8702 8678 8754 8730
rect 12194 8678 12246 8730
rect 12258 8678 12310 8730
rect 12322 8678 12374 8730
rect 12386 8678 12438 8730
rect 12450 8678 12502 8730
rect 5540 8576 5592 8628
rect 8208 8576 8260 8628
rect 9680 8576 9732 8628
rect 8300 8508 8352 8560
rect 7104 8372 7156 8424
rect 7656 8415 7708 8424
rect 7656 8381 7665 8415
rect 7665 8381 7699 8415
rect 7699 8381 7708 8415
rect 7656 8372 7708 8381
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 9864 8440 9916 8492
rect 8852 8372 8904 8424
rect 12716 8347 12768 8356
rect 12716 8313 12725 8347
rect 12725 8313 12759 8347
rect 12759 8313 12768 8347
rect 12716 8304 12768 8313
rect 8392 8236 8444 8288
rect 9496 8236 9548 8288
rect 2824 8134 2876 8186
rect 2888 8134 2940 8186
rect 2952 8134 3004 8186
rect 3016 8134 3068 8186
rect 3080 8134 3132 8186
rect 6572 8134 6624 8186
rect 6636 8134 6688 8186
rect 6700 8134 6752 8186
rect 6764 8134 6816 8186
rect 6828 8134 6880 8186
rect 10320 8134 10372 8186
rect 10384 8134 10436 8186
rect 10448 8134 10500 8186
rect 10512 8134 10564 8186
rect 10576 8134 10628 8186
rect 14068 8134 14120 8186
rect 14132 8134 14184 8186
rect 14196 8134 14248 8186
rect 14260 8134 14312 8186
rect 14324 8134 14376 8186
rect 5080 7896 5132 7948
rect 7288 7896 7340 7948
rect 4698 7590 4750 7642
rect 4762 7590 4814 7642
rect 4826 7590 4878 7642
rect 4890 7590 4942 7642
rect 4954 7590 5006 7642
rect 8446 7590 8498 7642
rect 8510 7590 8562 7642
rect 8574 7590 8626 7642
rect 8638 7590 8690 7642
rect 8702 7590 8754 7642
rect 12194 7590 12246 7642
rect 12258 7590 12310 7642
rect 12322 7590 12374 7642
rect 12386 7590 12438 7642
rect 12450 7590 12502 7642
rect 3332 7488 3384 7540
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 5080 7420 5132 7472
rect 7748 7488 7800 7540
rect 7932 7488 7984 7540
rect 9404 7488 9456 7540
rect 3240 7327 3292 7336
rect 3240 7293 3249 7327
rect 3249 7293 3283 7327
rect 3283 7293 3292 7327
rect 3240 7284 3292 7293
rect 9128 7284 9180 7336
rect 5080 7216 5132 7268
rect 4620 7191 4672 7200
rect 4620 7157 4629 7191
rect 4629 7157 4663 7191
rect 4663 7157 4672 7191
rect 4620 7148 4672 7157
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 7288 7216 7340 7268
rect 2824 7046 2876 7098
rect 2888 7046 2940 7098
rect 2952 7046 3004 7098
rect 3016 7046 3068 7098
rect 3080 7046 3132 7098
rect 6572 7046 6624 7098
rect 6636 7046 6688 7098
rect 6700 7046 6752 7098
rect 6764 7046 6816 7098
rect 6828 7046 6880 7098
rect 10320 7046 10372 7098
rect 10384 7046 10436 7098
rect 10448 7046 10500 7098
rect 10512 7046 10564 7098
rect 10576 7046 10628 7098
rect 14068 7046 14120 7098
rect 14132 7046 14184 7098
rect 14196 7046 14248 7098
rect 14260 7046 14312 7098
rect 14324 7046 14376 7098
rect 4698 6502 4750 6554
rect 4762 6502 4814 6554
rect 4826 6502 4878 6554
rect 4890 6502 4942 6554
rect 4954 6502 5006 6554
rect 8446 6502 8498 6554
rect 8510 6502 8562 6554
rect 8574 6502 8626 6554
rect 8638 6502 8690 6554
rect 8702 6502 8754 6554
rect 12194 6502 12246 6554
rect 12258 6502 12310 6554
rect 12322 6502 12374 6554
rect 12386 6502 12438 6554
rect 12450 6502 12502 6554
rect 2824 5958 2876 6010
rect 2888 5958 2940 6010
rect 2952 5958 3004 6010
rect 3016 5958 3068 6010
rect 3080 5958 3132 6010
rect 6572 5958 6624 6010
rect 6636 5958 6688 6010
rect 6700 5958 6752 6010
rect 6764 5958 6816 6010
rect 6828 5958 6880 6010
rect 10320 5958 10372 6010
rect 10384 5958 10436 6010
rect 10448 5958 10500 6010
rect 10512 5958 10564 6010
rect 10576 5958 10628 6010
rect 14068 5958 14120 6010
rect 14132 5958 14184 6010
rect 14196 5958 14248 6010
rect 14260 5958 14312 6010
rect 14324 5958 14376 6010
rect 4698 5414 4750 5466
rect 4762 5414 4814 5466
rect 4826 5414 4878 5466
rect 4890 5414 4942 5466
rect 4954 5414 5006 5466
rect 8446 5414 8498 5466
rect 8510 5414 8562 5466
rect 8574 5414 8626 5466
rect 8638 5414 8690 5466
rect 8702 5414 8754 5466
rect 12194 5414 12246 5466
rect 12258 5414 12310 5466
rect 12322 5414 12374 5466
rect 12386 5414 12438 5466
rect 12450 5414 12502 5466
rect 2824 4870 2876 4922
rect 2888 4870 2940 4922
rect 2952 4870 3004 4922
rect 3016 4870 3068 4922
rect 3080 4870 3132 4922
rect 6572 4870 6624 4922
rect 6636 4870 6688 4922
rect 6700 4870 6752 4922
rect 6764 4870 6816 4922
rect 6828 4870 6880 4922
rect 10320 4870 10372 4922
rect 10384 4870 10436 4922
rect 10448 4870 10500 4922
rect 10512 4870 10564 4922
rect 10576 4870 10628 4922
rect 14068 4870 14120 4922
rect 14132 4870 14184 4922
rect 14196 4870 14248 4922
rect 14260 4870 14312 4922
rect 14324 4870 14376 4922
rect 4698 4326 4750 4378
rect 4762 4326 4814 4378
rect 4826 4326 4878 4378
rect 4890 4326 4942 4378
rect 4954 4326 5006 4378
rect 8446 4326 8498 4378
rect 8510 4326 8562 4378
rect 8574 4326 8626 4378
rect 8638 4326 8690 4378
rect 8702 4326 8754 4378
rect 12194 4326 12246 4378
rect 12258 4326 12310 4378
rect 12322 4326 12374 4378
rect 12386 4326 12438 4378
rect 12450 4326 12502 4378
rect 3976 4088 4028 4140
rect 6460 4088 6512 4140
rect 7380 4088 7432 4140
rect 8852 4088 8904 4140
rect 9680 4088 9732 4140
rect 12072 4088 12124 4140
rect 12992 4088 13044 4140
rect 15752 4088 15804 4140
rect 5724 4020 5776 4072
rect 9128 4020 9180 4072
rect 9312 4020 9364 4072
rect 11704 4020 11756 4072
rect 13360 4020 13412 4072
rect 15016 4020 15068 4072
rect 3608 3952 3660 4004
rect 7012 3952 7064 4004
rect 8300 3952 8352 4004
rect 10968 3952 11020 4004
rect 4344 3884 4396 3936
rect 8116 3884 8168 3936
rect 2824 3782 2876 3834
rect 2888 3782 2940 3834
rect 2952 3782 3004 3834
rect 3016 3782 3068 3834
rect 3080 3782 3132 3834
rect 6572 3782 6624 3834
rect 6636 3782 6688 3834
rect 6700 3782 6752 3834
rect 6764 3782 6816 3834
rect 6828 3782 6880 3834
rect 10320 3782 10372 3834
rect 10384 3782 10436 3834
rect 10448 3782 10500 3834
rect 10512 3782 10564 3834
rect 10576 3782 10628 3834
rect 14068 3782 14120 3834
rect 14132 3782 14184 3834
rect 14196 3782 14248 3834
rect 14260 3782 14312 3834
rect 14324 3782 14376 3834
rect 1400 3680 1452 3732
rect 4620 3680 4672 3732
rect 6092 3680 6144 3732
rect 9864 3680 9916 3732
rect 11796 3680 11848 3732
rect 13912 3680 13964 3732
rect 10692 3612 10744 3664
rect 14648 3612 14700 3664
rect 4620 3544 4672 3596
rect 9036 3544 9088 3596
rect 9496 3544 9548 3596
rect 12532 3544 12584 3596
rect 2136 3476 2188 3528
rect 5172 3476 5224 3528
rect 7564 3476 7616 3528
rect 10968 3476 11020 3528
rect 1768 3408 1820 3460
rect 3792 3408 3844 3460
rect 6920 3408 6972 3460
rect 10876 3408 10928 3460
rect 11612 3408 11664 3460
rect 13820 3408 13872 3460
rect 10048 3340 10100 3392
rect 13176 3340 13228 3392
rect 4698 3238 4750 3290
rect 4762 3238 4814 3290
rect 4826 3238 4878 3290
rect 4890 3238 4942 3290
rect 4954 3238 5006 3290
rect 8446 3238 8498 3290
rect 8510 3238 8562 3290
rect 8574 3238 8626 3290
rect 8638 3238 8690 3290
rect 8702 3238 8754 3290
rect 12194 3238 12246 3290
rect 12258 3238 12310 3290
rect 12322 3238 12374 3290
rect 12386 3238 12438 3290
rect 12450 3238 12502 3290
rect 6276 3136 6328 3188
rect 10692 3136 10744 3188
rect 2504 3068 2556 3120
rect 5632 3068 5684 3120
rect 6184 3068 6236 3120
rect 10784 3068 10836 3120
rect 5816 2796 5868 2848
rect 9956 2796 10008 2848
rect 2824 2694 2876 2746
rect 2888 2694 2940 2746
rect 2952 2694 3004 2746
rect 3016 2694 3068 2746
rect 3080 2694 3132 2746
rect 6572 2694 6624 2746
rect 6636 2694 6688 2746
rect 6700 2694 6752 2746
rect 6764 2694 6816 2746
rect 6828 2694 6880 2746
rect 10320 2694 10372 2746
rect 10384 2694 10436 2746
rect 10448 2694 10500 2746
rect 10512 2694 10564 2746
rect 10576 2694 10628 2746
rect 14068 2694 14120 2746
rect 14132 2694 14184 2746
rect 14196 2694 14248 2746
rect 14260 2694 14312 2746
rect 14324 2694 14376 2746
rect 2872 2592 2924 2644
rect 3332 2592 3384 2644
rect 6368 2592 6420 2644
rect 12440 2592 12492 2644
rect 4698 2150 4750 2202
rect 4762 2150 4814 2202
rect 4826 2150 4878 2202
rect 4890 2150 4942 2202
rect 4954 2150 5006 2202
rect 8446 2150 8498 2202
rect 8510 2150 8562 2202
rect 8574 2150 8626 2202
rect 8638 2150 8690 2202
rect 8702 2150 8754 2202
rect 12194 2150 12246 2202
rect 12258 2150 12310 2202
rect 12322 2150 12374 2202
rect 12386 2150 12438 2202
rect 12450 2150 12502 2202
<< metal2 >>
rect 1214 19200 1270 20000
rect 1582 19200 1638 20000
rect 1688 19230 1900 19258
rect 1228 14074 1256 19200
rect 1596 15366 1624 19200
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1216 14068 1268 14074
rect 1216 14010 1268 14016
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1504 8838 1532 9454
rect 1688 9382 1716 19230
rect 1872 19122 1900 19230
rect 1950 19200 2006 20000
rect 2318 19200 2374 20000
rect 2686 19200 2742 20000
rect 3054 19200 3110 20000
rect 3422 19200 3478 20000
rect 3790 19200 3846 20000
rect 4158 19200 4214 20000
rect 4264 19230 4476 19258
rect 1964 19122 1992 19200
rect 1872 19094 1992 19122
rect 2332 15502 2360 19200
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 1766 14920 1822 14929
rect 1766 14855 1822 14864
rect 1780 9518 1808 14855
rect 2700 10470 2728 19200
rect 3068 17898 3096 19200
rect 3068 17870 3188 17898
rect 2824 16892 3132 16901
rect 2824 16890 2830 16892
rect 2886 16890 2910 16892
rect 2966 16890 2990 16892
rect 3046 16890 3070 16892
rect 3126 16890 3132 16892
rect 2886 16838 2888 16890
rect 3068 16838 3070 16890
rect 2824 16836 2830 16838
rect 2886 16836 2910 16838
rect 2966 16836 2990 16838
rect 3046 16836 3070 16838
rect 3126 16836 3132 16838
rect 2824 16827 3132 16836
rect 2824 15804 3132 15813
rect 2824 15802 2830 15804
rect 2886 15802 2910 15804
rect 2966 15802 2990 15804
rect 3046 15802 3070 15804
rect 3126 15802 3132 15804
rect 2886 15750 2888 15802
rect 3068 15750 3070 15802
rect 2824 15748 2830 15750
rect 2886 15748 2910 15750
rect 2966 15748 2990 15750
rect 3046 15748 3070 15750
rect 3126 15748 3132 15750
rect 2824 15739 3132 15748
rect 3160 15434 3188 17870
rect 3436 15570 3464 19200
rect 3804 16046 3832 19200
rect 4066 18184 4122 18193
rect 4066 18119 4122 18128
rect 4080 17762 4108 18119
rect 4172 17950 4200 19200
rect 4160 17944 4212 17950
rect 4160 17886 4212 17892
rect 4080 17734 4200 17762
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 2824 14716 3132 14725
rect 2824 14714 2830 14716
rect 2886 14714 2910 14716
rect 2966 14714 2990 14716
rect 3046 14714 3070 14716
rect 3126 14714 3132 14716
rect 2886 14662 2888 14714
rect 3068 14662 3070 14714
rect 2824 14660 2830 14662
rect 2886 14660 2910 14662
rect 2966 14660 2990 14662
rect 3046 14660 3070 14662
rect 3126 14660 3132 14662
rect 2824 14651 3132 14660
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 2824 13628 3132 13637
rect 2824 13626 2830 13628
rect 2886 13626 2910 13628
rect 2966 13626 2990 13628
rect 3046 13626 3070 13628
rect 3126 13626 3132 13628
rect 2886 13574 2888 13626
rect 3068 13574 3070 13626
rect 2824 13572 2830 13574
rect 2886 13572 2910 13574
rect 2966 13572 2990 13574
rect 3046 13572 3070 13574
rect 3126 13572 3132 13574
rect 2824 13563 3132 13572
rect 2824 12540 3132 12549
rect 2824 12538 2830 12540
rect 2886 12538 2910 12540
rect 2966 12538 2990 12540
rect 3046 12538 3070 12540
rect 3126 12538 3132 12540
rect 2886 12486 2888 12538
rect 3068 12486 3070 12538
rect 2824 12484 2830 12486
rect 2886 12484 2910 12486
rect 2966 12484 2990 12486
rect 3046 12484 3070 12486
rect 3126 12484 3132 12486
rect 2824 12475 3132 12484
rect 2824 11452 3132 11461
rect 2824 11450 2830 11452
rect 2886 11450 2910 11452
rect 2966 11450 2990 11452
rect 3046 11450 3070 11452
rect 3126 11450 3132 11452
rect 2886 11398 2888 11450
rect 3068 11398 3070 11450
rect 2824 11396 2830 11398
rect 2886 11396 2910 11398
rect 2966 11396 2990 11398
rect 3046 11396 3070 11398
rect 3126 11396 3132 11398
rect 2824 11387 3132 11396
rect 3528 10674 3556 13806
rect 3988 12374 4016 15438
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 4080 12442 4108 15302
rect 4172 12986 4200 17734
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 4158 11656 4214 11665
rect 4158 11591 4214 11600
rect 4172 10810 4200 11591
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2824 10364 3132 10373
rect 2824 10362 2830 10364
rect 2886 10362 2910 10364
rect 2966 10362 2990 10364
rect 3046 10362 3070 10364
rect 3126 10362 3132 10364
rect 2886 10310 2888 10362
rect 3068 10310 3070 10362
rect 2824 10308 2830 10310
rect 2886 10308 2910 10310
rect 2966 10308 2990 10310
rect 3046 10308 3070 10310
rect 3126 10308 3132 10310
rect 2824 10299 3132 10308
rect 3252 9654 3280 10610
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 2824 9276 3132 9285
rect 2824 9274 2830 9276
rect 2886 9274 2910 9276
rect 2966 9274 2990 9276
rect 3046 9274 3070 9276
rect 3126 9274 3132 9276
rect 2886 9222 2888 9274
rect 3068 9222 3070 9274
rect 2824 9220 2830 9222
rect 2886 9220 2910 9222
rect 2966 9220 2990 9222
rect 3046 9220 3070 9222
rect 3126 9220 3132 9222
rect 2824 9211 3132 9220
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 2824 8188 3132 8197
rect 2824 8186 2830 8188
rect 2886 8186 2910 8188
rect 2966 8186 2990 8188
rect 3046 8186 3070 8188
rect 3126 8186 3132 8188
rect 2886 8134 2888 8186
rect 3068 8134 3070 8186
rect 2824 8132 2830 8134
rect 2886 8132 2910 8134
rect 2966 8132 2990 8134
rect 3046 8132 3070 8134
rect 3126 8132 3132 8134
rect 2824 8123 3132 8132
rect 2824 7100 3132 7109
rect 2824 7098 2830 7100
rect 2886 7098 2910 7100
rect 2966 7098 2990 7100
rect 3046 7098 3070 7100
rect 3126 7098 3132 7100
rect 2886 7046 2888 7098
rect 3068 7046 3070 7098
rect 2824 7044 2830 7046
rect 2886 7044 2910 7046
rect 2966 7044 2990 7046
rect 3046 7044 3070 7046
rect 3126 7044 3132 7046
rect 2824 7035 3132 7044
rect 2824 6012 3132 6021
rect 2824 6010 2830 6012
rect 2886 6010 2910 6012
rect 2966 6010 2990 6012
rect 3046 6010 3070 6012
rect 3126 6010 3132 6012
rect 2886 5958 2888 6010
rect 3068 5958 3070 6010
rect 2824 5956 2830 5958
rect 2886 5956 2910 5958
rect 2966 5956 2990 5958
rect 3046 5956 3070 5958
rect 3126 5956 3132 5958
rect 2824 5947 3132 5956
rect 2824 4924 3132 4933
rect 2824 4922 2830 4924
rect 2886 4922 2910 4924
rect 2966 4922 2990 4924
rect 3046 4922 3070 4924
rect 3126 4922 3132 4924
rect 2886 4870 2888 4922
rect 3068 4870 3070 4922
rect 2824 4868 2830 4870
rect 2886 4868 2910 4870
rect 2966 4868 2990 4870
rect 3046 4868 3070 4870
rect 3126 4868 3132 4870
rect 2824 4859 3132 4868
rect 2824 3836 3132 3845
rect 2824 3834 2830 3836
rect 2886 3834 2910 3836
rect 2966 3834 2990 3836
rect 3046 3834 3070 3836
rect 3126 3834 3132 3836
rect 2886 3782 2888 3834
rect 3068 3782 3070 3834
rect 2824 3780 2830 3782
rect 2886 3780 2910 3782
rect 2966 3780 2990 3782
rect 3046 3780 3070 3782
rect 3126 3780 3132 3782
rect 2824 3771 3132 3780
rect 1400 3732 1452 3738
rect 1400 3674 1452 3680
rect 1412 800 1440 3674
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 1768 3460 1820 3466
rect 1768 3402 1820 3408
rect 1780 800 1808 3402
rect 2148 800 2176 3470
rect 2504 3120 2556 3126
rect 2504 3062 2556 3068
rect 2516 800 2544 3062
rect 2824 2748 3132 2757
rect 2824 2746 2830 2748
rect 2886 2746 2910 2748
rect 2966 2746 2990 2748
rect 3046 2746 3070 2748
rect 3126 2746 3132 2748
rect 2886 2694 2888 2746
rect 3068 2694 3070 2746
rect 2824 2692 2830 2694
rect 2886 2692 2910 2694
rect 2966 2692 2990 2694
rect 3046 2692 3070 2694
rect 3126 2692 3132 2694
rect 2824 2683 3132 2692
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2884 800 2912 2586
rect 3160 1873 3188 8774
rect 3252 8401 3280 9590
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 3238 8392 3294 8401
rect 3238 8327 3294 8336
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3252 5137 3280 7278
rect 3238 5128 3294 5137
rect 3238 5063 3294 5072
rect 3344 2650 3372 7482
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3436 2530 3464 9386
rect 3528 7410 3556 10134
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3252 2502 3464 2530
rect 3146 1864 3202 1873
rect 3146 1799 3202 1808
rect 3252 800 3280 2502
rect 3620 800 3648 3946
rect 3804 3466 3832 9862
rect 4264 9654 4292 19230
rect 4448 19122 4476 19230
rect 4526 19200 4582 20000
rect 4632 19230 4844 19258
rect 4540 19122 4568 19200
rect 4448 19094 4568 19122
rect 4344 17944 4396 17950
rect 4344 17886 4396 17892
rect 4356 15638 4384 17886
rect 4344 15632 4396 15638
rect 4344 15574 4396 15580
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4356 9110 4384 12718
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4632 8906 4660 19230
rect 4816 19122 4844 19230
rect 4894 19200 4950 20000
rect 5262 19200 5318 20000
rect 5630 19200 5686 20000
rect 5998 19200 6054 20000
rect 6104 19230 6316 19258
rect 4908 19122 4936 19200
rect 4816 19094 4936 19122
rect 4698 17436 5006 17445
rect 4698 17434 4704 17436
rect 4760 17434 4784 17436
rect 4840 17434 4864 17436
rect 4920 17434 4944 17436
rect 5000 17434 5006 17436
rect 4760 17382 4762 17434
rect 4942 17382 4944 17434
rect 4698 17380 4704 17382
rect 4760 17380 4784 17382
rect 4840 17380 4864 17382
rect 4920 17380 4944 17382
rect 5000 17380 5006 17382
rect 4698 17371 5006 17380
rect 4698 16348 5006 16357
rect 4698 16346 4704 16348
rect 4760 16346 4784 16348
rect 4840 16346 4864 16348
rect 4920 16346 4944 16348
rect 5000 16346 5006 16348
rect 4760 16294 4762 16346
rect 4942 16294 4944 16346
rect 4698 16292 4704 16294
rect 4760 16292 4784 16294
rect 4840 16292 4864 16294
rect 4920 16292 4944 16294
rect 5000 16292 5006 16294
rect 4698 16283 5006 16292
rect 5276 15366 5304 19200
rect 5644 16574 5672 19200
rect 5552 16546 5672 16574
rect 5724 16584 5776 16590
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 4698 15260 5006 15269
rect 4698 15258 4704 15260
rect 4760 15258 4784 15260
rect 4840 15258 4864 15260
rect 4920 15258 4944 15260
rect 5000 15258 5006 15260
rect 4760 15206 4762 15258
rect 4942 15206 4944 15258
rect 4698 15204 4704 15206
rect 4760 15204 4784 15206
rect 4840 15204 4864 15206
rect 4920 15204 4944 15206
rect 5000 15204 5006 15206
rect 4698 15195 5006 15204
rect 4698 14172 5006 14181
rect 4698 14170 4704 14172
rect 4760 14170 4784 14172
rect 4840 14170 4864 14172
rect 4920 14170 4944 14172
rect 5000 14170 5006 14172
rect 4760 14118 4762 14170
rect 4942 14118 4944 14170
rect 4698 14116 4704 14118
rect 4760 14116 4784 14118
rect 4840 14116 4864 14118
rect 4920 14116 4944 14118
rect 5000 14116 5006 14118
rect 4698 14107 5006 14116
rect 4698 13084 5006 13093
rect 4698 13082 4704 13084
rect 4760 13082 4784 13084
rect 4840 13082 4864 13084
rect 4920 13082 4944 13084
rect 5000 13082 5006 13084
rect 4760 13030 4762 13082
rect 4942 13030 4944 13082
rect 4698 13028 4704 13030
rect 4760 13028 4784 13030
rect 4840 13028 4864 13030
rect 4920 13028 4944 13030
rect 5000 13028 5006 13030
rect 4698 13019 5006 13028
rect 4698 11996 5006 12005
rect 4698 11994 4704 11996
rect 4760 11994 4784 11996
rect 4840 11994 4864 11996
rect 4920 11994 4944 11996
rect 5000 11994 5006 11996
rect 4760 11942 4762 11994
rect 4942 11942 4944 11994
rect 4698 11940 4704 11942
rect 4760 11940 4784 11942
rect 4840 11940 4864 11942
rect 4920 11940 4944 11942
rect 5000 11940 5006 11942
rect 4698 11931 5006 11940
rect 5368 11898 5396 15982
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5552 11393 5580 16546
rect 5724 16526 5776 16532
rect 5736 16402 5764 16526
rect 5644 16374 5764 16402
rect 5538 11384 5594 11393
rect 5538 11319 5594 11328
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 4698 10908 5006 10917
rect 4698 10906 4704 10908
rect 4760 10906 4784 10908
rect 4840 10906 4864 10908
rect 4920 10906 4944 10908
rect 5000 10906 5006 10908
rect 4760 10854 4762 10906
rect 4942 10854 4944 10906
rect 4698 10852 4704 10854
rect 4760 10852 4784 10854
rect 4840 10852 4864 10854
rect 4920 10852 4944 10854
rect 5000 10852 5006 10854
rect 4698 10843 5006 10852
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 5000 10062 5028 10678
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5276 9994 5304 10406
rect 5368 10130 5396 10746
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5552 10062 5580 11222
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 4698 9820 5006 9829
rect 4698 9818 4704 9820
rect 4760 9818 4784 9820
rect 4840 9818 4864 9820
rect 4920 9818 4944 9820
rect 5000 9818 5006 9820
rect 4760 9766 4762 9818
rect 4942 9766 4944 9818
rect 4698 9764 4704 9766
rect 4760 9764 4784 9766
rect 4840 9764 4864 9766
rect 4920 9764 4944 9766
rect 5000 9764 5006 9766
rect 4698 9755 5006 9764
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5368 9178 5396 9454
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4698 8732 5006 8741
rect 4698 8730 4704 8732
rect 4760 8730 4784 8732
rect 4840 8730 4864 8732
rect 4920 8730 4944 8732
rect 5000 8730 5006 8732
rect 4760 8678 4762 8730
rect 4942 8678 4944 8730
rect 4698 8676 4704 8678
rect 4760 8676 4784 8678
rect 4840 8676 4864 8678
rect 4920 8676 4944 8678
rect 5000 8676 5006 8678
rect 4698 8667 5006 8676
rect 5552 8634 5580 9862
rect 5644 9625 5672 16374
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5736 11558 5764 16050
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5722 11384 5778 11393
rect 5722 11319 5778 11328
rect 5736 10418 5764 11319
rect 5828 10810 5856 15506
rect 5908 15428 5960 15434
rect 5908 15370 5960 15376
rect 5920 12986 5948 15370
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5920 10538 5948 12038
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5736 10390 5948 10418
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5630 9616 5686 9625
rect 5630 9551 5686 9560
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 4698 7644 5006 7653
rect 4698 7642 4704 7644
rect 4760 7642 4784 7644
rect 4840 7642 4864 7644
rect 4920 7642 4944 7644
rect 5000 7642 5006 7644
rect 4760 7590 4762 7642
rect 4942 7590 4944 7642
rect 4698 7588 4704 7590
rect 4760 7588 4784 7590
rect 4840 7588 4864 7590
rect 4920 7588 4944 7590
rect 5000 7588 5006 7590
rect 4698 7579 5006 7588
rect 5092 7478 5120 7890
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 3988 800 4016 4082
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4356 800 4384 3878
rect 4632 3738 4660 7142
rect 4698 6556 5006 6565
rect 4698 6554 4704 6556
rect 4760 6554 4784 6556
rect 4840 6554 4864 6556
rect 4920 6554 4944 6556
rect 5000 6554 5006 6556
rect 4760 6502 4762 6554
rect 4942 6502 4944 6554
rect 4698 6500 4704 6502
rect 4760 6500 4784 6502
rect 4840 6500 4864 6502
rect 4920 6500 4944 6502
rect 5000 6500 5006 6502
rect 4698 6491 5006 6500
rect 4698 5468 5006 5477
rect 4698 5466 4704 5468
rect 4760 5466 4784 5468
rect 4840 5466 4864 5468
rect 4920 5466 4944 5468
rect 5000 5466 5006 5468
rect 4760 5414 4762 5466
rect 4942 5414 4944 5466
rect 4698 5412 4704 5414
rect 4760 5412 4784 5414
rect 4840 5412 4864 5414
rect 4920 5412 4944 5414
rect 5000 5412 5006 5414
rect 4698 5403 5006 5412
rect 4698 4380 5006 4389
rect 4698 4378 4704 4380
rect 4760 4378 4784 4380
rect 4840 4378 4864 4380
rect 4920 4378 4944 4380
rect 5000 4378 5006 4380
rect 4760 4326 4762 4378
rect 4942 4326 4944 4378
rect 4698 4324 4704 4326
rect 4760 4324 4784 4326
rect 4840 4324 4864 4326
rect 4920 4324 4944 4326
rect 5000 4324 5006 4326
rect 4698 4315 5006 4324
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4632 1850 4660 3538
rect 4698 3292 5006 3301
rect 4698 3290 4704 3292
rect 4760 3290 4784 3292
rect 4840 3290 4864 3292
rect 4920 3290 4944 3292
rect 5000 3290 5006 3292
rect 4760 3238 4762 3290
rect 4942 3238 4944 3290
rect 4698 3236 4704 3238
rect 4760 3236 4784 3238
rect 4840 3236 4864 3238
rect 4920 3236 4944 3238
rect 5000 3236 5006 3238
rect 4698 3227 5006 3236
rect 4698 2204 5006 2213
rect 4698 2202 4704 2204
rect 4760 2202 4784 2204
rect 4840 2202 4864 2204
rect 4920 2202 4944 2204
rect 5000 2202 5006 2204
rect 4760 2150 4762 2202
rect 4942 2150 4944 2202
rect 4698 2148 4704 2150
rect 4760 2148 4784 2150
rect 4840 2148 4864 2150
rect 4920 2148 4944 2150
rect 5000 2148 5006 2150
rect 4698 2139 5006 2148
rect 4632 1822 4752 1850
rect 4724 800 4752 1822
rect 5092 800 5120 7210
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 3534 5212 7142
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5644 3126 5672 9318
rect 5736 8838 5764 9522
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5736 4078 5764 8774
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5828 2938 5856 10202
rect 5920 8906 5948 10390
rect 6012 9489 6040 19200
rect 6104 16590 6132 19230
rect 6288 19122 6316 19230
rect 6366 19200 6422 20000
rect 6472 19230 6684 19258
rect 6380 19122 6408 19200
rect 6288 19094 6408 19122
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6472 16114 6500 19230
rect 6656 19122 6684 19230
rect 6734 19200 6790 20000
rect 7102 19200 7158 20000
rect 7470 19200 7526 20000
rect 7838 19200 7894 20000
rect 8206 19200 8262 20000
rect 8574 19200 8630 20000
rect 8680 19230 8892 19258
rect 6748 19122 6776 19200
rect 6656 19094 6776 19122
rect 6572 16892 6880 16901
rect 6572 16890 6578 16892
rect 6634 16890 6658 16892
rect 6714 16890 6738 16892
rect 6794 16890 6818 16892
rect 6874 16890 6880 16892
rect 6634 16838 6636 16890
rect 6816 16838 6818 16890
rect 6572 16836 6578 16838
rect 6634 16836 6658 16838
rect 6714 16836 6738 16838
rect 6794 16836 6818 16838
rect 6874 16836 6880 16838
rect 6572 16827 6880 16836
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6104 10674 6132 10950
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 5998 9480 6054 9489
rect 5998 9415 6054 9424
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6012 8945 6040 9114
rect 5998 8936 6054 8945
rect 5908 8900 5960 8906
rect 5998 8871 6054 8880
rect 5908 8842 5960 8848
rect 6104 3738 6132 10610
rect 6196 9081 6224 11494
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6288 10674 6316 10950
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6182 9072 6238 9081
rect 6182 9007 6238 9016
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6288 3194 6316 10610
rect 6380 10606 6408 12582
rect 6472 11354 6500 15914
rect 6572 15804 6880 15813
rect 6572 15802 6578 15804
rect 6634 15802 6658 15804
rect 6714 15802 6738 15804
rect 6794 15802 6818 15804
rect 6874 15802 6880 15804
rect 6634 15750 6636 15802
rect 6816 15750 6818 15802
rect 6572 15748 6578 15750
rect 6634 15748 6658 15750
rect 6714 15748 6738 15750
rect 6794 15748 6818 15750
rect 6874 15748 6880 15750
rect 6572 15739 6880 15748
rect 7116 15706 7144 19200
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 6572 14716 6880 14725
rect 6572 14714 6578 14716
rect 6634 14714 6658 14716
rect 6714 14714 6738 14716
rect 6794 14714 6818 14716
rect 6874 14714 6880 14716
rect 6634 14662 6636 14714
rect 6816 14662 6818 14714
rect 6572 14660 6578 14662
rect 6634 14660 6658 14662
rect 6714 14660 6738 14662
rect 6794 14660 6818 14662
rect 6874 14660 6880 14662
rect 6572 14651 6880 14660
rect 6572 13628 6880 13637
rect 6572 13626 6578 13628
rect 6634 13626 6658 13628
rect 6714 13626 6738 13628
rect 6794 13626 6818 13628
rect 6874 13626 6880 13628
rect 6634 13574 6636 13626
rect 6816 13574 6818 13626
rect 6572 13572 6578 13574
rect 6634 13572 6658 13574
rect 6714 13572 6738 13574
rect 6794 13572 6818 13574
rect 6874 13572 6880 13574
rect 6572 13563 6880 13572
rect 6572 12540 6880 12549
rect 6572 12538 6578 12540
rect 6634 12538 6658 12540
rect 6714 12538 6738 12540
rect 6794 12538 6818 12540
rect 6874 12538 6880 12540
rect 6634 12486 6636 12538
rect 6816 12486 6818 12538
rect 6572 12484 6578 12486
rect 6634 12484 6658 12486
rect 6714 12484 6738 12486
rect 6794 12484 6818 12486
rect 6874 12484 6880 12486
rect 6572 12475 6880 12484
rect 7208 12434 7236 15846
rect 7484 15502 7512 19200
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7484 12442 7512 15302
rect 7116 12406 7236 12434
rect 7472 12436 7524 12442
rect 6572 11452 6880 11461
rect 6572 11450 6578 11452
rect 6634 11450 6658 11452
rect 6714 11450 6738 11452
rect 6794 11450 6818 11452
rect 6874 11450 6880 11452
rect 6634 11398 6636 11450
rect 6816 11398 6818 11450
rect 6572 11396 6578 11398
rect 6634 11396 6658 11398
rect 6714 11396 6738 11398
rect 6794 11396 6818 11398
rect 6874 11396 6880 11398
rect 6572 11387 6880 11396
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6472 10674 6500 11290
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 5460 2910 5856 2938
rect 5460 800 5488 2910
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5828 800 5856 2790
rect 6196 800 6224 3062
rect 6380 2650 6408 9930
rect 6472 4146 6500 10406
rect 6572 10364 6880 10373
rect 6572 10362 6578 10364
rect 6634 10362 6658 10364
rect 6714 10362 6738 10364
rect 6794 10362 6818 10364
rect 6874 10362 6880 10364
rect 6634 10310 6636 10362
rect 6816 10310 6818 10362
rect 6572 10308 6578 10310
rect 6634 10308 6658 10310
rect 6714 10308 6738 10310
rect 6794 10308 6818 10310
rect 6874 10308 6880 10310
rect 6572 10299 6880 10308
rect 6826 10024 6882 10033
rect 6826 9959 6828 9968
rect 6880 9959 6882 9968
rect 6828 9930 6880 9936
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6572 9276 6880 9285
rect 6572 9274 6578 9276
rect 6634 9274 6658 9276
rect 6714 9274 6738 9276
rect 6794 9274 6818 9276
rect 6874 9274 6880 9276
rect 6634 9222 6636 9274
rect 6816 9222 6818 9274
rect 6572 9220 6578 9222
rect 6634 9220 6658 9222
rect 6714 9220 6738 9222
rect 6794 9220 6818 9222
rect 6874 9220 6880 9222
rect 6572 9211 6880 9220
rect 6932 8974 6960 9590
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6572 8188 6880 8197
rect 6572 8186 6578 8188
rect 6634 8186 6658 8188
rect 6714 8186 6738 8188
rect 6794 8186 6818 8188
rect 6874 8186 6880 8188
rect 6634 8134 6636 8186
rect 6816 8134 6818 8186
rect 6572 8132 6578 8134
rect 6634 8132 6658 8134
rect 6714 8132 6738 8134
rect 6794 8132 6818 8134
rect 6874 8132 6880 8134
rect 6572 8123 6880 8132
rect 6572 7100 6880 7109
rect 6572 7098 6578 7100
rect 6634 7098 6658 7100
rect 6714 7098 6738 7100
rect 6794 7098 6818 7100
rect 6874 7098 6880 7100
rect 6634 7046 6636 7098
rect 6816 7046 6818 7098
rect 6572 7044 6578 7046
rect 6634 7044 6658 7046
rect 6714 7044 6738 7046
rect 6794 7044 6818 7046
rect 6874 7044 6880 7046
rect 6572 7035 6880 7044
rect 6572 6012 6880 6021
rect 6572 6010 6578 6012
rect 6634 6010 6658 6012
rect 6714 6010 6738 6012
rect 6794 6010 6818 6012
rect 6874 6010 6880 6012
rect 6634 5958 6636 6010
rect 6816 5958 6818 6010
rect 6572 5956 6578 5958
rect 6634 5956 6658 5958
rect 6714 5956 6738 5958
rect 6794 5956 6818 5958
rect 6874 5956 6880 5958
rect 6572 5947 6880 5956
rect 6572 4924 6880 4933
rect 6572 4922 6578 4924
rect 6634 4922 6658 4924
rect 6714 4922 6738 4924
rect 6794 4922 6818 4924
rect 6874 4922 6880 4924
rect 6634 4870 6636 4922
rect 6816 4870 6818 4922
rect 6572 4868 6578 4870
rect 6634 4868 6658 4870
rect 6714 4868 6738 4870
rect 6794 4868 6818 4870
rect 6874 4868 6880 4870
rect 6572 4859 6880 4868
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 7024 4010 7052 11290
rect 7116 9654 7144 12406
rect 7472 12378 7524 12384
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7208 11150 7236 12310
rect 7668 11898 7696 15574
rect 7852 15434 7880 19200
rect 8220 15638 8248 19200
rect 8588 19122 8616 19200
rect 8680 19122 8708 19230
rect 8588 19094 8708 19122
rect 8446 17436 8754 17445
rect 8446 17434 8452 17436
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8748 17434 8754 17436
rect 8508 17382 8510 17434
rect 8690 17382 8692 17434
rect 8446 17380 8452 17382
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8748 17380 8754 17382
rect 8446 17371 8754 17380
rect 8446 16348 8754 16357
rect 8446 16346 8452 16348
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8748 16346 8754 16348
rect 8508 16294 8510 16346
rect 8690 16294 8692 16346
rect 8446 16292 8452 16294
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8748 16292 8754 16294
rect 8446 16283 8754 16292
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8864 15570 8892 19230
rect 8942 19200 8998 20000
rect 9310 19200 9366 20000
rect 9678 19200 9734 20000
rect 10046 19200 10102 20000
rect 10414 19200 10470 20000
rect 10782 19200 10838 20000
rect 11150 19200 11206 20000
rect 11518 19200 11574 20000
rect 11886 19200 11942 20000
rect 12254 19200 12310 20000
rect 12622 19200 12678 20000
rect 12990 19200 13046 20000
rect 13358 19200 13414 20000
rect 13726 19200 13782 20000
rect 14094 19200 14150 20000
rect 14462 19200 14518 20000
rect 14830 19200 14886 20000
rect 15198 19200 15254 20000
rect 15566 19200 15622 20000
rect 15934 19200 15990 20000
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 8446 15260 8754 15269
rect 8446 15258 8452 15260
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8748 15258 8754 15260
rect 8508 15206 8510 15258
rect 8690 15206 8692 15258
rect 8446 15204 8452 15206
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8748 15204 8754 15206
rect 8446 15195 8754 15204
rect 8446 14172 8754 14181
rect 8446 14170 8452 14172
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8748 14170 8754 14172
rect 8508 14118 8510 14170
rect 8690 14118 8692 14170
rect 8446 14116 8452 14118
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8748 14116 8754 14118
rect 8446 14107 8754 14116
rect 8446 13084 8754 13093
rect 8446 13082 8452 13084
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8748 13082 8754 13084
rect 8508 13030 8510 13082
rect 8690 13030 8692 13082
rect 8446 13028 8452 13030
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8748 13028 8754 13030
rect 8446 13019 8754 13028
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7760 12102 7788 12174
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7208 10062 7236 10406
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 9722 7236 9998
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7116 8974 7144 9318
rect 7208 9178 7236 9658
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7116 8430 7144 8910
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7300 7954 7328 10746
rect 7484 10674 7512 10950
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6572 3836 6880 3845
rect 6572 3834 6578 3836
rect 6634 3834 6658 3836
rect 6714 3834 6738 3836
rect 6794 3834 6818 3836
rect 6874 3834 6880 3836
rect 6634 3782 6636 3834
rect 6816 3782 6818 3834
rect 6572 3780 6578 3782
rect 6634 3780 6658 3782
rect 6714 3780 6738 3782
rect 6794 3780 6818 3782
rect 6874 3780 6880 3782
rect 6572 3771 6880 3780
rect 6458 3632 6514 3641
rect 6458 3567 6514 3576
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6472 1850 6500 3567
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6572 2748 6880 2757
rect 6572 2746 6578 2748
rect 6634 2746 6658 2748
rect 6714 2746 6738 2748
rect 6794 2746 6818 2748
rect 6874 2746 6880 2748
rect 6634 2694 6636 2746
rect 6816 2694 6818 2746
rect 6572 2692 6578 2694
rect 6634 2692 6658 2694
rect 6714 2692 6738 2694
rect 6794 2692 6818 2694
rect 6874 2692 6880 2694
rect 6572 2683 6880 2692
rect 6472 1822 6592 1850
rect 6564 800 6592 1822
rect 6932 800 6960 3402
rect 7300 800 7328 7210
rect 7392 4146 7420 10542
rect 7484 9994 7512 10610
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7484 8974 7512 9522
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7576 3534 7604 11698
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7668 8430 7696 11154
rect 7760 10169 7788 12038
rect 7944 11762 7972 12038
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7746 10160 7802 10169
rect 7746 10095 7802 10104
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7760 9353 7788 9590
rect 7746 9344 7802 9353
rect 7746 9279 7802 9288
rect 7852 9194 7880 11086
rect 8036 11014 8064 11154
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8036 10062 8064 10610
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7760 9166 7880 9194
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7760 7546 7788 9166
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7852 2774 7880 9046
rect 7944 7546 7972 9862
rect 8036 9178 8064 9998
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 8022 4040 8078 4049
rect 8022 3975 8078 3984
rect 7668 2746 7880 2774
rect 7668 800 7696 2746
rect 8036 800 8064 3975
rect 8128 3942 8156 11494
rect 8220 9217 8248 12582
rect 8956 12442 8984 19200
rect 9324 16574 9352 19200
rect 9232 16546 9352 16574
rect 9692 16574 9720 19200
rect 9692 16546 9812 16574
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 8312 10810 8340 12378
rect 8446 11996 8754 12005
rect 8446 11994 8452 11996
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8748 11994 8754 11996
rect 8508 11942 8510 11994
rect 8690 11942 8692 11994
rect 8446 11940 8452 11942
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8748 11940 8754 11942
rect 8446 11931 8754 11940
rect 9048 11257 9076 15302
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 9140 11762 9168 12106
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9034 11248 9090 11257
rect 9034 11183 9090 11192
rect 9140 11082 9168 11698
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 8446 10908 8754 10917
rect 8446 10906 8452 10908
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8748 10906 8754 10908
rect 8508 10854 8510 10906
rect 8690 10854 8692 10906
rect 8446 10852 8452 10854
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8748 10852 8754 10854
rect 8446 10843 8754 10852
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8312 10130 8340 10746
rect 9048 10674 9076 11018
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8760 10532 8812 10538
rect 8760 10474 8812 10480
rect 8772 10266 8800 10474
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8404 10010 8432 10134
rect 8864 10062 8892 10406
rect 9034 10160 9090 10169
rect 9140 10146 9168 11018
rect 9232 10742 9260 16546
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9416 12442 9444 15438
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9600 12646 9628 13874
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9324 11150 9352 11630
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9324 10266 9352 10610
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9416 10146 9444 11086
rect 9140 10118 9260 10146
rect 9034 10095 9090 10104
rect 8312 9982 8432 10010
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8852 10056 8904 10062
rect 9048 10044 9076 10095
rect 9048 10016 9168 10044
rect 8852 9998 8904 10004
rect 8312 9704 8340 9982
rect 8772 9908 8800 9998
rect 8772 9880 9076 9908
rect 8446 9820 8754 9829
rect 8446 9818 8452 9820
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8748 9818 8754 9820
rect 8508 9766 8510 9818
rect 8690 9766 8692 9818
rect 8446 9764 8452 9766
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8748 9764 8754 9766
rect 8446 9755 8754 9764
rect 8850 9752 8906 9761
rect 8392 9716 8444 9722
rect 8312 9676 8392 9704
rect 8850 9687 8906 9696
rect 8944 9716 8996 9722
rect 8392 9658 8444 9664
rect 8576 9648 8628 9654
rect 8496 9608 8576 9636
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8206 9208 8262 9217
rect 8206 9143 8262 9152
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8220 8634 8248 8910
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8312 8566 8340 9454
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8404 8974 8432 9386
rect 8496 9353 8524 9608
rect 8576 9590 8628 9596
rect 8668 9648 8720 9654
rect 8864 9602 8892 9687
rect 8944 9658 8996 9664
rect 8668 9590 8720 9596
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8482 9344 8538 9353
rect 8482 9279 8538 9288
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8588 8906 8616 9454
rect 8680 9217 8708 9590
rect 8772 9586 8892 9602
rect 8760 9580 8892 9586
rect 8812 9574 8892 9580
rect 8760 9522 8812 9528
rect 8666 9208 8722 9217
rect 8772 9178 8800 9522
rect 8666 9143 8722 9152
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8446 8732 8754 8741
rect 8446 8730 8452 8732
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8748 8730 8754 8732
rect 8508 8678 8510 8730
rect 8690 8678 8692 8730
rect 8446 8676 8452 8678
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8748 8676 8754 8678
rect 8446 8667 8754 8676
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8404 8294 8432 8434
rect 8852 8424 8904 8430
rect 8956 8412 8984 9658
rect 9048 9518 9076 9880
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9140 9382 9168 10016
rect 9128 9376 9180 9382
rect 9034 9344 9090 9353
rect 9128 9318 9180 9324
rect 9034 9279 9090 9288
rect 9048 8945 9076 9279
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9034 8936 9090 8945
rect 9034 8871 9090 8880
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8904 8384 8984 8412
rect 8852 8366 8904 8372
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8446 7644 8754 7653
rect 8446 7642 8452 7644
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8748 7642 8754 7644
rect 8508 7590 8510 7642
rect 8690 7590 8692 7642
rect 8446 7588 8452 7590
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8748 7588 8754 7590
rect 8446 7579 8754 7588
rect 8446 6556 8754 6565
rect 8446 6554 8452 6556
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8748 6554 8754 6556
rect 8508 6502 8510 6554
rect 8690 6502 8692 6554
rect 8446 6500 8452 6502
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8748 6500 8754 6502
rect 8446 6491 8754 6500
rect 8446 5468 8754 5477
rect 8446 5466 8452 5468
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8748 5466 8754 5468
rect 8508 5414 8510 5466
rect 8690 5414 8692 5466
rect 8446 5412 8452 5414
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8748 5412 8754 5414
rect 8446 5403 8754 5412
rect 8446 4380 8754 4389
rect 8446 4378 8452 4380
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8748 4378 8754 4380
rect 8508 4326 8510 4378
rect 8690 4326 8692 4378
rect 8446 4324 8452 4326
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8748 4324 8754 4326
rect 8446 4315 8754 4324
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8312 1986 8340 3946
rect 8446 3292 8754 3301
rect 8446 3290 8452 3292
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8748 3290 8754 3292
rect 8508 3238 8510 3290
rect 8690 3238 8692 3290
rect 8446 3236 8452 3238
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8748 3236 8754 3238
rect 8446 3227 8754 3236
rect 8446 2204 8754 2213
rect 8446 2202 8452 2204
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8748 2202 8754 2204
rect 8508 2150 8510 2202
rect 8690 2150 8692 2202
rect 8446 2148 8452 2150
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8748 2148 8754 2150
rect 8446 2139 8754 2148
rect 8864 1986 8892 4082
rect 9048 3602 9076 8774
rect 9140 7342 9168 9114
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8312 1958 8432 1986
rect 8404 800 8432 1958
rect 8772 1958 8892 1986
rect 8772 800 8800 1958
rect 9140 800 9168 4014
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2134 0 2190 800
rect 2502 0 2558 800
rect 2870 0 2926 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9232 762 9260 10118
rect 9324 10118 9444 10146
rect 9508 10130 9536 11154
rect 9600 10810 9628 12582
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9496 10124 9548 10130
rect 9324 9194 9352 10118
rect 9496 10066 9548 10072
rect 9508 9722 9536 10066
rect 9600 9926 9628 10202
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9353 9444 9454
rect 9402 9344 9458 9353
rect 9402 9279 9458 9288
rect 9324 9166 9444 9194
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9324 4078 9352 8978
rect 9416 7546 9444 9166
rect 9508 9042 9536 9522
rect 9692 9518 9720 15642
rect 9784 12306 9812 16546
rect 10060 12434 10088 19200
rect 10428 17898 10456 19200
rect 10244 17870 10456 17898
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 9876 12406 10088 12434
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9784 10538 9812 12038
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9876 10146 9904 12406
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9968 11830 9996 12242
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 9968 11286 9996 11766
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9784 10118 9904 10146
rect 9784 9586 9812 10118
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9770 9480 9826 9489
rect 9770 9415 9826 9424
rect 9784 9382 9812 9415
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9600 8922 9628 9318
rect 9508 8894 9628 8922
rect 9680 8900 9732 8906
rect 9508 8294 9536 8894
rect 9680 8842 9732 8848
rect 9692 8634 9720 8842
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9508 3602 9536 8230
rect 9692 4146 9720 8570
rect 9876 8498 9904 9862
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9416 870 9536 898
rect 9416 762 9444 870
rect 9508 800 9536 870
rect 9876 800 9904 3674
rect 9968 2854 9996 10406
rect 10060 10266 10088 10406
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10060 8838 10088 9522
rect 10152 9178 10180 15438
rect 10244 15366 10272 17870
rect 10320 16892 10628 16901
rect 10320 16890 10326 16892
rect 10382 16890 10406 16892
rect 10462 16890 10486 16892
rect 10542 16890 10566 16892
rect 10622 16890 10628 16892
rect 10382 16838 10384 16890
rect 10564 16838 10566 16890
rect 10320 16836 10326 16838
rect 10382 16836 10406 16838
rect 10462 16836 10486 16838
rect 10542 16836 10566 16838
rect 10622 16836 10628 16838
rect 10320 16827 10628 16836
rect 10796 15910 10824 19200
rect 11164 16574 11192 19200
rect 10980 16546 11192 16574
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10320 15804 10628 15813
rect 10320 15802 10326 15804
rect 10382 15802 10406 15804
rect 10462 15802 10486 15804
rect 10542 15802 10566 15804
rect 10622 15802 10628 15804
rect 10382 15750 10384 15802
rect 10564 15750 10566 15802
rect 10320 15748 10326 15750
rect 10382 15748 10406 15750
rect 10462 15748 10486 15750
rect 10542 15748 10566 15750
rect 10622 15748 10628 15750
rect 10320 15739 10628 15748
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10320 14716 10628 14725
rect 10320 14714 10326 14716
rect 10382 14714 10406 14716
rect 10462 14714 10486 14716
rect 10542 14714 10566 14716
rect 10622 14714 10628 14716
rect 10382 14662 10384 14714
rect 10564 14662 10566 14714
rect 10320 14660 10326 14662
rect 10382 14660 10406 14662
rect 10462 14660 10486 14662
rect 10542 14660 10566 14662
rect 10622 14660 10628 14662
rect 10320 14651 10628 14660
rect 10320 13628 10628 13637
rect 10320 13626 10326 13628
rect 10382 13626 10406 13628
rect 10462 13626 10486 13628
rect 10542 13626 10566 13628
rect 10622 13626 10628 13628
rect 10382 13574 10384 13626
rect 10564 13574 10566 13626
rect 10320 13572 10326 13574
rect 10382 13572 10406 13574
rect 10462 13572 10486 13574
rect 10542 13572 10566 13574
rect 10622 13572 10628 13574
rect 10320 13563 10628 13572
rect 10320 12540 10628 12549
rect 10320 12538 10326 12540
rect 10382 12538 10406 12540
rect 10462 12538 10486 12540
rect 10542 12538 10566 12540
rect 10622 12538 10628 12540
rect 10382 12486 10384 12538
rect 10564 12486 10566 12538
rect 10320 12484 10326 12486
rect 10382 12484 10406 12486
rect 10462 12484 10486 12486
rect 10542 12484 10566 12486
rect 10622 12484 10628 12486
rect 10320 12475 10628 12484
rect 10320 11452 10628 11461
rect 10320 11450 10326 11452
rect 10382 11450 10406 11452
rect 10462 11450 10486 11452
rect 10542 11450 10566 11452
rect 10622 11450 10628 11452
rect 10382 11398 10384 11450
rect 10564 11398 10566 11450
rect 10320 11396 10326 11398
rect 10382 11396 10406 11398
rect 10462 11396 10486 11398
rect 10542 11396 10566 11398
rect 10622 11396 10628 11398
rect 10320 11387 10628 11396
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10244 10062 10272 11290
rect 10704 10810 10732 15302
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10320 10364 10628 10373
rect 10320 10362 10326 10364
rect 10382 10362 10406 10364
rect 10462 10362 10486 10364
rect 10542 10362 10566 10364
rect 10622 10362 10628 10364
rect 10382 10310 10384 10362
rect 10564 10310 10566 10362
rect 10320 10308 10326 10310
rect 10382 10308 10406 10310
rect 10462 10308 10486 10310
rect 10542 10308 10566 10310
rect 10622 10308 10628 10310
rect 10320 10299 10628 10308
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10600 9920 10652 9926
rect 10704 9908 10732 10474
rect 10796 10266 10824 15370
rect 10980 12374 11008 16546
rect 11532 15978 11560 19200
rect 11520 15972 11572 15978
rect 11520 15914 11572 15920
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 10652 9880 10732 9908
rect 10600 9862 10652 9868
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10322 9616 10378 9625
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10152 8974 10180 9114
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10244 8906 10272 9590
rect 10322 9551 10378 9560
rect 10336 9382 10364 9551
rect 10506 9480 10562 9489
rect 10506 9415 10562 9424
rect 10520 9382 10548 9415
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10320 9276 10628 9285
rect 10320 9274 10326 9276
rect 10382 9274 10406 9276
rect 10462 9274 10486 9276
rect 10542 9274 10566 9276
rect 10622 9274 10628 9276
rect 10382 9222 10384 9274
rect 10564 9222 10566 9274
rect 10320 9220 10326 9222
rect 10382 9220 10406 9222
rect 10462 9220 10486 9222
rect 10542 9220 10566 9222
rect 10622 9220 10628 9222
rect 10320 9211 10628 9220
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 10060 3398 10088 8774
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 10244 800 10272 8842
rect 10320 8188 10628 8197
rect 10320 8186 10326 8188
rect 10382 8186 10406 8188
rect 10462 8186 10486 8188
rect 10542 8186 10566 8188
rect 10622 8186 10628 8188
rect 10382 8134 10384 8186
rect 10564 8134 10566 8186
rect 10320 8132 10326 8134
rect 10382 8132 10406 8134
rect 10462 8132 10486 8134
rect 10542 8132 10566 8134
rect 10622 8132 10628 8134
rect 10320 8123 10628 8132
rect 10320 7100 10628 7109
rect 10320 7098 10326 7100
rect 10382 7098 10406 7100
rect 10462 7098 10486 7100
rect 10542 7098 10566 7100
rect 10622 7098 10628 7100
rect 10382 7046 10384 7098
rect 10564 7046 10566 7098
rect 10320 7044 10326 7046
rect 10382 7044 10406 7046
rect 10462 7044 10486 7046
rect 10542 7044 10566 7046
rect 10622 7044 10628 7046
rect 10320 7035 10628 7044
rect 10320 6012 10628 6021
rect 10320 6010 10326 6012
rect 10382 6010 10406 6012
rect 10462 6010 10486 6012
rect 10542 6010 10566 6012
rect 10622 6010 10628 6012
rect 10382 5958 10384 6010
rect 10564 5958 10566 6010
rect 10320 5956 10326 5958
rect 10382 5956 10406 5958
rect 10462 5956 10486 5958
rect 10542 5956 10566 5958
rect 10622 5956 10628 5958
rect 10320 5947 10628 5956
rect 10320 4924 10628 4933
rect 10320 4922 10326 4924
rect 10382 4922 10406 4924
rect 10462 4922 10486 4924
rect 10542 4922 10566 4924
rect 10622 4922 10628 4924
rect 10382 4870 10384 4922
rect 10564 4870 10566 4922
rect 10320 4868 10326 4870
rect 10382 4868 10406 4870
rect 10462 4868 10486 4870
rect 10542 4868 10566 4870
rect 10622 4868 10628 4870
rect 10320 4859 10628 4868
rect 10320 3836 10628 3845
rect 10320 3834 10326 3836
rect 10382 3834 10406 3836
rect 10462 3834 10486 3836
rect 10542 3834 10566 3836
rect 10622 3834 10628 3836
rect 10382 3782 10384 3834
rect 10564 3782 10566 3834
rect 10320 3780 10326 3782
rect 10382 3780 10406 3782
rect 10462 3780 10486 3782
rect 10542 3780 10566 3782
rect 10622 3780 10628 3782
rect 10320 3771 10628 3780
rect 10704 3670 10732 9880
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10320 2748 10628 2757
rect 10320 2746 10326 2748
rect 10382 2746 10406 2748
rect 10462 2746 10486 2748
rect 10542 2746 10566 2748
rect 10622 2746 10628 2748
rect 10382 2694 10384 2746
rect 10564 2694 10566 2746
rect 10320 2692 10326 2694
rect 10382 2692 10406 2694
rect 10462 2692 10486 2694
rect 10542 2692 10566 2694
rect 10622 2692 10628 2694
rect 10320 2683 10628 2692
rect 10704 1714 10732 3130
rect 10796 3126 10824 9862
rect 10888 3466 10916 10134
rect 10980 10062 11008 10610
rect 11072 10606 11100 15370
rect 11164 11218 11192 15642
rect 11900 11898 11928 19200
rect 12268 17898 12296 19200
rect 12084 17870 12296 17898
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 10980 4010 11008 9862
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 11164 3641 11192 9862
rect 11150 3632 11206 3641
rect 11150 3567 11206 3576
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 10612 1686 10732 1714
rect 10612 800 10640 1686
rect 10980 800 11008 3470
rect 11256 2774 11284 11562
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11348 10062 11376 10746
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11716 10062 11744 10542
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11808 9382 11836 9522
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11624 3466 11652 9318
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 11256 2746 11376 2774
rect 11348 800 11376 2746
rect 11716 800 11744 4014
rect 11808 3738 11836 9318
rect 11900 9110 11928 9862
rect 11992 9450 12020 15574
rect 12084 15502 12112 17870
rect 12194 17436 12502 17445
rect 12194 17434 12200 17436
rect 12256 17434 12280 17436
rect 12336 17434 12360 17436
rect 12416 17434 12440 17436
rect 12496 17434 12502 17436
rect 12256 17382 12258 17434
rect 12438 17382 12440 17434
rect 12194 17380 12200 17382
rect 12256 17380 12280 17382
rect 12336 17380 12360 17382
rect 12416 17380 12440 17382
rect 12496 17380 12502 17382
rect 12194 17371 12502 17380
rect 12636 16574 12664 19200
rect 12544 16546 12664 16574
rect 12194 16348 12502 16357
rect 12194 16346 12200 16348
rect 12256 16346 12280 16348
rect 12336 16346 12360 16348
rect 12416 16346 12440 16348
rect 12496 16346 12502 16348
rect 12256 16294 12258 16346
rect 12438 16294 12440 16346
rect 12194 16292 12200 16294
rect 12256 16292 12280 16294
rect 12336 16292 12360 16294
rect 12416 16292 12440 16294
rect 12496 16292 12502 16294
rect 12194 16283 12502 16292
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12194 15260 12502 15269
rect 12194 15258 12200 15260
rect 12256 15258 12280 15260
rect 12336 15258 12360 15260
rect 12416 15258 12440 15260
rect 12496 15258 12502 15260
rect 12256 15206 12258 15258
rect 12438 15206 12440 15258
rect 12194 15204 12200 15206
rect 12256 15204 12280 15206
rect 12336 15204 12360 15206
rect 12416 15204 12440 15206
rect 12496 15204 12502 15206
rect 12194 15195 12502 15204
rect 12194 14172 12502 14181
rect 12194 14170 12200 14172
rect 12256 14170 12280 14172
rect 12336 14170 12360 14172
rect 12416 14170 12440 14172
rect 12496 14170 12502 14172
rect 12256 14118 12258 14170
rect 12438 14118 12440 14170
rect 12194 14116 12200 14118
rect 12256 14116 12280 14118
rect 12336 14116 12360 14118
rect 12416 14116 12440 14118
rect 12496 14116 12502 14118
rect 12194 14107 12502 14116
rect 12194 13084 12502 13093
rect 12194 13082 12200 13084
rect 12256 13082 12280 13084
rect 12336 13082 12360 13084
rect 12416 13082 12440 13084
rect 12496 13082 12502 13084
rect 12256 13030 12258 13082
rect 12438 13030 12440 13082
rect 12194 13028 12200 13030
rect 12256 13028 12280 13030
rect 12336 13028 12360 13030
rect 12416 13028 12440 13030
rect 12496 13028 12502 13030
rect 12194 13019 12502 13028
rect 12438 12744 12494 12753
rect 12438 12679 12494 12688
rect 12452 12646 12480 12679
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12194 11996 12502 12005
rect 12194 11994 12200 11996
rect 12256 11994 12280 11996
rect 12336 11994 12360 11996
rect 12416 11994 12440 11996
rect 12496 11994 12502 11996
rect 12256 11942 12258 11994
rect 12438 11942 12440 11994
rect 12194 11940 12200 11942
rect 12256 11940 12280 11942
rect 12336 11940 12360 11942
rect 12416 11940 12440 11942
rect 12496 11940 12502 11942
rect 12194 11931 12502 11940
rect 12194 10908 12502 10917
rect 12194 10906 12200 10908
rect 12256 10906 12280 10908
rect 12336 10906 12360 10908
rect 12416 10906 12440 10908
rect 12496 10906 12502 10908
rect 12256 10854 12258 10906
rect 12438 10854 12440 10906
rect 12194 10852 12200 10854
rect 12256 10852 12280 10854
rect 12336 10852 12360 10854
rect 12416 10852 12440 10854
rect 12496 10852 12502 10854
rect 12194 10843 12502 10852
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12084 10062 12112 10678
rect 12544 10538 12572 16546
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12194 9820 12502 9829
rect 12194 9818 12200 9820
rect 12256 9818 12280 9820
rect 12336 9818 12360 9820
rect 12416 9818 12440 9820
rect 12496 9818 12502 9820
rect 12256 9766 12258 9818
rect 12438 9766 12440 9818
rect 12194 9764 12200 9766
rect 12256 9764 12280 9766
rect 12336 9764 12360 9766
rect 12416 9764 12440 9766
rect 12496 9764 12502 9766
rect 12194 9755 12502 9764
rect 11980 9444 12032 9450
rect 11980 9386 12032 9392
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 12194 8732 12502 8741
rect 12194 8730 12200 8732
rect 12256 8730 12280 8732
rect 12336 8730 12360 8732
rect 12416 8730 12440 8732
rect 12496 8730 12502 8732
rect 12256 8678 12258 8730
rect 12438 8678 12440 8730
rect 12194 8676 12200 8678
rect 12256 8676 12280 8678
rect 12336 8676 12360 8678
rect 12416 8676 12440 8678
rect 12496 8676 12502 8678
rect 12194 8667 12502 8676
rect 12194 7644 12502 7653
rect 12194 7642 12200 7644
rect 12256 7642 12280 7644
rect 12336 7642 12360 7644
rect 12416 7642 12440 7644
rect 12496 7642 12502 7644
rect 12256 7590 12258 7642
rect 12438 7590 12440 7642
rect 12194 7588 12200 7590
rect 12256 7588 12280 7590
rect 12336 7588 12360 7590
rect 12416 7588 12440 7590
rect 12496 7588 12502 7590
rect 12194 7579 12502 7588
rect 12194 6556 12502 6565
rect 12194 6554 12200 6556
rect 12256 6554 12280 6556
rect 12336 6554 12360 6556
rect 12416 6554 12440 6556
rect 12496 6554 12502 6556
rect 12256 6502 12258 6554
rect 12438 6502 12440 6554
rect 12194 6500 12200 6502
rect 12256 6500 12280 6502
rect 12336 6500 12360 6502
rect 12416 6500 12440 6502
rect 12496 6500 12502 6502
rect 12194 6491 12502 6500
rect 12194 5468 12502 5477
rect 12194 5466 12200 5468
rect 12256 5466 12280 5468
rect 12336 5466 12360 5468
rect 12416 5466 12440 5468
rect 12496 5466 12502 5468
rect 12256 5414 12258 5466
rect 12438 5414 12440 5466
rect 12194 5412 12200 5414
rect 12256 5412 12280 5414
rect 12336 5412 12360 5414
rect 12416 5412 12440 5414
rect 12496 5412 12502 5414
rect 12194 5403 12502 5412
rect 12194 4380 12502 4389
rect 12194 4378 12200 4380
rect 12256 4378 12280 4380
rect 12336 4378 12360 4380
rect 12416 4378 12440 4380
rect 12496 4378 12502 4380
rect 12256 4326 12258 4378
rect 12438 4326 12440 4378
rect 12194 4324 12200 4326
rect 12256 4324 12280 4326
rect 12336 4324 12360 4326
rect 12416 4324 12440 4326
rect 12496 4324 12502 4326
rect 12194 4315 12502 4324
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 12084 800 12112 4082
rect 12544 4049 12572 9862
rect 12636 9450 12664 15506
rect 13004 15434 13032 19200
rect 12992 15428 13044 15434
rect 12992 15370 13044 15376
rect 13372 15366 13400 19200
rect 13740 17898 13768 19200
rect 14108 17898 14136 19200
rect 13648 17870 13768 17898
rect 13924 17870 14136 17898
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13648 10674 13676 17870
rect 13726 17368 13782 17377
rect 13726 17303 13782 17312
rect 13740 12986 13768 17303
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13832 10266 13860 15370
rect 13924 10810 13952 17870
rect 14068 16892 14376 16901
rect 14068 16890 14074 16892
rect 14130 16890 14154 16892
rect 14210 16890 14234 16892
rect 14290 16890 14314 16892
rect 14370 16890 14376 16892
rect 14130 16838 14132 16890
rect 14312 16838 14314 16890
rect 14068 16836 14074 16838
rect 14130 16836 14154 16838
rect 14210 16836 14234 16838
rect 14290 16836 14314 16838
rect 14370 16836 14376 16838
rect 14068 16827 14376 16836
rect 14476 16574 14504 19200
rect 14476 16546 14596 16574
rect 14068 15804 14376 15813
rect 14068 15802 14074 15804
rect 14130 15802 14154 15804
rect 14210 15802 14234 15804
rect 14290 15802 14314 15804
rect 14370 15802 14376 15804
rect 14130 15750 14132 15802
rect 14312 15750 14314 15802
rect 14068 15748 14074 15750
rect 14130 15748 14154 15750
rect 14210 15748 14234 15750
rect 14290 15748 14314 15750
rect 14370 15748 14376 15750
rect 14068 15739 14376 15748
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14068 14716 14376 14725
rect 14068 14714 14074 14716
rect 14130 14714 14154 14716
rect 14210 14714 14234 14716
rect 14290 14714 14314 14716
rect 14370 14714 14376 14716
rect 14130 14662 14132 14714
rect 14312 14662 14314 14714
rect 14068 14660 14074 14662
rect 14130 14660 14154 14662
rect 14210 14660 14234 14662
rect 14290 14660 14314 14662
rect 14370 14660 14376 14662
rect 14068 14651 14376 14660
rect 14068 13628 14376 13637
rect 14068 13626 14074 13628
rect 14130 13626 14154 13628
rect 14210 13626 14234 13628
rect 14290 13626 14314 13628
rect 14370 13626 14376 13628
rect 14130 13574 14132 13626
rect 14312 13574 14314 13626
rect 14068 13572 14074 13574
rect 14130 13572 14154 13574
rect 14210 13572 14234 13574
rect 14290 13572 14314 13574
rect 14370 13572 14376 13574
rect 14068 13563 14376 13572
rect 14068 12540 14376 12549
rect 14068 12538 14074 12540
rect 14130 12538 14154 12540
rect 14210 12538 14234 12540
rect 14290 12538 14314 12540
rect 14370 12538 14376 12540
rect 14130 12486 14132 12538
rect 14312 12486 14314 12538
rect 14068 12484 14074 12486
rect 14130 12484 14154 12486
rect 14210 12484 14234 12486
rect 14290 12484 14314 12486
rect 14370 12484 14376 12486
rect 14068 12475 14376 12484
rect 14068 11452 14376 11461
rect 14068 11450 14074 11452
rect 14130 11450 14154 11452
rect 14210 11450 14234 11452
rect 14290 11450 14314 11452
rect 14370 11450 14376 11452
rect 14130 11398 14132 11450
rect 14312 11398 14314 11450
rect 14068 11396 14074 11398
rect 14130 11396 14154 11398
rect 14210 11396 14234 11398
rect 14290 11396 14314 11398
rect 14370 11396 14376 11398
rect 14068 11387 14376 11396
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 14068 10364 14376 10373
rect 14068 10362 14074 10364
rect 14130 10362 14154 10364
rect 14210 10362 14234 10364
rect 14290 10362 14314 10364
rect 14370 10362 14376 10364
rect 14130 10310 14132 10362
rect 14312 10310 14314 10362
rect 14068 10308 14074 10310
rect 14130 10308 14154 10310
rect 14210 10308 14234 10310
rect 14290 10308 14314 10310
rect 14370 10308 14376 10310
rect 14068 10299 14376 10308
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 14476 10198 14504 15302
rect 14568 10606 14596 16546
rect 14844 15706 14872 19200
rect 15212 16574 15240 19200
rect 15120 16546 15240 16574
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14464 10192 14516 10198
rect 14464 10134 14516 10140
rect 14660 10033 14688 12582
rect 15120 10742 15148 16546
rect 15580 15434 15608 19200
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15948 15366 15976 19200
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15108 10736 15160 10742
rect 15108 10678 15160 10684
rect 14646 10024 14702 10033
rect 14646 9959 14702 9968
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 13004 9382 13032 9522
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12728 7585 12756 8298
rect 12714 7576 12770 7585
rect 12714 7511 12770 7520
rect 12530 4040 12586 4049
rect 12530 3975 12586 3984
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12194 3292 12502 3301
rect 12194 3290 12200 3292
rect 12256 3290 12280 3292
rect 12336 3290 12360 3292
rect 12416 3290 12440 3292
rect 12496 3290 12502 3292
rect 12256 3238 12258 3290
rect 12438 3238 12440 3290
rect 12194 3236 12200 3238
rect 12256 3236 12280 3238
rect 12336 3236 12360 3238
rect 12416 3236 12440 3238
rect 12496 3236 12502 3238
rect 12194 3227 12502 3236
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12452 2553 12480 2586
rect 12438 2544 12494 2553
rect 12438 2479 12494 2488
rect 12194 2204 12502 2213
rect 12194 2202 12200 2204
rect 12256 2202 12280 2204
rect 12336 2202 12360 2204
rect 12416 2202 12440 2204
rect 12496 2202 12502 2204
rect 12256 2150 12258 2202
rect 12438 2150 12440 2202
rect 12194 2148 12200 2150
rect 12256 2148 12280 2150
rect 12336 2148 12360 2150
rect 12416 2148 12440 2150
rect 12496 2148 12502 2150
rect 12194 2139 12502 2148
rect 12544 1986 12572 3538
rect 12452 1958 12572 1986
rect 12452 800 12480 1958
rect 12820 800 12848 8978
rect 13004 4146 13032 9318
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13372 4078 13400 9862
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13188 800 13216 3334
rect 13556 800 13584 9590
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 14068 9276 14376 9285
rect 14068 9274 14074 9276
rect 14130 9274 14154 9276
rect 14210 9274 14234 9276
rect 14290 9274 14314 9276
rect 14370 9274 14376 9276
rect 14130 9222 14132 9274
rect 14312 9222 14314 9274
rect 14068 9220 14074 9222
rect 14130 9220 14154 9222
rect 14210 9220 14234 9222
rect 14290 9220 14314 9222
rect 14370 9220 14376 9222
rect 14068 9211 14376 9220
rect 14068 8188 14376 8197
rect 14068 8186 14074 8188
rect 14130 8186 14154 8188
rect 14210 8186 14234 8188
rect 14290 8186 14314 8188
rect 14370 8186 14376 8188
rect 14130 8134 14132 8186
rect 14312 8134 14314 8186
rect 14068 8132 14074 8134
rect 14130 8132 14154 8134
rect 14210 8132 14234 8134
rect 14290 8132 14314 8134
rect 14370 8132 14376 8134
rect 14068 8123 14376 8132
rect 14068 7100 14376 7109
rect 14068 7098 14074 7100
rect 14130 7098 14154 7100
rect 14210 7098 14234 7100
rect 14290 7098 14314 7100
rect 14370 7098 14376 7100
rect 14130 7046 14132 7098
rect 14312 7046 14314 7098
rect 14068 7044 14074 7046
rect 14130 7044 14154 7046
rect 14210 7044 14234 7046
rect 14290 7044 14314 7046
rect 14370 7044 14376 7046
rect 14068 7035 14376 7044
rect 14068 6012 14376 6021
rect 14068 6010 14074 6012
rect 14130 6010 14154 6012
rect 14210 6010 14234 6012
rect 14290 6010 14314 6012
rect 14370 6010 14376 6012
rect 14130 5958 14132 6010
rect 14312 5958 14314 6010
rect 14068 5956 14074 5958
rect 14130 5956 14154 5958
rect 14210 5956 14234 5958
rect 14290 5956 14314 5958
rect 14370 5956 14376 5958
rect 14068 5947 14376 5956
rect 14068 4924 14376 4933
rect 14068 4922 14074 4924
rect 14130 4922 14154 4924
rect 14210 4922 14234 4924
rect 14290 4922 14314 4924
rect 14370 4922 14376 4924
rect 14130 4870 14132 4922
rect 14312 4870 14314 4922
rect 14068 4868 14074 4870
rect 14130 4868 14154 4870
rect 14210 4868 14234 4870
rect 14290 4868 14314 4870
rect 14370 4868 14376 4870
rect 14068 4859 14376 4868
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 14068 3836 14376 3845
rect 14068 3834 14074 3836
rect 14130 3834 14154 3836
rect 14210 3834 14234 3836
rect 14290 3834 14314 3836
rect 14370 3834 14376 3836
rect 14130 3782 14132 3834
rect 14312 3782 14314 3834
rect 14068 3780 14074 3782
rect 14130 3780 14154 3782
rect 14210 3780 14234 3782
rect 14290 3780 14314 3782
rect 14370 3780 14376 3782
rect 14068 3771 14376 3780
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 13832 898 13860 3402
rect 13924 1170 13952 3674
rect 14648 3664 14700 3670
rect 14648 3606 14700 3612
rect 14068 2748 14376 2757
rect 14068 2746 14074 2748
rect 14130 2746 14154 2748
rect 14210 2746 14234 2748
rect 14290 2746 14314 2748
rect 14370 2746 14376 2748
rect 14130 2694 14132 2746
rect 14312 2694 14314 2746
rect 14068 2692 14074 2694
rect 14130 2692 14154 2694
rect 14210 2692 14234 2694
rect 14290 2692 14314 2694
rect 14370 2692 14376 2694
rect 14068 2683 14376 2692
rect 13924 1142 14044 1170
rect 13832 870 13952 898
rect 13924 800 13952 870
rect 9232 734 9444 762
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14016 762 14044 1142
rect 14200 870 14320 898
rect 14200 762 14228 870
rect 14292 800 14320 870
rect 14660 800 14688 3606
rect 15028 800 15056 4014
rect 15120 2774 15148 9386
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15120 2746 15424 2774
rect 15396 800 15424 2746
rect 15764 800 15792 4082
rect 14016 734 14228 762
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
<< via2 >>
rect 1766 14864 1822 14920
rect 2830 16890 2886 16892
rect 2910 16890 2966 16892
rect 2990 16890 3046 16892
rect 3070 16890 3126 16892
rect 2830 16838 2876 16890
rect 2876 16838 2886 16890
rect 2910 16838 2940 16890
rect 2940 16838 2952 16890
rect 2952 16838 2966 16890
rect 2990 16838 3004 16890
rect 3004 16838 3016 16890
rect 3016 16838 3046 16890
rect 3070 16838 3080 16890
rect 3080 16838 3126 16890
rect 2830 16836 2886 16838
rect 2910 16836 2966 16838
rect 2990 16836 3046 16838
rect 3070 16836 3126 16838
rect 2830 15802 2886 15804
rect 2910 15802 2966 15804
rect 2990 15802 3046 15804
rect 3070 15802 3126 15804
rect 2830 15750 2876 15802
rect 2876 15750 2886 15802
rect 2910 15750 2940 15802
rect 2940 15750 2952 15802
rect 2952 15750 2966 15802
rect 2990 15750 3004 15802
rect 3004 15750 3016 15802
rect 3016 15750 3046 15802
rect 3070 15750 3080 15802
rect 3080 15750 3126 15802
rect 2830 15748 2886 15750
rect 2910 15748 2966 15750
rect 2990 15748 3046 15750
rect 3070 15748 3126 15750
rect 4066 18128 4122 18184
rect 2830 14714 2886 14716
rect 2910 14714 2966 14716
rect 2990 14714 3046 14716
rect 3070 14714 3126 14716
rect 2830 14662 2876 14714
rect 2876 14662 2886 14714
rect 2910 14662 2940 14714
rect 2940 14662 2952 14714
rect 2952 14662 2966 14714
rect 2990 14662 3004 14714
rect 3004 14662 3016 14714
rect 3016 14662 3046 14714
rect 3070 14662 3080 14714
rect 3080 14662 3126 14714
rect 2830 14660 2886 14662
rect 2910 14660 2966 14662
rect 2990 14660 3046 14662
rect 3070 14660 3126 14662
rect 2830 13626 2886 13628
rect 2910 13626 2966 13628
rect 2990 13626 3046 13628
rect 3070 13626 3126 13628
rect 2830 13574 2876 13626
rect 2876 13574 2886 13626
rect 2910 13574 2940 13626
rect 2940 13574 2952 13626
rect 2952 13574 2966 13626
rect 2990 13574 3004 13626
rect 3004 13574 3016 13626
rect 3016 13574 3046 13626
rect 3070 13574 3080 13626
rect 3080 13574 3126 13626
rect 2830 13572 2886 13574
rect 2910 13572 2966 13574
rect 2990 13572 3046 13574
rect 3070 13572 3126 13574
rect 2830 12538 2886 12540
rect 2910 12538 2966 12540
rect 2990 12538 3046 12540
rect 3070 12538 3126 12540
rect 2830 12486 2876 12538
rect 2876 12486 2886 12538
rect 2910 12486 2940 12538
rect 2940 12486 2952 12538
rect 2952 12486 2966 12538
rect 2990 12486 3004 12538
rect 3004 12486 3016 12538
rect 3016 12486 3046 12538
rect 3070 12486 3080 12538
rect 3080 12486 3126 12538
rect 2830 12484 2886 12486
rect 2910 12484 2966 12486
rect 2990 12484 3046 12486
rect 3070 12484 3126 12486
rect 2830 11450 2886 11452
rect 2910 11450 2966 11452
rect 2990 11450 3046 11452
rect 3070 11450 3126 11452
rect 2830 11398 2876 11450
rect 2876 11398 2886 11450
rect 2910 11398 2940 11450
rect 2940 11398 2952 11450
rect 2952 11398 2966 11450
rect 2990 11398 3004 11450
rect 3004 11398 3016 11450
rect 3016 11398 3046 11450
rect 3070 11398 3080 11450
rect 3080 11398 3126 11450
rect 2830 11396 2886 11398
rect 2910 11396 2966 11398
rect 2990 11396 3046 11398
rect 3070 11396 3126 11398
rect 4158 11600 4214 11656
rect 2830 10362 2886 10364
rect 2910 10362 2966 10364
rect 2990 10362 3046 10364
rect 3070 10362 3126 10364
rect 2830 10310 2876 10362
rect 2876 10310 2886 10362
rect 2910 10310 2940 10362
rect 2940 10310 2952 10362
rect 2952 10310 2966 10362
rect 2990 10310 3004 10362
rect 3004 10310 3016 10362
rect 3016 10310 3046 10362
rect 3070 10310 3080 10362
rect 3080 10310 3126 10362
rect 2830 10308 2886 10310
rect 2910 10308 2966 10310
rect 2990 10308 3046 10310
rect 3070 10308 3126 10310
rect 2830 9274 2886 9276
rect 2910 9274 2966 9276
rect 2990 9274 3046 9276
rect 3070 9274 3126 9276
rect 2830 9222 2876 9274
rect 2876 9222 2886 9274
rect 2910 9222 2940 9274
rect 2940 9222 2952 9274
rect 2952 9222 2966 9274
rect 2990 9222 3004 9274
rect 3004 9222 3016 9274
rect 3016 9222 3046 9274
rect 3070 9222 3080 9274
rect 3080 9222 3126 9274
rect 2830 9220 2886 9222
rect 2910 9220 2966 9222
rect 2990 9220 3046 9222
rect 3070 9220 3126 9222
rect 2830 8186 2886 8188
rect 2910 8186 2966 8188
rect 2990 8186 3046 8188
rect 3070 8186 3126 8188
rect 2830 8134 2876 8186
rect 2876 8134 2886 8186
rect 2910 8134 2940 8186
rect 2940 8134 2952 8186
rect 2952 8134 2966 8186
rect 2990 8134 3004 8186
rect 3004 8134 3016 8186
rect 3016 8134 3046 8186
rect 3070 8134 3080 8186
rect 3080 8134 3126 8186
rect 2830 8132 2886 8134
rect 2910 8132 2966 8134
rect 2990 8132 3046 8134
rect 3070 8132 3126 8134
rect 2830 7098 2886 7100
rect 2910 7098 2966 7100
rect 2990 7098 3046 7100
rect 3070 7098 3126 7100
rect 2830 7046 2876 7098
rect 2876 7046 2886 7098
rect 2910 7046 2940 7098
rect 2940 7046 2952 7098
rect 2952 7046 2966 7098
rect 2990 7046 3004 7098
rect 3004 7046 3016 7098
rect 3016 7046 3046 7098
rect 3070 7046 3080 7098
rect 3080 7046 3126 7098
rect 2830 7044 2886 7046
rect 2910 7044 2966 7046
rect 2990 7044 3046 7046
rect 3070 7044 3126 7046
rect 2830 6010 2886 6012
rect 2910 6010 2966 6012
rect 2990 6010 3046 6012
rect 3070 6010 3126 6012
rect 2830 5958 2876 6010
rect 2876 5958 2886 6010
rect 2910 5958 2940 6010
rect 2940 5958 2952 6010
rect 2952 5958 2966 6010
rect 2990 5958 3004 6010
rect 3004 5958 3016 6010
rect 3016 5958 3046 6010
rect 3070 5958 3080 6010
rect 3080 5958 3126 6010
rect 2830 5956 2886 5958
rect 2910 5956 2966 5958
rect 2990 5956 3046 5958
rect 3070 5956 3126 5958
rect 2830 4922 2886 4924
rect 2910 4922 2966 4924
rect 2990 4922 3046 4924
rect 3070 4922 3126 4924
rect 2830 4870 2876 4922
rect 2876 4870 2886 4922
rect 2910 4870 2940 4922
rect 2940 4870 2952 4922
rect 2952 4870 2966 4922
rect 2990 4870 3004 4922
rect 3004 4870 3016 4922
rect 3016 4870 3046 4922
rect 3070 4870 3080 4922
rect 3080 4870 3126 4922
rect 2830 4868 2886 4870
rect 2910 4868 2966 4870
rect 2990 4868 3046 4870
rect 3070 4868 3126 4870
rect 2830 3834 2886 3836
rect 2910 3834 2966 3836
rect 2990 3834 3046 3836
rect 3070 3834 3126 3836
rect 2830 3782 2876 3834
rect 2876 3782 2886 3834
rect 2910 3782 2940 3834
rect 2940 3782 2952 3834
rect 2952 3782 2966 3834
rect 2990 3782 3004 3834
rect 3004 3782 3016 3834
rect 3016 3782 3046 3834
rect 3070 3782 3080 3834
rect 3080 3782 3126 3834
rect 2830 3780 2886 3782
rect 2910 3780 2966 3782
rect 2990 3780 3046 3782
rect 3070 3780 3126 3782
rect 2830 2746 2886 2748
rect 2910 2746 2966 2748
rect 2990 2746 3046 2748
rect 3070 2746 3126 2748
rect 2830 2694 2876 2746
rect 2876 2694 2886 2746
rect 2910 2694 2940 2746
rect 2940 2694 2952 2746
rect 2952 2694 2966 2746
rect 2990 2694 3004 2746
rect 3004 2694 3016 2746
rect 3016 2694 3046 2746
rect 3070 2694 3080 2746
rect 3080 2694 3126 2746
rect 2830 2692 2886 2694
rect 2910 2692 2966 2694
rect 2990 2692 3046 2694
rect 3070 2692 3126 2694
rect 3238 8336 3294 8392
rect 3238 5072 3294 5128
rect 3146 1808 3202 1864
rect 4704 17434 4760 17436
rect 4784 17434 4840 17436
rect 4864 17434 4920 17436
rect 4944 17434 5000 17436
rect 4704 17382 4750 17434
rect 4750 17382 4760 17434
rect 4784 17382 4814 17434
rect 4814 17382 4826 17434
rect 4826 17382 4840 17434
rect 4864 17382 4878 17434
rect 4878 17382 4890 17434
rect 4890 17382 4920 17434
rect 4944 17382 4954 17434
rect 4954 17382 5000 17434
rect 4704 17380 4760 17382
rect 4784 17380 4840 17382
rect 4864 17380 4920 17382
rect 4944 17380 5000 17382
rect 4704 16346 4760 16348
rect 4784 16346 4840 16348
rect 4864 16346 4920 16348
rect 4944 16346 5000 16348
rect 4704 16294 4750 16346
rect 4750 16294 4760 16346
rect 4784 16294 4814 16346
rect 4814 16294 4826 16346
rect 4826 16294 4840 16346
rect 4864 16294 4878 16346
rect 4878 16294 4890 16346
rect 4890 16294 4920 16346
rect 4944 16294 4954 16346
rect 4954 16294 5000 16346
rect 4704 16292 4760 16294
rect 4784 16292 4840 16294
rect 4864 16292 4920 16294
rect 4944 16292 5000 16294
rect 4704 15258 4760 15260
rect 4784 15258 4840 15260
rect 4864 15258 4920 15260
rect 4944 15258 5000 15260
rect 4704 15206 4750 15258
rect 4750 15206 4760 15258
rect 4784 15206 4814 15258
rect 4814 15206 4826 15258
rect 4826 15206 4840 15258
rect 4864 15206 4878 15258
rect 4878 15206 4890 15258
rect 4890 15206 4920 15258
rect 4944 15206 4954 15258
rect 4954 15206 5000 15258
rect 4704 15204 4760 15206
rect 4784 15204 4840 15206
rect 4864 15204 4920 15206
rect 4944 15204 5000 15206
rect 4704 14170 4760 14172
rect 4784 14170 4840 14172
rect 4864 14170 4920 14172
rect 4944 14170 5000 14172
rect 4704 14118 4750 14170
rect 4750 14118 4760 14170
rect 4784 14118 4814 14170
rect 4814 14118 4826 14170
rect 4826 14118 4840 14170
rect 4864 14118 4878 14170
rect 4878 14118 4890 14170
rect 4890 14118 4920 14170
rect 4944 14118 4954 14170
rect 4954 14118 5000 14170
rect 4704 14116 4760 14118
rect 4784 14116 4840 14118
rect 4864 14116 4920 14118
rect 4944 14116 5000 14118
rect 4704 13082 4760 13084
rect 4784 13082 4840 13084
rect 4864 13082 4920 13084
rect 4944 13082 5000 13084
rect 4704 13030 4750 13082
rect 4750 13030 4760 13082
rect 4784 13030 4814 13082
rect 4814 13030 4826 13082
rect 4826 13030 4840 13082
rect 4864 13030 4878 13082
rect 4878 13030 4890 13082
rect 4890 13030 4920 13082
rect 4944 13030 4954 13082
rect 4954 13030 5000 13082
rect 4704 13028 4760 13030
rect 4784 13028 4840 13030
rect 4864 13028 4920 13030
rect 4944 13028 5000 13030
rect 4704 11994 4760 11996
rect 4784 11994 4840 11996
rect 4864 11994 4920 11996
rect 4944 11994 5000 11996
rect 4704 11942 4750 11994
rect 4750 11942 4760 11994
rect 4784 11942 4814 11994
rect 4814 11942 4826 11994
rect 4826 11942 4840 11994
rect 4864 11942 4878 11994
rect 4878 11942 4890 11994
rect 4890 11942 4920 11994
rect 4944 11942 4954 11994
rect 4954 11942 5000 11994
rect 4704 11940 4760 11942
rect 4784 11940 4840 11942
rect 4864 11940 4920 11942
rect 4944 11940 5000 11942
rect 5538 11328 5594 11384
rect 4704 10906 4760 10908
rect 4784 10906 4840 10908
rect 4864 10906 4920 10908
rect 4944 10906 5000 10908
rect 4704 10854 4750 10906
rect 4750 10854 4760 10906
rect 4784 10854 4814 10906
rect 4814 10854 4826 10906
rect 4826 10854 4840 10906
rect 4864 10854 4878 10906
rect 4878 10854 4890 10906
rect 4890 10854 4920 10906
rect 4944 10854 4954 10906
rect 4954 10854 5000 10906
rect 4704 10852 4760 10854
rect 4784 10852 4840 10854
rect 4864 10852 4920 10854
rect 4944 10852 5000 10854
rect 4704 9818 4760 9820
rect 4784 9818 4840 9820
rect 4864 9818 4920 9820
rect 4944 9818 5000 9820
rect 4704 9766 4750 9818
rect 4750 9766 4760 9818
rect 4784 9766 4814 9818
rect 4814 9766 4826 9818
rect 4826 9766 4840 9818
rect 4864 9766 4878 9818
rect 4878 9766 4890 9818
rect 4890 9766 4920 9818
rect 4944 9766 4954 9818
rect 4954 9766 5000 9818
rect 4704 9764 4760 9766
rect 4784 9764 4840 9766
rect 4864 9764 4920 9766
rect 4944 9764 5000 9766
rect 4704 8730 4760 8732
rect 4784 8730 4840 8732
rect 4864 8730 4920 8732
rect 4944 8730 5000 8732
rect 4704 8678 4750 8730
rect 4750 8678 4760 8730
rect 4784 8678 4814 8730
rect 4814 8678 4826 8730
rect 4826 8678 4840 8730
rect 4864 8678 4878 8730
rect 4878 8678 4890 8730
rect 4890 8678 4920 8730
rect 4944 8678 4954 8730
rect 4954 8678 5000 8730
rect 4704 8676 4760 8678
rect 4784 8676 4840 8678
rect 4864 8676 4920 8678
rect 4944 8676 5000 8678
rect 5722 11328 5778 11384
rect 5630 9560 5686 9616
rect 4704 7642 4760 7644
rect 4784 7642 4840 7644
rect 4864 7642 4920 7644
rect 4944 7642 5000 7644
rect 4704 7590 4750 7642
rect 4750 7590 4760 7642
rect 4784 7590 4814 7642
rect 4814 7590 4826 7642
rect 4826 7590 4840 7642
rect 4864 7590 4878 7642
rect 4878 7590 4890 7642
rect 4890 7590 4920 7642
rect 4944 7590 4954 7642
rect 4954 7590 5000 7642
rect 4704 7588 4760 7590
rect 4784 7588 4840 7590
rect 4864 7588 4920 7590
rect 4944 7588 5000 7590
rect 4704 6554 4760 6556
rect 4784 6554 4840 6556
rect 4864 6554 4920 6556
rect 4944 6554 5000 6556
rect 4704 6502 4750 6554
rect 4750 6502 4760 6554
rect 4784 6502 4814 6554
rect 4814 6502 4826 6554
rect 4826 6502 4840 6554
rect 4864 6502 4878 6554
rect 4878 6502 4890 6554
rect 4890 6502 4920 6554
rect 4944 6502 4954 6554
rect 4954 6502 5000 6554
rect 4704 6500 4760 6502
rect 4784 6500 4840 6502
rect 4864 6500 4920 6502
rect 4944 6500 5000 6502
rect 4704 5466 4760 5468
rect 4784 5466 4840 5468
rect 4864 5466 4920 5468
rect 4944 5466 5000 5468
rect 4704 5414 4750 5466
rect 4750 5414 4760 5466
rect 4784 5414 4814 5466
rect 4814 5414 4826 5466
rect 4826 5414 4840 5466
rect 4864 5414 4878 5466
rect 4878 5414 4890 5466
rect 4890 5414 4920 5466
rect 4944 5414 4954 5466
rect 4954 5414 5000 5466
rect 4704 5412 4760 5414
rect 4784 5412 4840 5414
rect 4864 5412 4920 5414
rect 4944 5412 5000 5414
rect 4704 4378 4760 4380
rect 4784 4378 4840 4380
rect 4864 4378 4920 4380
rect 4944 4378 5000 4380
rect 4704 4326 4750 4378
rect 4750 4326 4760 4378
rect 4784 4326 4814 4378
rect 4814 4326 4826 4378
rect 4826 4326 4840 4378
rect 4864 4326 4878 4378
rect 4878 4326 4890 4378
rect 4890 4326 4920 4378
rect 4944 4326 4954 4378
rect 4954 4326 5000 4378
rect 4704 4324 4760 4326
rect 4784 4324 4840 4326
rect 4864 4324 4920 4326
rect 4944 4324 5000 4326
rect 4704 3290 4760 3292
rect 4784 3290 4840 3292
rect 4864 3290 4920 3292
rect 4944 3290 5000 3292
rect 4704 3238 4750 3290
rect 4750 3238 4760 3290
rect 4784 3238 4814 3290
rect 4814 3238 4826 3290
rect 4826 3238 4840 3290
rect 4864 3238 4878 3290
rect 4878 3238 4890 3290
rect 4890 3238 4920 3290
rect 4944 3238 4954 3290
rect 4954 3238 5000 3290
rect 4704 3236 4760 3238
rect 4784 3236 4840 3238
rect 4864 3236 4920 3238
rect 4944 3236 5000 3238
rect 4704 2202 4760 2204
rect 4784 2202 4840 2204
rect 4864 2202 4920 2204
rect 4944 2202 5000 2204
rect 4704 2150 4750 2202
rect 4750 2150 4760 2202
rect 4784 2150 4814 2202
rect 4814 2150 4826 2202
rect 4826 2150 4840 2202
rect 4864 2150 4878 2202
rect 4878 2150 4890 2202
rect 4890 2150 4920 2202
rect 4944 2150 4954 2202
rect 4954 2150 5000 2202
rect 4704 2148 4760 2150
rect 4784 2148 4840 2150
rect 4864 2148 4920 2150
rect 4944 2148 5000 2150
rect 6578 16890 6634 16892
rect 6658 16890 6714 16892
rect 6738 16890 6794 16892
rect 6818 16890 6874 16892
rect 6578 16838 6624 16890
rect 6624 16838 6634 16890
rect 6658 16838 6688 16890
rect 6688 16838 6700 16890
rect 6700 16838 6714 16890
rect 6738 16838 6752 16890
rect 6752 16838 6764 16890
rect 6764 16838 6794 16890
rect 6818 16838 6828 16890
rect 6828 16838 6874 16890
rect 6578 16836 6634 16838
rect 6658 16836 6714 16838
rect 6738 16836 6794 16838
rect 6818 16836 6874 16838
rect 5998 9424 6054 9480
rect 5998 8880 6054 8936
rect 6182 9016 6238 9072
rect 6578 15802 6634 15804
rect 6658 15802 6714 15804
rect 6738 15802 6794 15804
rect 6818 15802 6874 15804
rect 6578 15750 6624 15802
rect 6624 15750 6634 15802
rect 6658 15750 6688 15802
rect 6688 15750 6700 15802
rect 6700 15750 6714 15802
rect 6738 15750 6752 15802
rect 6752 15750 6764 15802
rect 6764 15750 6794 15802
rect 6818 15750 6828 15802
rect 6828 15750 6874 15802
rect 6578 15748 6634 15750
rect 6658 15748 6714 15750
rect 6738 15748 6794 15750
rect 6818 15748 6874 15750
rect 6578 14714 6634 14716
rect 6658 14714 6714 14716
rect 6738 14714 6794 14716
rect 6818 14714 6874 14716
rect 6578 14662 6624 14714
rect 6624 14662 6634 14714
rect 6658 14662 6688 14714
rect 6688 14662 6700 14714
rect 6700 14662 6714 14714
rect 6738 14662 6752 14714
rect 6752 14662 6764 14714
rect 6764 14662 6794 14714
rect 6818 14662 6828 14714
rect 6828 14662 6874 14714
rect 6578 14660 6634 14662
rect 6658 14660 6714 14662
rect 6738 14660 6794 14662
rect 6818 14660 6874 14662
rect 6578 13626 6634 13628
rect 6658 13626 6714 13628
rect 6738 13626 6794 13628
rect 6818 13626 6874 13628
rect 6578 13574 6624 13626
rect 6624 13574 6634 13626
rect 6658 13574 6688 13626
rect 6688 13574 6700 13626
rect 6700 13574 6714 13626
rect 6738 13574 6752 13626
rect 6752 13574 6764 13626
rect 6764 13574 6794 13626
rect 6818 13574 6828 13626
rect 6828 13574 6874 13626
rect 6578 13572 6634 13574
rect 6658 13572 6714 13574
rect 6738 13572 6794 13574
rect 6818 13572 6874 13574
rect 6578 12538 6634 12540
rect 6658 12538 6714 12540
rect 6738 12538 6794 12540
rect 6818 12538 6874 12540
rect 6578 12486 6624 12538
rect 6624 12486 6634 12538
rect 6658 12486 6688 12538
rect 6688 12486 6700 12538
rect 6700 12486 6714 12538
rect 6738 12486 6752 12538
rect 6752 12486 6764 12538
rect 6764 12486 6794 12538
rect 6818 12486 6828 12538
rect 6828 12486 6874 12538
rect 6578 12484 6634 12486
rect 6658 12484 6714 12486
rect 6738 12484 6794 12486
rect 6818 12484 6874 12486
rect 6578 11450 6634 11452
rect 6658 11450 6714 11452
rect 6738 11450 6794 11452
rect 6818 11450 6874 11452
rect 6578 11398 6624 11450
rect 6624 11398 6634 11450
rect 6658 11398 6688 11450
rect 6688 11398 6700 11450
rect 6700 11398 6714 11450
rect 6738 11398 6752 11450
rect 6752 11398 6764 11450
rect 6764 11398 6794 11450
rect 6818 11398 6828 11450
rect 6828 11398 6874 11450
rect 6578 11396 6634 11398
rect 6658 11396 6714 11398
rect 6738 11396 6794 11398
rect 6818 11396 6874 11398
rect 6578 10362 6634 10364
rect 6658 10362 6714 10364
rect 6738 10362 6794 10364
rect 6818 10362 6874 10364
rect 6578 10310 6624 10362
rect 6624 10310 6634 10362
rect 6658 10310 6688 10362
rect 6688 10310 6700 10362
rect 6700 10310 6714 10362
rect 6738 10310 6752 10362
rect 6752 10310 6764 10362
rect 6764 10310 6794 10362
rect 6818 10310 6828 10362
rect 6828 10310 6874 10362
rect 6578 10308 6634 10310
rect 6658 10308 6714 10310
rect 6738 10308 6794 10310
rect 6818 10308 6874 10310
rect 6826 9988 6882 10024
rect 6826 9968 6828 9988
rect 6828 9968 6880 9988
rect 6880 9968 6882 9988
rect 6578 9274 6634 9276
rect 6658 9274 6714 9276
rect 6738 9274 6794 9276
rect 6818 9274 6874 9276
rect 6578 9222 6624 9274
rect 6624 9222 6634 9274
rect 6658 9222 6688 9274
rect 6688 9222 6700 9274
rect 6700 9222 6714 9274
rect 6738 9222 6752 9274
rect 6752 9222 6764 9274
rect 6764 9222 6794 9274
rect 6818 9222 6828 9274
rect 6828 9222 6874 9274
rect 6578 9220 6634 9222
rect 6658 9220 6714 9222
rect 6738 9220 6794 9222
rect 6818 9220 6874 9222
rect 6578 8186 6634 8188
rect 6658 8186 6714 8188
rect 6738 8186 6794 8188
rect 6818 8186 6874 8188
rect 6578 8134 6624 8186
rect 6624 8134 6634 8186
rect 6658 8134 6688 8186
rect 6688 8134 6700 8186
rect 6700 8134 6714 8186
rect 6738 8134 6752 8186
rect 6752 8134 6764 8186
rect 6764 8134 6794 8186
rect 6818 8134 6828 8186
rect 6828 8134 6874 8186
rect 6578 8132 6634 8134
rect 6658 8132 6714 8134
rect 6738 8132 6794 8134
rect 6818 8132 6874 8134
rect 6578 7098 6634 7100
rect 6658 7098 6714 7100
rect 6738 7098 6794 7100
rect 6818 7098 6874 7100
rect 6578 7046 6624 7098
rect 6624 7046 6634 7098
rect 6658 7046 6688 7098
rect 6688 7046 6700 7098
rect 6700 7046 6714 7098
rect 6738 7046 6752 7098
rect 6752 7046 6764 7098
rect 6764 7046 6794 7098
rect 6818 7046 6828 7098
rect 6828 7046 6874 7098
rect 6578 7044 6634 7046
rect 6658 7044 6714 7046
rect 6738 7044 6794 7046
rect 6818 7044 6874 7046
rect 6578 6010 6634 6012
rect 6658 6010 6714 6012
rect 6738 6010 6794 6012
rect 6818 6010 6874 6012
rect 6578 5958 6624 6010
rect 6624 5958 6634 6010
rect 6658 5958 6688 6010
rect 6688 5958 6700 6010
rect 6700 5958 6714 6010
rect 6738 5958 6752 6010
rect 6752 5958 6764 6010
rect 6764 5958 6794 6010
rect 6818 5958 6828 6010
rect 6828 5958 6874 6010
rect 6578 5956 6634 5958
rect 6658 5956 6714 5958
rect 6738 5956 6794 5958
rect 6818 5956 6874 5958
rect 6578 4922 6634 4924
rect 6658 4922 6714 4924
rect 6738 4922 6794 4924
rect 6818 4922 6874 4924
rect 6578 4870 6624 4922
rect 6624 4870 6634 4922
rect 6658 4870 6688 4922
rect 6688 4870 6700 4922
rect 6700 4870 6714 4922
rect 6738 4870 6752 4922
rect 6752 4870 6764 4922
rect 6764 4870 6794 4922
rect 6818 4870 6828 4922
rect 6828 4870 6874 4922
rect 6578 4868 6634 4870
rect 6658 4868 6714 4870
rect 6738 4868 6794 4870
rect 6818 4868 6874 4870
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8498 17434
rect 8498 17382 8508 17434
rect 8532 17382 8562 17434
rect 8562 17382 8574 17434
rect 8574 17382 8588 17434
rect 8612 17382 8626 17434
rect 8626 17382 8638 17434
rect 8638 17382 8668 17434
rect 8692 17382 8702 17434
rect 8702 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8498 16346
rect 8498 16294 8508 16346
rect 8532 16294 8562 16346
rect 8562 16294 8574 16346
rect 8574 16294 8588 16346
rect 8612 16294 8626 16346
rect 8626 16294 8638 16346
rect 8638 16294 8668 16346
rect 8692 16294 8702 16346
rect 8702 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8498 15258
rect 8498 15206 8508 15258
rect 8532 15206 8562 15258
rect 8562 15206 8574 15258
rect 8574 15206 8588 15258
rect 8612 15206 8626 15258
rect 8626 15206 8638 15258
rect 8638 15206 8668 15258
rect 8692 15206 8702 15258
rect 8702 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8498 14170
rect 8498 14118 8508 14170
rect 8532 14118 8562 14170
rect 8562 14118 8574 14170
rect 8574 14118 8588 14170
rect 8612 14118 8626 14170
rect 8626 14118 8638 14170
rect 8638 14118 8668 14170
rect 8692 14118 8702 14170
rect 8702 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8498 13082
rect 8498 13030 8508 13082
rect 8532 13030 8562 13082
rect 8562 13030 8574 13082
rect 8574 13030 8588 13082
rect 8612 13030 8626 13082
rect 8626 13030 8638 13082
rect 8638 13030 8668 13082
rect 8692 13030 8702 13082
rect 8702 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 6578 3834 6634 3836
rect 6658 3834 6714 3836
rect 6738 3834 6794 3836
rect 6818 3834 6874 3836
rect 6578 3782 6624 3834
rect 6624 3782 6634 3834
rect 6658 3782 6688 3834
rect 6688 3782 6700 3834
rect 6700 3782 6714 3834
rect 6738 3782 6752 3834
rect 6752 3782 6764 3834
rect 6764 3782 6794 3834
rect 6818 3782 6828 3834
rect 6828 3782 6874 3834
rect 6578 3780 6634 3782
rect 6658 3780 6714 3782
rect 6738 3780 6794 3782
rect 6818 3780 6874 3782
rect 6458 3576 6514 3632
rect 6578 2746 6634 2748
rect 6658 2746 6714 2748
rect 6738 2746 6794 2748
rect 6818 2746 6874 2748
rect 6578 2694 6624 2746
rect 6624 2694 6634 2746
rect 6658 2694 6688 2746
rect 6688 2694 6700 2746
rect 6700 2694 6714 2746
rect 6738 2694 6752 2746
rect 6752 2694 6764 2746
rect 6764 2694 6794 2746
rect 6818 2694 6828 2746
rect 6828 2694 6874 2746
rect 6578 2692 6634 2694
rect 6658 2692 6714 2694
rect 6738 2692 6794 2694
rect 6818 2692 6874 2694
rect 7746 10104 7802 10160
rect 7746 9288 7802 9344
rect 8022 3984 8078 4040
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8498 11994
rect 8498 11942 8508 11994
rect 8532 11942 8562 11994
rect 8562 11942 8574 11994
rect 8574 11942 8588 11994
rect 8612 11942 8626 11994
rect 8626 11942 8638 11994
rect 8638 11942 8668 11994
rect 8692 11942 8702 11994
rect 8702 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 9034 11192 9090 11248
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8498 10906
rect 8498 10854 8508 10906
rect 8532 10854 8562 10906
rect 8562 10854 8574 10906
rect 8574 10854 8588 10906
rect 8612 10854 8626 10906
rect 8626 10854 8638 10906
rect 8638 10854 8668 10906
rect 8692 10854 8702 10906
rect 8702 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 9034 10104 9090 10160
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8498 9818
rect 8498 9766 8508 9818
rect 8532 9766 8562 9818
rect 8562 9766 8574 9818
rect 8574 9766 8588 9818
rect 8612 9766 8626 9818
rect 8626 9766 8638 9818
rect 8638 9766 8668 9818
rect 8692 9766 8702 9818
rect 8702 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8850 9696 8906 9752
rect 8206 9152 8262 9208
rect 8482 9288 8538 9344
rect 8666 9152 8722 9208
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8498 8730
rect 8498 8678 8508 8730
rect 8532 8678 8562 8730
rect 8562 8678 8574 8730
rect 8574 8678 8588 8730
rect 8612 8678 8626 8730
rect 8626 8678 8638 8730
rect 8638 8678 8668 8730
rect 8692 8678 8702 8730
rect 8702 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 9034 9288 9090 9344
rect 9034 8880 9090 8936
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8498 7642
rect 8498 7590 8508 7642
rect 8532 7590 8562 7642
rect 8562 7590 8574 7642
rect 8574 7590 8588 7642
rect 8612 7590 8626 7642
rect 8626 7590 8638 7642
rect 8638 7590 8668 7642
rect 8692 7590 8702 7642
rect 8702 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8498 6554
rect 8498 6502 8508 6554
rect 8532 6502 8562 6554
rect 8562 6502 8574 6554
rect 8574 6502 8588 6554
rect 8612 6502 8626 6554
rect 8626 6502 8638 6554
rect 8638 6502 8668 6554
rect 8692 6502 8702 6554
rect 8702 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8498 5466
rect 8498 5414 8508 5466
rect 8532 5414 8562 5466
rect 8562 5414 8574 5466
rect 8574 5414 8588 5466
rect 8612 5414 8626 5466
rect 8626 5414 8638 5466
rect 8638 5414 8668 5466
rect 8692 5414 8702 5466
rect 8702 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8498 4378
rect 8498 4326 8508 4378
rect 8532 4326 8562 4378
rect 8562 4326 8574 4378
rect 8574 4326 8588 4378
rect 8612 4326 8626 4378
rect 8626 4326 8638 4378
rect 8638 4326 8668 4378
rect 8692 4326 8702 4378
rect 8702 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8498 3290
rect 8498 3238 8508 3290
rect 8532 3238 8562 3290
rect 8562 3238 8574 3290
rect 8574 3238 8588 3290
rect 8612 3238 8626 3290
rect 8626 3238 8638 3290
rect 8638 3238 8668 3290
rect 8692 3238 8702 3290
rect 8702 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8498 2202
rect 8498 2150 8508 2202
rect 8532 2150 8562 2202
rect 8562 2150 8574 2202
rect 8574 2150 8588 2202
rect 8612 2150 8626 2202
rect 8626 2150 8638 2202
rect 8638 2150 8668 2202
rect 8692 2150 8702 2202
rect 8702 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 9402 9288 9458 9344
rect 9770 9424 9826 9480
rect 10326 16890 10382 16892
rect 10406 16890 10462 16892
rect 10486 16890 10542 16892
rect 10566 16890 10622 16892
rect 10326 16838 10372 16890
rect 10372 16838 10382 16890
rect 10406 16838 10436 16890
rect 10436 16838 10448 16890
rect 10448 16838 10462 16890
rect 10486 16838 10500 16890
rect 10500 16838 10512 16890
rect 10512 16838 10542 16890
rect 10566 16838 10576 16890
rect 10576 16838 10622 16890
rect 10326 16836 10382 16838
rect 10406 16836 10462 16838
rect 10486 16836 10542 16838
rect 10566 16836 10622 16838
rect 10326 15802 10382 15804
rect 10406 15802 10462 15804
rect 10486 15802 10542 15804
rect 10566 15802 10622 15804
rect 10326 15750 10372 15802
rect 10372 15750 10382 15802
rect 10406 15750 10436 15802
rect 10436 15750 10448 15802
rect 10448 15750 10462 15802
rect 10486 15750 10500 15802
rect 10500 15750 10512 15802
rect 10512 15750 10542 15802
rect 10566 15750 10576 15802
rect 10576 15750 10622 15802
rect 10326 15748 10382 15750
rect 10406 15748 10462 15750
rect 10486 15748 10542 15750
rect 10566 15748 10622 15750
rect 10326 14714 10382 14716
rect 10406 14714 10462 14716
rect 10486 14714 10542 14716
rect 10566 14714 10622 14716
rect 10326 14662 10372 14714
rect 10372 14662 10382 14714
rect 10406 14662 10436 14714
rect 10436 14662 10448 14714
rect 10448 14662 10462 14714
rect 10486 14662 10500 14714
rect 10500 14662 10512 14714
rect 10512 14662 10542 14714
rect 10566 14662 10576 14714
rect 10576 14662 10622 14714
rect 10326 14660 10382 14662
rect 10406 14660 10462 14662
rect 10486 14660 10542 14662
rect 10566 14660 10622 14662
rect 10326 13626 10382 13628
rect 10406 13626 10462 13628
rect 10486 13626 10542 13628
rect 10566 13626 10622 13628
rect 10326 13574 10372 13626
rect 10372 13574 10382 13626
rect 10406 13574 10436 13626
rect 10436 13574 10448 13626
rect 10448 13574 10462 13626
rect 10486 13574 10500 13626
rect 10500 13574 10512 13626
rect 10512 13574 10542 13626
rect 10566 13574 10576 13626
rect 10576 13574 10622 13626
rect 10326 13572 10382 13574
rect 10406 13572 10462 13574
rect 10486 13572 10542 13574
rect 10566 13572 10622 13574
rect 10326 12538 10382 12540
rect 10406 12538 10462 12540
rect 10486 12538 10542 12540
rect 10566 12538 10622 12540
rect 10326 12486 10372 12538
rect 10372 12486 10382 12538
rect 10406 12486 10436 12538
rect 10436 12486 10448 12538
rect 10448 12486 10462 12538
rect 10486 12486 10500 12538
rect 10500 12486 10512 12538
rect 10512 12486 10542 12538
rect 10566 12486 10576 12538
rect 10576 12486 10622 12538
rect 10326 12484 10382 12486
rect 10406 12484 10462 12486
rect 10486 12484 10542 12486
rect 10566 12484 10622 12486
rect 10326 11450 10382 11452
rect 10406 11450 10462 11452
rect 10486 11450 10542 11452
rect 10566 11450 10622 11452
rect 10326 11398 10372 11450
rect 10372 11398 10382 11450
rect 10406 11398 10436 11450
rect 10436 11398 10448 11450
rect 10448 11398 10462 11450
rect 10486 11398 10500 11450
rect 10500 11398 10512 11450
rect 10512 11398 10542 11450
rect 10566 11398 10576 11450
rect 10576 11398 10622 11450
rect 10326 11396 10382 11398
rect 10406 11396 10462 11398
rect 10486 11396 10542 11398
rect 10566 11396 10622 11398
rect 10326 10362 10382 10364
rect 10406 10362 10462 10364
rect 10486 10362 10542 10364
rect 10566 10362 10622 10364
rect 10326 10310 10372 10362
rect 10372 10310 10382 10362
rect 10406 10310 10436 10362
rect 10436 10310 10448 10362
rect 10448 10310 10462 10362
rect 10486 10310 10500 10362
rect 10500 10310 10512 10362
rect 10512 10310 10542 10362
rect 10566 10310 10576 10362
rect 10576 10310 10622 10362
rect 10326 10308 10382 10310
rect 10406 10308 10462 10310
rect 10486 10308 10542 10310
rect 10566 10308 10622 10310
rect 10322 9560 10378 9616
rect 10506 9424 10562 9480
rect 10326 9274 10382 9276
rect 10406 9274 10462 9276
rect 10486 9274 10542 9276
rect 10566 9274 10622 9276
rect 10326 9222 10372 9274
rect 10372 9222 10382 9274
rect 10406 9222 10436 9274
rect 10436 9222 10448 9274
rect 10448 9222 10462 9274
rect 10486 9222 10500 9274
rect 10500 9222 10512 9274
rect 10512 9222 10542 9274
rect 10566 9222 10576 9274
rect 10576 9222 10622 9274
rect 10326 9220 10382 9222
rect 10406 9220 10462 9222
rect 10486 9220 10542 9222
rect 10566 9220 10622 9222
rect 10326 8186 10382 8188
rect 10406 8186 10462 8188
rect 10486 8186 10542 8188
rect 10566 8186 10622 8188
rect 10326 8134 10372 8186
rect 10372 8134 10382 8186
rect 10406 8134 10436 8186
rect 10436 8134 10448 8186
rect 10448 8134 10462 8186
rect 10486 8134 10500 8186
rect 10500 8134 10512 8186
rect 10512 8134 10542 8186
rect 10566 8134 10576 8186
rect 10576 8134 10622 8186
rect 10326 8132 10382 8134
rect 10406 8132 10462 8134
rect 10486 8132 10542 8134
rect 10566 8132 10622 8134
rect 10326 7098 10382 7100
rect 10406 7098 10462 7100
rect 10486 7098 10542 7100
rect 10566 7098 10622 7100
rect 10326 7046 10372 7098
rect 10372 7046 10382 7098
rect 10406 7046 10436 7098
rect 10436 7046 10448 7098
rect 10448 7046 10462 7098
rect 10486 7046 10500 7098
rect 10500 7046 10512 7098
rect 10512 7046 10542 7098
rect 10566 7046 10576 7098
rect 10576 7046 10622 7098
rect 10326 7044 10382 7046
rect 10406 7044 10462 7046
rect 10486 7044 10542 7046
rect 10566 7044 10622 7046
rect 10326 6010 10382 6012
rect 10406 6010 10462 6012
rect 10486 6010 10542 6012
rect 10566 6010 10622 6012
rect 10326 5958 10372 6010
rect 10372 5958 10382 6010
rect 10406 5958 10436 6010
rect 10436 5958 10448 6010
rect 10448 5958 10462 6010
rect 10486 5958 10500 6010
rect 10500 5958 10512 6010
rect 10512 5958 10542 6010
rect 10566 5958 10576 6010
rect 10576 5958 10622 6010
rect 10326 5956 10382 5958
rect 10406 5956 10462 5958
rect 10486 5956 10542 5958
rect 10566 5956 10622 5958
rect 10326 4922 10382 4924
rect 10406 4922 10462 4924
rect 10486 4922 10542 4924
rect 10566 4922 10622 4924
rect 10326 4870 10372 4922
rect 10372 4870 10382 4922
rect 10406 4870 10436 4922
rect 10436 4870 10448 4922
rect 10448 4870 10462 4922
rect 10486 4870 10500 4922
rect 10500 4870 10512 4922
rect 10512 4870 10542 4922
rect 10566 4870 10576 4922
rect 10576 4870 10622 4922
rect 10326 4868 10382 4870
rect 10406 4868 10462 4870
rect 10486 4868 10542 4870
rect 10566 4868 10622 4870
rect 10326 3834 10382 3836
rect 10406 3834 10462 3836
rect 10486 3834 10542 3836
rect 10566 3834 10622 3836
rect 10326 3782 10372 3834
rect 10372 3782 10382 3834
rect 10406 3782 10436 3834
rect 10436 3782 10448 3834
rect 10448 3782 10462 3834
rect 10486 3782 10500 3834
rect 10500 3782 10512 3834
rect 10512 3782 10542 3834
rect 10566 3782 10576 3834
rect 10576 3782 10622 3834
rect 10326 3780 10382 3782
rect 10406 3780 10462 3782
rect 10486 3780 10542 3782
rect 10566 3780 10622 3782
rect 10326 2746 10382 2748
rect 10406 2746 10462 2748
rect 10486 2746 10542 2748
rect 10566 2746 10622 2748
rect 10326 2694 10372 2746
rect 10372 2694 10382 2746
rect 10406 2694 10436 2746
rect 10436 2694 10448 2746
rect 10448 2694 10462 2746
rect 10486 2694 10500 2746
rect 10500 2694 10512 2746
rect 10512 2694 10542 2746
rect 10566 2694 10576 2746
rect 10576 2694 10622 2746
rect 10326 2692 10382 2694
rect 10406 2692 10462 2694
rect 10486 2692 10542 2694
rect 10566 2692 10622 2694
rect 11150 3576 11206 3632
rect 12200 17434 12256 17436
rect 12280 17434 12336 17436
rect 12360 17434 12416 17436
rect 12440 17434 12496 17436
rect 12200 17382 12246 17434
rect 12246 17382 12256 17434
rect 12280 17382 12310 17434
rect 12310 17382 12322 17434
rect 12322 17382 12336 17434
rect 12360 17382 12374 17434
rect 12374 17382 12386 17434
rect 12386 17382 12416 17434
rect 12440 17382 12450 17434
rect 12450 17382 12496 17434
rect 12200 17380 12256 17382
rect 12280 17380 12336 17382
rect 12360 17380 12416 17382
rect 12440 17380 12496 17382
rect 12200 16346 12256 16348
rect 12280 16346 12336 16348
rect 12360 16346 12416 16348
rect 12440 16346 12496 16348
rect 12200 16294 12246 16346
rect 12246 16294 12256 16346
rect 12280 16294 12310 16346
rect 12310 16294 12322 16346
rect 12322 16294 12336 16346
rect 12360 16294 12374 16346
rect 12374 16294 12386 16346
rect 12386 16294 12416 16346
rect 12440 16294 12450 16346
rect 12450 16294 12496 16346
rect 12200 16292 12256 16294
rect 12280 16292 12336 16294
rect 12360 16292 12416 16294
rect 12440 16292 12496 16294
rect 12200 15258 12256 15260
rect 12280 15258 12336 15260
rect 12360 15258 12416 15260
rect 12440 15258 12496 15260
rect 12200 15206 12246 15258
rect 12246 15206 12256 15258
rect 12280 15206 12310 15258
rect 12310 15206 12322 15258
rect 12322 15206 12336 15258
rect 12360 15206 12374 15258
rect 12374 15206 12386 15258
rect 12386 15206 12416 15258
rect 12440 15206 12450 15258
rect 12450 15206 12496 15258
rect 12200 15204 12256 15206
rect 12280 15204 12336 15206
rect 12360 15204 12416 15206
rect 12440 15204 12496 15206
rect 12200 14170 12256 14172
rect 12280 14170 12336 14172
rect 12360 14170 12416 14172
rect 12440 14170 12496 14172
rect 12200 14118 12246 14170
rect 12246 14118 12256 14170
rect 12280 14118 12310 14170
rect 12310 14118 12322 14170
rect 12322 14118 12336 14170
rect 12360 14118 12374 14170
rect 12374 14118 12386 14170
rect 12386 14118 12416 14170
rect 12440 14118 12450 14170
rect 12450 14118 12496 14170
rect 12200 14116 12256 14118
rect 12280 14116 12336 14118
rect 12360 14116 12416 14118
rect 12440 14116 12496 14118
rect 12200 13082 12256 13084
rect 12280 13082 12336 13084
rect 12360 13082 12416 13084
rect 12440 13082 12496 13084
rect 12200 13030 12246 13082
rect 12246 13030 12256 13082
rect 12280 13030 12310 13082
rect 12310 13030 12322 13082
rect 12322 13030 12336 13082
rect 12360 13030 12374 13082
rect 12374 13030 12386 13082
rect 12386 13030 12416 13082
rect 12440 13030 12450 13082
rect 12450 13030 12496 13082
rect 12200 13028 12256 13030
rect 12280 13028 12336 13030
rect 12360 13028 12416 13030
rect 12440 13028 12496 13030
rect 12438 12688 12494 12744
rect 12200 11994 12256 11996
rect 12280 11994 12336 11996
rect 12360 11994 12416 11996
rect 12440 11994 12496 11996
rect 12200 11942 12246 11994
rect 12246 11942 12256 11994
rect 12280 11942 12310 11994
rect 12310 11942 12322 11994
rect 12322 11942 12336 11994
rect 12360 11942 12374 11994
rect 12374 11942 12386 11994
rect 12386 11942 12416 11994
rect 12440 11942 12450 11994
rect 12450 11942 12496 11994
rect 12200 11940 12256 11942
rect 12280 11940 12336 11942
rect 12360 11940 12416 11942
rect 12440 11940 12496 11942
rect 12200 10906 12256 10908
rect 12280 10906 12336 10908
rect 12360 10906 12416 10908
rect 12440 10906 12496 10908
rect 12200 10854 12246 10906
rect 12246 10854 12256 10906
rect 12280 10854 12310 10906
rect 12310 10854 12322 10906
rect 12322 10854 12336 10906
rect 12360 10854 12374 10906
rect 12374 10854 12386 10906
rect 12386 10854 12416 10906
rect 12440 10854 12450 10906
rect 12450 10854 12496 10906
rect 12200 10852 12256 10854
rect 12280 10852 12336 10854
rect 12360 10852 12416 10854
rect 12440 10852 12496 10854
rect 12200 9818 12256 9820
rect 12280 9818 12336 9820
rect 12360 9818 12416 9820
rect 12440 9818 12496 9820
rect 12200 9766 12246 9818
rect 12246 9766 12256 9818
rect 12280 9766 12310 9818
rect 12310 9766 12322 9818
rect 12322 9766 12336 9818
rect 12360 9766 12374 9818
rect 12374 9766 12386 9818
rect 12386 9766 12416 9818
rect 12440 9766 12450 9818
rect 12450 9766 12496 9818
rect 12200 9764 12256 9766
rect 12280 9764 12336 9766
rect 12360 9764 12416 9766
rect 12440 9764 12496 9766
rect 12200 8730 12256 8732
rect 12280 8730 12336 8732
rect 12360 8730 12416 8732
rect 12440 8730 12496 8732
rect 12200 8678 12246 8730
rect 12246 8678 12256 8730
rect 12280 8678 12310 8730
rect 12310 8678 12322 8730
rect 12322 8678 12336 8730
rect 12360 8678 12374 8730
rect 12374 8678 12386 8730
rect 12386 8678 12416 8730
rect 12440 8678 12450 8730
rect 12450 8678 12496 8730
rect 12200 8676 12256 8678
rect 12280 8676 12336 8678
rect 12360 8676 12416 8678
rect 12440 8676 12496 8678
rect 12200 7642 12256 7644
rect 12280 7642 12336 7644
rect 12360 7642 12416 7644
rect 12440 7642 12496 7644
rect 12200 7590 12246 7642
rect 12246 7590 12256 7642
rect 12280 7590 12310 7642
rect 12310 7590 12322 7642
rect 12322 7590 12336 7642
rect 12360 7590 12374 7642
rect 12374 7590 12386 7642
rect 12386 7590 12416 7642
rect 12440 7590 12450 7642
rect 12450 7590 12496 7642
rect 12200 7588 12256 7590
rect 12280 7588 12336 7590
rect 12360 7588 12416 7590
rect 12440 7588 12496 7590
rect 12200 6554 12256 6556
rect 12280 6554 12336 6556
rect 12360 6554 12416 6556
rect 12440 6554 12496 6556
rect 12200 6502 12246 6554
rect 12246 6502 12256 6554
rect 12280 6502 12310 6554
rect 12310 6502 12322 6554
rect 12322 6502 12336 6554
rect 12360 6502 12374 6554
rect 12374 6502 12386 6554
rect 12386 6502 12416 6554
rect 12440 6502 12450 6554
rect 12450 6502 12496 6554
rect 12200 6500 12256 6502
rect 12280 6500 12336 6502
rect 12360 6500 12416 6502
rect 12440 6500 12496 6502
rect 12200 5466 12256 5468
rect 12280 5466 12336 5468
rect 12360 5466 12416 5468
rect 12440 5466 12496 5468
rect 12200 5414 12246 5466
rect 12246 5414 12256 5466
rect 12280 5414 12310 5466
rect 12310 5414 12322 5466
rect 12322 5414 12336 5466
rect 12360 5414 12374 5466
rect 12374 5414 12386 5466
rect 12386 5414 12416 5466
rect 12440 5414 12450 5466
rect 12450 5414 12496 5466
rect 12200 5412 12256 5414
rect 12280 5412 12336 5414
rect 12360 5412 12416 5414
rect 12440 5412 12496 5414
rect 12200 4378 12256 4380
rect 12280 4378 12336 4380
rect 12360 4378 12416 4380
rect 12440 4378 12496 4380
rect 12200 4326 12246 4378
rect 12246 4326 12256 4378
rect 12280 4326 12310 4378
rect 12310 4326 12322 4378
rect 12322 4326 12336 4378
rect 12360 4326 12374 4378
rect 12374 4326 12386 4378
rect 12386 4326 12416 4378
rect 12440 4326 12450 4378
rect 12450 4326 12496 4378
rect 12200 4324 12256 4326
rect 12280 4324 12336 4326
rect 12360 4324 12416 4326
rect 12440 4324 12496 4326
rect 13726 17312 13782 17368
rect 14074 16890 14130 16892
rect 14154 16890 14210 16892
rect 14234 16890 14290 16892
rect 14314 16890 14370 16892
rect 14074 16838 14120 16890
rect 14120 16838 14130 16890
rect 14154 16838 14184 16890
rect 14184 16838 14196 16890
rect 14196 16838 14210 16890
rect 14234 16838 14248 16890
rect 14248 16838 14260 16890
rect 14260 16838 14290 16890
rect 14314 16838 14324 16890
rect 14324 16838 14370 16890
rect 14074 16836 14130 16838
rect 14154 16836 14210 16838
rect 14234 16836 14290 16838
rect 14314 16836 14370 16838
rect 14074 15802 14130 15804
rect 14154 15802 14210 15804
rect 14234 15802 14290 15804
rect 14314 15802 14370 15804
rect 14074 15750 14120 15802
rect 14120 15750 14130 15802
rect 14154 15750 14184 15802
rect 14184 15750 14196 15802
rect 14196 15750 14210 15802
rect 14234 15750 14248 15802
rect 14248 15750 14260 15802
rect 14260 15750 14290 15802
rect 14314 15750 14324 15802
rect 14324 15750 14370 15802
rect 14074 15748 14130 15750
rect 14154 15748 14210 15750
rect 14234 15748 14290 15750
rect 14314 15748 14370 15750
rect 14074 14714 14130 14716
rect 14154 14714 14210 14716
rect 14234 14714 14290 14716
rect 14314 14714 14370 14716
rect 14074 14662 14120 14714
rect 14120 14662 14130 14714
rect 14154 14662 14184 14714
rect 14184 14662 14196 14714
rect 14196 14662 14210 14714
rect 14234 14662 14248 14714
rect 14248 14662 14260 14714
rect 14260 14662 14290 14714
rect 14314 14662 14324 14714
rect 14324 14662 14370 14714
rect 14074 14660 14130 14662
rect 14154 14660 14210 14662
rect 14234 14660 14290 14662
rect 14314 14660 14370 14662
rect 14074 13626 14130 13628
rect 14154 13626 14210 13628
rect 14234 13626 14290 13628
rect 14314 13626 14370 13628
rect 14074 13574 14120 13626
rect 14120 13574 14130 13626
rect 14154 13574 14184 13626
rect 14184 13574 14196 13626
rect 14196 13574 14210 13626
rect 14234 13574 14248 13626
rect 14248 13574 14260 13626
rect 14260 13574 14290 13626
rect 14314 13574 14324 13626
rect 14324 13574 14370 13626
rect 14074 13572 14130 13574
rect 14154 13572 14210 13574
rect 14234 13572 14290 13574
rect 14314 13572 14370 13574
rect 14074 12538 14130 12540
rect 14154 12538 14210 12540
rect 14234 12538 14290 12540
rect 14314 12538 14370 12540
rect 14074 12486 14120 12538
rect 14120 12486 14130 12538
rect 14154 12486 14184 12538
rect 14184 12486 14196 12538
rect 14196 12486 14210 12538
rect 14234 12486 14248 12538
rect 14248 12486 14260 12538
rect 14260 12486 14290 12538
rect 14314 12486 14324 12538
rect 14324 12486 14370 12538
rect 14074 12484 14130 12486
rect 14154 12484 14210 12486
rect 14234 12484 14290 12486
rect 14314 12484 14370 12486
rect 14074 11450 14130 11452
rect 14154 11450 14210 11452
rect 14234 11450 14290 11452
rect 14314 11450 14370 11452
rect 14074 11398 14120 11450
rect 14120 11398 14130 11450
rect 14154 11398 14184 11450
rect 14184 11398 14196 11450
rect 14196 11398 14210 11450
rect 14234 11398 14248 11450
rect 14248 11398 14260 11450
rect 14260 11398 14290 11450
rect 14314 11398 14324 11450
rect 14324 11398 14370 11450
rect 14074 11396 14130 11398
rect 14154 11396 14210 11398
rect 14234 11396 14290 11398
rect 14314 11396 14370 11398
rect 14074 10362 14130 10364
rect 14154 10362 14210 10364
rect 14234 10362 14290 10364
rect 14314 10362 14370 10364
rect 14074 10310 14120 10362
rect 14120 10310 14130 10362
rect 14154 10310 14184 10362
rect 14184 10310 14196 10362
rect 14196 10310 14210 10362
rect 14234 10310 14248 10362
rect 14248 10310 14260 10362
rect 14260 10310 14290 10362
rect 14314 10310 14324 10362
rect 14324 10310 14370 10362
rect 14074 10308 14130 10310
rect 14154 10308 14210 10310
rect 14234 10308 14290 10310
rect 14314 10308 14370 10310
rect 14646 9968 14702 10024
rect 12714 7520 12770 7576
rect 12530 3984 12586 4040
rect 12200 3290 12256 3292
rect 12280 3290 12336 3292
rect 12360 3290 12416 3292
rect 12440 3290 12496 3292
rect 12200 3238 12246 3290
rect 12246 3238 12256 3290
rect 12280 3238 12310 3290
rect 12310 3238 12322 3290
rect 12322 3238 12336 3290
rect 12360 3238 12374 3290
rect 12374 3238 12386 3290
rect 12386 3238 12416 3290
rect 12440 3238 12450 3290
rect 12450 3238 12496 3290
rect 12200 3236 12256 3238
rect 12280 3236 12336 3238
rect 12360 3236 12416 3238
rect 12440 3236 12496 3238
rect 12438 2488 12494 2544
rect 12200 2202 12256 2204
rect 12280 2202 12336 2204
rect 12360 2202 12416 2204
rect 12440 2202 12496 2204
rect 12200 2150 12246 2202
rect 12246 2150 12256 2202
rect 12280 2150 12310 2202
rect 12310 2150 12322 2202
rect 12322 2150 12336 2202
rect 12360 2150 12374 2202
rect 12374 2150 12386 2202
rect 12386 2150 12416 2202
rect 12440 2150 12450 2202
rect 12450 2150 12496 2202
rect 12200 2148 12256 2150
rect 12280 2148 12336 2150
rect 12360 2148 12416 2150
rect 12440 2148 12496 2150
rect 14074 9274 14130 9276
rect 14154 9274 14210 9276
rect 14234 9274 14290 9276
rect 14314 9274 14370 9276
rect 14074 9222 14120 9274
rect 14120 9222 14130 9274
rect 14154 9222 14184 9274
rect 14184 9222 14196 9274
rect 14196 9222 14210 9274
rect 14234 9222 14248 9274
rect 14248 9222 14260 9274
rect 14260 9222 14290 9274
rect 14314 9222 14324 9274
rect 14324 9222 14370 9274
rect 14074 9220 14130 9222
rect 14154 9220 14210 9222
rect 14234 9220 14290 9222
rect 14314 9220 14370 9222
rect 14074 8186 14130 8188
rect 14154 8186 14210 8188
rect 14234 8186 14290 8188
rect 14314 8186 14370 8188
rect 14074 8134 14120 8186
rect 14120 8134 14130 8186
rect 14154 8134 14184 8186
rect 14184 8134 14196 8186
rect 14196 8134 14210 8186
rect 14234 8134 14248 8186
rect 14248 8134 14260 8186
rect 14260 8134 14290 8186
rect 14314 8134 14324 8186
rect 14324 8134 14370 8186
rect 14074 8132 14130 8134
rect 14154 8132 14210 8134
rect 14234 8132 14290 8134
rect 14314 8132 14370 8134
rect 14074 7098 14130 7100
rect 14154 7098 14210 7100
rect 14234 7098 14290 7100
rect 14314 7098 14370 7100
rect 14074 7046 14120 7098
rect 14120 7046 14130 7098
rect 14154 7046 14184 7098
rect 14184 7046 14196 7098
rect 14196 7046 14210 7098
rect 14234 7046 14248 7098
rect 14248 7046 14260 7098
rect 14260 7046 14290 7098
rect 14314 7046 14324 7098
rect 14324 7046 14370 7098
rect 14074 7044 14130 7046
rect 14154 7044 14210 7046
rect 14234 7044 14290 7046
rect 14314 7044 14370 7046
rect 14074 6010 14130 6012
rect 14154 6010 14210 6012
rect 14234 6010 14290 6012
rect 14314 6010 14370 6012
rect 14074 5958 14120 6010
rect 14120 5958 14130 6010
rect 14154 5958 14184 6010
rect 14184 5958 14196 6010
rect 14196 5958 14210 6010
rect 14234 5958 14248 6010
rect 14248 5958 14260 6010
rect 14260 5958 14290 6010
rect 14314 5958 14324 6010
rect 14324 5958 14370 6010
rect 14074 5956 14130 5958
rect 14154 5956 14210 5958
rect 14234 5956 14290 5958
rect 14314 5956 14370 5958
rect 14074 4922 14130 4924
rect 14154 4922 14210 4924
rect 14234 4922 14290 4924
rect 14314 4922 14370 4924
rect 14074 4870 14120 4922
rect 14120 4870 14130 4922
rect 14154 4870 14184 4922
rect 14184 4870 14196 4922
rect 14196 4870 14210 4922
rect 14234 4870 14248 4922
rect 14248 4870 14260 4922
rect 14260 4870 14290 4922
rect 14314 4870 14324 4922
rect 14324 4870 14370 4922
rect 14074 4868 14130 4870
rect 14154 4868 14210 4870
rect 14234 4868 14290 4870
rect 14314 4868 14370 4870
rect 14074 3834 14130 3836
rect 14154 3834 14210 3836
rect 14234 3834 14290 3836
rect 14314 3834 14370 3836
rect 14074 3782 14120 3834
rect 14120 3782 14130 3834
rect 14154 3782 14184 3834
rect 14184 3782 14196 3834
rect 14196 3782 14210 3834
rect 14234 3782 14248 3834
rect 14248 3782 14260 3834
rect 14260 3782 14290 3834
rect 14314 3782 14324 3834
rect 14324 3782 14370 3834
rect 14074 3780 14130 3782
rect 14154 3780 14210 3782
rect 14234 3780 14290 3782
rect 14314 3780 14370 3782
rect 14074 2746 14130 2748
rect 14154 2746 14210 2748
rect 14234 2746 14290 2748
rect 14314 2746 14370 2748
rect 14074 2694 14120 2746
rect 14120 2694 14130 2746
rect 14154 2694 14184 2746
rect 14184 2694 14196 2746
rect 14196 2694 14210 2746
rect 14234 2694 14248 2746
rect 14248 2694 14260 2746
rect 14260 2694 14290 2746
rect 14314 2694 14324 2746
rect 14324 2694 14370 2746
rect 14074 2692 14130 2694
rect 14154 2692 14210 2694
rect 14234 2692 14290 2694
rect 14314 2692 14370 2694
<< metal3 >>
rect 0 18186 800 18216
rect 4061 18186 4127 18189
rect 0 18184 4127 18186
rect 0 18128 4066 18184
rect 4122 18128 4127 18184
rect 0 18126 4127 18128
rect 0 18096 800 18126
rect 4061 18123 4127 18126
rect 4694 17440 5010 17441
rect 4694 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5010 17440
rect 4694 17375 5010 17376
rect 8442 17440 8758 17441
rect 8442 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8758 17440
rect 8442 17375 8758 17376
rect 12190 17440 12506 17441
rect 12190 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12506 17440
rect 12190 17375 12506 17376
rect 13721 17370 13787 17373
rect 16400 17370 17200 17400
rect 13721 17368 17200 17370
rect 13721 17312 13726 17368
rect 13782 17312 17200 17368
rect 13721 17310 17200 17312
rect 13721 17307 13787 17310
rect 16400 17280 17200 17310
rect 2820 16896 3136 16897
rect 2820 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3136 16896
rect 2820 16831 3136 16832
rect 6568 16896 6884 16897
rect 6568 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6884 16896
rect 6568 16831 6884 16832
rect 10316 16896 10632 16897
rect 10316 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10632 16896
rect 10316 16831 10632 16832
rect 14064 16896 14380 16897
rect 14064 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14380 16896
rect 14064 16831 14380 16832
rect 4694 16352 5010 16353
rect 4694 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5010 16352
rect 4694 16287 5010 16288
rect 8442 16352 8758 16353
rect 8442 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8758 16352
rect 8442 16287 8758 16288
rect 12190 16352 12506 16353
rect 12190 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12506 16352
rect 12190 16287 12506 16288
rect 2820 15808 3136 15809
rect 2820 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3136 15808
rect 2820 15743 3136 15744
rect 6568 15808 6884 15809
rect 6568 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6884 15808
rect 6568 15743 6884 15744
rect 10316 15808 10632 15809
rect 10316 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10632 15808
rect 10316 15743 10632 15744
rect 14064 15808 14380 15809
rect 14064 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14380 15808
rect 14064 15743 14380 15744
rect 4694 15264 5010 15265
rect 4694 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5010 15264
rect 4694 15199 5010 15200
rect 8442 15264 8758 15265
rect 8442 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8758 15264
rect 8442 15199 8758 15200
rect 12190 15264 12506 15265
rect 12190 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12506 15264
rect 12190 15199 12506 15200
rect 0 14922 800 14952
rect 1761 14922 1827 14925
rect 0 14920 1827 14922
rect 0 14864 1766 14920
rect 1822 14864 1827 14920
rect 0 14862 1827 14864
rect 0 14832 800 14862
rect 1761 14859 1827 14862
rect 2820 14720 3136 14721
rect 2820 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3136 14720
rect 2820 14655 3136 14656
rect 6568 14720 6884 14721
rect 6568 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6884 14720
rect 6568 14655 6884 14656
rect 10316 14720 10632 14721
rect 10316 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10632 14720
rect 10316 14655 10632 14656
rect 14064 14720 14380 14721
rect 14064 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14380 14720
rect 14064 14655 14380 14656
rect 4694 14176 5010 14177
rect 4694 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5010 14176
rect 4694 14111 5010 14112
rect 8442 14176 8758 14177
rect 8442 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8758 14176
rect 8442 14111 8758 14112
rect 12190 14176 12506 14177
rect 12190 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12506 14176
rect 12190 14111 12506 14112
rect 2820 13632 3136 13633
rect 2820 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3136 13632
rect 2820 13567 3136 13568
rect 6568 13632 6884 13633
rect 6568 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6884 13632
rect 6568 13567 6884 13568
rect 10316 13632 10632 13633
rect 10316 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10632 13632
rect 10316 13567 10632 13568
rect 14064 13632 14380 13633
rect 14064 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14380 13632
rect 14064 13567 14380 13568
rect 4694 13088 5010 13089
rect 4694 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5010 13088
rect 4694 13023 5010 13024
rect 8442 13088 8758 13089
rect 8442 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8758 13088
rect 8442 13023 8758 13024
rect 12190 13088 12506 13089
rect 12190 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12506 13088
rect 12190 13023 12506 13024
rect 12433 12746 12499 12749
rect 12433 12744 14658 12746
rect 12433 12688 12438 12744
rect 12494 12688 14658 12744
rect 12433 12686 14658 12688
rect 12433 12683 12499 12686
rect 2820 12544 3136 12545
rect 2820 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3136 12544
rect 2820 12479 3136 12480
rect 6568 12544 6884 12545
rect 6568 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6884 12544
rect 6568 12479 6884 12480
rect 10316 12544 10632 12545
rect 10316 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10632 12544
rect 10316 12479 10632 12480
rect 14064 12544 14380 12545
rect 14064 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14380 12544
rect 14064 12479 14380 12480
rect 14598 12474 14658 12686
rect 16400 12474 17200 12504
rect 14598 12414 17200 12474
rect 16400 12384 17200 12414
rect 4694 12000 5010 12001
rect 4694 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5010 12000
rect 4694 11935 5010 11936
rect 8442 12000 8758 12001
rect 8442 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8758 12000
rect 8442 11935 8758 11936
rect 12190 12000 12506 12001
rect 12190 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12506 12000
rect 12190 11935 12506 11936
rect 0 11658 800 11688
rect 4153 11658 4219 11661
rect 0 11656 4219 11658
rect 0 11600 4158 11656
rect 4214 11600 4219 11656
rect 0 11598 4219 11600
rect 0 11568 800 11598
rect 4153 11595 4219 11598
rect 2820 11456 3136 11457
rect 2820 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3136 11456
rect 2820 11391 3136 11392
rect 6568 11456 6884 11457
rect 6568 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6884 11456
rect 6568 11391 6884 11392
rect 10316 11456 10632 11457
rect 10316 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10632 11456
rect 10316 11391 10632 11392
rect 14064 11456 14380 11457
rect 14064 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14380 11456
rect 14064 11391 14380 11392
rect 5533 11386 5599 11389
rect 5717 11386 5783 11389
rect 5533 11384 5783 11386
rect 5533 11328 5538 11384
rect 5594 11328 5722 11384
rect 5778 11328 5783 11384
rect 5533 11326 5783 11328
rect 5533 11323 5599 11326
rect 5717 11323 5783 11326
rect 8886 11188 8892 11252
rect 8956 11250 8962 11252
rect 9029 11250 9095 11253
rect 8956 11248 9095 11250
rect 8956 11192 9034 11248
rect 9090 11192 9095 11248
rect 8956 11190 9095 11192
rect 8956 11188 8962 11190
rect 9029 11187 9095 11190
rect 4694 10912 5010 10913
rect 4694 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5010 10912
rect 4694 10847 5010 10848
rect 8442 10912 8758 10913
rect 8442 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8758 10912
rect 8442 10847 8758 10848
rect 12190 10912 12506 10913
rect 12190 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12506 10912
rect 12190 10847 12506 10848
rect 2820 10368 3136 10369
rect 2820 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3136 10368
rect 2820 10303 3136 10304
rect 6568 10368 6884 10369
rect 6568 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6884 10368
rect 6568 10303 6884 10304
rect 10316 10368 10632 10369
rect 10316 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10632 10368
rect 10316 10303 10632 10304
rect 14064 10368 14380 10369
rect 14064 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14380 10368
rect 14064 10303 14380 10304
rect 7741 10162 7807 10165
rect 9029 10162 9095 10165
rect 7741 10160 9095 10162
rect 7741 10104 7746 10160
rect 7802 10104 9034 10160
rect 9090 10104 9095 10160
rect 7741 10102 9095 10104
rect 7741 10099 7807 10102
rect 9029 10099 9095 10102
rect 6821 10026 6887 10029
rect 14641 10026 14707 10029
rect 6821 10024 14707 10026
rect 6821 9968 6826 10024
rect 6882 9968 14646 10024
rect 14702 9968 14707 10024
rect 6821 9966 14707 9968
rect 6821 9963 6887 9966
rect 14641 9963 14707 9966
rect 4694 9824 5010 9825
rect 4694 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5010 9824
rect 4694 9759 5010 9760
rect 8442 9824 8758 9825
rect 8442 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8758 9824
rect 8442 9759 8758 9760
rect 12190 9824 12506 9825
rect 12190 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12506 9824
rect 12190 9759 12506 9760
rect 8845 9756 8911 9757
rect 8845 9752 8892 9756
rect 8956 9754 8962 9756
rect 8845 9696 8850 9752
rect 8845 9692 8892 9696
rect 8956 9694 9002 9754
rect 8956 9692 8962 9694
rect 8845 9691 8911 9692
rect 5625 9618 5691 9621
rect 10317 9618 10383 9621
rect 5625 9616 10383 9618
rect 5625 9560 5630 9616
rect 5686 9560 10322 9616
rect 10378 9560 10383 9616
rect 5625 9558 10383 9560
rect 5625 9555 5691 9558
rect 10317 9555 10383 9558
rect 5993 9482 6059 9485
rect 9765 9482 9831 9485
rect 10501 9482 10567 9485
rect 5993 9480 9831 9482
rect 5993 9424 5998 9480
rect 6054 9424 9770 9480
rect 9826 9424 9831 9480
rect 5993 9422 9831 9424
rect 5993 9419 6059 9422
rect 9765 9419 9831 9422
rect 9998 9480 10567 9482
rect 9998 9424 10506 9480
rect 10562 9424 10567 9480
rect 9998 9422 10567 9424
rect 7741 9346 7807 9349
rect 8477 9346 8543 9349
rect 7741 9344 8543 9346
rect 7741 9288 7746 9344
rect 7802 9288 8482 9344
rect 8538 9288 8543 9344
rect 7741 9286 8543 9288
rect 7741 9283 7807 9286
rect 8477 9283 8543 9286
rect 9029 9346 9095 9349
rect 9397 9346 9463 9349
rect 9029 9344 9463 9346
rect 9029 9288 9034 9344
rect 9090 9288 9402 9344
rect 9458 9288 9463 9344
rect 9029 9286 9463 9288
rect 9029 9283 9095 9286
rect 9397 9283 9463 9286
rect 2820 9280 3136 9281
rect 2820 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3136 9280
rect 2820 9215 3136 9216
rect 6568 9280 6884 9281
rect 6568 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6884 9280
rect 6568 9215 6884 9216
rect 8201 9210 8267 9213
rect 8661 9210 8727 9213
rect 8201 9208 8727 9210
rect 8201 9152 8206 9208
rect 8262 9152 8666 9208
rect 8722 9152 8727 9208
rect 8201 9150 8727 9152
rect 8201 9147 8267 9150
rect 8661 9147 8727 9150
rect 6177 9074 6243 9077
rect 9998 9074 10058 9422
rect 10501 9419 10567 9422
rect 10316 9280 10632 9281
rect 10316 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10632 9280
rect 10316 9215 10632 9216
rect 14064 9280 14380 9281
rect 14064 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14380 9280
rect 14064 9215 14380 9216
rect 6177 9072 10058 9074
rect 6177 9016 6182 9072
rect 6238 9016 10058 9072
rect 6177 9014 10058 9016
rect 6177 9011 6243 9014
rect 5993 8938 6059 8941
rect 9029 8938 9095 8941
rect 5993 8936 9095 8938
rect 5993 8880 5998 8936
rect 6054 8880 9034 8936
rect 9090 8880 9095 8936
rect 5993 8878 9095 8880
rect 5993 8875 6059 8878
rect 9029 8875 9095 8878
rect 4694 8736 5010 8737
rect 4694 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5010 8736
rect 4694 8671 5010 8672
rect 8442 8736 8758 8737
rect 8442 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8758 8736
rect 8442 8671 8758 8672
rect 12190 8736 12506 8737
rect 12190 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12506 8736
rect 12190 8671 12506 8672
rect 0 8394 800 8424
rect 3233 8394 3299 8397
rect 0 8392 3299 8394
rect 0 8336 3238 8392
rect 3294 8336 3299 8392
rect 0 8334 3299 8336
rect 0 8304 800 8334
rect 3233 8331 3299 8334
rect 2820 8192 3136 8193
rect 2820 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3136 8192
rect 2820 8127 3136 8128
rect 6568 8192 6884 8193
rect 6568 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6884 8192
rect 6568 8127 6884 8128
rect 10316 8192 10632 8193
rect 10316 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10632 8192
rect 10316 8127 10632 8128
rect 14064 8192 14380 8193
rect 14064 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14380 8192
rect 14064 8127 14380 8128
rect 4694 7648 5010 7649
rect 4694 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5010 7648
rect 4694 7583 5010 7584
rect 8442 7648 8758 7649
rect 8442 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8758 7648
rect 8442 7583 8758 7584
rect 12190 7648 12506 7649
rect 12190 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12506 7648
rect 12190 7583 12506 7584
rect 12709 7578 12775 7581
rect 16400 7578 17200 7608
rect 12709 7576 17200 7578
rect 12709 7520 12714 7576
rect 12770 7520 17200 7576
rect 12709 7518 17200 7520
rect 12709 7515 12775 7518
rect 16400 7488 17200 7518
rect 2820 7104 3136 7105
rect 2820 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3136 7104
rect 2820 7039 3136 7040
rect 6568 7104 6884 7105
rect 6568 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6884 7104
rect 6568 7039 6884 7040
rect 10316 7104 10632 7105
rect 10316 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10632 7104
rect 10316 7039 10632 7040
rect 14064 7104 14380 7105
rect 14064 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14380 7104
rect 14064 7039 14380 7040
rect 4694 6560 5010 6561
rect 4694 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5010 6560
rect 4694 6495 5010 6496
rect 8442 6560 8758 6561
rect 8442 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8758 6560
rect 8442 6495 8758 6496
rect 12190 6560 12506 6561
rect 12190 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12506 6560
rect 12190 6495 12506 6496
rect 2820 6016 3136 6017
rect 2820 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3136 6016
rect 2820 5951 3136 5952
rect 6568 6016 6884 6017
rect 6568 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6884 6016
rect 6568 5951 6884 5952
rect 10316 6016 10632 6017
rect 10316 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10632 6016
rect 10316 5951 10632 5952
rect 14064 6016 14380 6017
rect 14064 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14380 6016
rect 14064 5951 14380 5952
rect 4694 5472 5010 5473
rect 4694 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5010 5472
rect 4694 5407 5010 5408
rect 8442 5472 8758 5473
rect 8442 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8758 5472
rect 8442 5407 8758 5408
rect 12190 5472 12506 5473
rect 12190 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12506 5472
rect 12190 5407 12506 5408
rect 0 5130 800 5160
rect 3233 5130 3299 5133
rect 0 5128 3299 5130
rect 0 5072 3238 5128
rect 3294 5072 3299 5128
rect 0 5070 3299 5072
rect 0 5040 800 5070
rect 3233 5067 3299 5070
rect 2820 4928 3136 4929
rect 2820 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3136 4928
rect 2820 4863 3136 4864
rect 6568 4928 6884 4929
rect 6568 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6884 4928
rect 6568 4863 6884 4864
rect 10316 4928 10632 4929
rect 10316 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10632 4928
rect 10316 4863 10632 4864
rect 14064 4928 14380 4929
rect 14064 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14380 4928
rect 14064 4863 14380 4864
rect 4694 4384 5010 4385
rect 4694 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5010 4384
rect 4694 4319 5010 4320
rect 8442 4384 8758 4385
rect 8442 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8758 4384
rect 8442 4319 8758 4320
rect 12190 4384 12506 4385
rect 12190 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12506 4384
rect 12190 4319 12506 4320
rect 8017 4042 8083 4045
rect 12525 4042 12591 4045
rect 8017 4040 12591 4042
rect 8017 3984 8022 4040
rect 8078 3984 12530 4040
rect 12586 3984 12591 4040
rect 8017 3982 12591 3984
rect 8017 3979 8083 3982
rect 12525 3979 12591 3982
rect 2820 3840 3136 3841
rect 2820 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3136 3840
rect 2820 3775 3136 3776
rect 6568 3840 6884 3841
rect 6568 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6884 3840
rect 6568 3775 6884 3776
rect 10316 3840 10632 3841
rect 10316 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10632 3840
rect 10316 3775 10632 3776
rect 14064 3840 14380 3841
rect 14064 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14380 3840
rect 14064 3775 14380 3776
rect 6453 3634 6519 3637
rect 11145 3634 11211 3637
rect 6453 3632 11211 3634
rect 6453 3576 6458 3632
rect 6514 3576 11150 3632
rect 11206 3576 11211 3632
rect 6453 3574 11211 3576
rect 6453 3571 6519 3574
rect 11145 3571 11211 3574
rect 4694 3296 5010 3297
rect 4694 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5010 3296
rect 4694 3231 5010 3232
rect 8442 3296 8758 3297
rect 8442 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8758 3296
rect 8442 3231 8758 3232
rect 12190 3296 12506 3297
rect 12190 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12506 3296
rect 12190 3231 12506 3232
rect 2820 2752 3136 2753
rect 2820 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3136 2752
rect 2820 2687 3136 2688
rect 6568 2752 6884 2753
rect 6568 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6884 2752
rect 6568 2687 6884 2688
rect 10316 2752 10632 2753
rect 10316 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10632 2752
rect 10316 2687 10632 2688
rect 14064 2752 14380 2753
rect 14064 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14380 2752
rect 14064 2687 14380 2688
rect 16400 2682 17200 2712
rect 14598 2622 17200 2682
rect 12433 2546 12499 2549
rect 14598 2546 14658 2622
rect 16400 2592 17200 2622
rect 12433 2544 14658 2546
rect 12433 2488 12438 2544
rect 12494 2488 14658 2544
rect 12433 2486 14658 2488
rect 12433 2483 12499 2486
rect 4694 2208 5010 2209
rect 4694 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5010 2208
rect 4694 2143 5010 2144
rect 8442 2208 8758 2209
rect 8442 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8758 2208
rect 8442 2143 8758 2144
rect 12190 2208 12506 2209
rect 12190 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12506 2208
rect 12190 2143 12506 2144
rect 0 1866 800 1896
rect 3141 1866 3207 1869
rect 0 1864 3207 1866
rect 0 1808 3146 1864
rect 3202 1808 3207 1864
rect 0 1806 3207 1808
rect 0 1776 800 1806
rect 3141 1803 3207 1806
<< via3 >>
rect 4700 17436 4764 17440
rect 4700 17380 4704 17436
rect 4704 17380 4760 17436
rect 4760 17380 4764 17436
rect 4700 17376 4764 17380
rect 4780 17436 4844 17440
rect 4780 17380 4784 17436
rect 4784 17380 4840 17436
rect 4840 17380 4844 17436
rect 4780 17376 4844 17380
rect 4860 17436 4924 17440
rect 4860 17380 4864 17436
rect 4864 17380 4920 17436
rect 4920 17380 4924 17436
rect 4860 17376 4924 17380
rect 4940 17436 5004 17440
rect 4940 17380 4944 17436
rect 4944 17380 5000 17436
rect 5000 17380 5004 17436
rect 4940 17376 5004 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 12196 17436 12260 17440
rect 12196 17380 12200 17436
rect 12200 17380 12256 17436
rect 12256 17380 12260 17436
rect 12196 17376 12260 17380
rect 12276 17436 12340 17440
rect 12276 17380 12280 17436
rect 12280 17380 12336 17436
rect 12336 17380 12340 17436
rect 12276 17376 12340 17380
rect 12356 17436 12420 17440
rect 12356 17380 12360 17436
rect 12360 17380 12416 17436
rect 12416 17380 12420 17436
rect 12356 17376 12420 17380
rect 12436 17436 12500 17440
rect 12436 17380 12440 17436
rect 12440 17380 12496 17436
rect 12496 17380 12500 17436
rect 12436 17376 12500 17380
rect 2826 16892 2890 16896
rect 2826 16836 2830 16892
rect 2830 16836 2886 16892
rect 2886 16836 2890 16892
rect 2826 16832 2890 16836
rect 2906 16892 2970 16896
rect 2906 16836 2910 16892
rect 2910 16836 2966 16892
rect 2966 16836 2970 16892
rect 2906 16832 2970 16836
rect 2986 16892 3050 16896
rect 2986 16836 2990 16892
rect 2990 16836 3046 16892
rect 3046 16836 3050 16892
rect 2986 16832 3050 16836
rect 3066 16892 3130 16896
rect 3066 16836 3070 16892
rect 3070 16836 3126 16892
rect 3126 16836 3130 16892
rect 3066 16832 3130 16836
rect 6574 16892 6638 16896
rect 6574 16836 6578 16892
rect 6578 16836 6634 16892
rect 6634 16836 6638 16892
rect 6574 16832 6638 16836
rect 6654 16892 6718 16896
rect 6654 16836 6658 16892
rect 6658 16836 6714 16892
rect 6714 16836 6718 16892
rect 6654 16832 6718 16836
rect 6734 16892 6798 16896
rect 6734 16836 6738 16892
rect 6738 16836 6794 16892
rect 6794 16836 6798 16892
rect 6734 16832 6798 16836
rect 6814 16892 6878 16896
rect 6814 16836 6818 16892
rect 6818 16836 6874 16892
rect 6874 16836 6878 16892
rect 6814 16832 6878 16836
rect 10322 16892 10386 16896
rect 10322 16836 10326 16892
rect 10326 16836 10382 16892
rect 10382 16836 10386 16892
rect 10322 16832 10386 16836
rect 10402 16892 10466 16896
rect 10402 16836 10406 16892
rect 10406 16836 10462 16892
rect 10462 16836 10466 16892
rect 10402 16832 10466 16836
rect 10482 16892 10546 16896
rect 10482 16836 10486 16892
rect 10486 16836 10542 16892
rect 10542 16836 10546 16892
rect 10482 16832 10546 16836
rect 10562 16892 10626 16896
rect 10562 16836 10566 16892
rect 10566 16836 10622 16892
rect 10622 16836 10626 16892
rect 10562 16832 10626 16836
rect 14070 16892 14134 16896
rect 14070 16836 14074 16892
rect 14074 16836 14130 16892
rect 14130 16836 14134 16892
rect 14070 16832 14134 16836
rect 14150 16892 14214 16896
rect 14150 16836 14154 16892
rect 14154 16836 14210 16892
rect 14210 16836 14214 16892
rect 14150 16832 14214 16836
rect 14230 16892 14294 16896
rect 14230 16836 14234 16892
rect 14234 16836 14290 16892
rect 14290 16836 14294 16892
rect 14230 16832 14294 16836
rect 14310 16892 14374 16896
rect 14310 16836 14314 16892
rect 14314 16836 14370 16892
rect 14370 16836 14374 16892
rect 14310 16832 14374 16836
rect 4700 16348 4764 16352
rect 4700 16292 4704 16348
rect 4704 16292 4760 16348
rect 4760 16292 4764 16348
rect 4700 16288 4764 16292
rect 4780 16348 4844 16352
rect 4780 16292 4784 16348
rect 4784 16292 4840 16348
rect 4840 16292 4844 16348
rect 4780 16288 4844 16292
rect 4860 16348 4924 16352
rect 4860 16292 4864 16348
rect 4864 16292 4920 16348
rect 4920 16292 4924 16348
rect 4860 16288 4924 16292
rect 4940 16348 5004 16352
rect 4940 16292 4944 16348
rect 4944 16292 5000 16348
rect 5000 16292 5004 16348
rect 4940 16288 5004 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 12196 16348 12260 16352
rect 12196 16292 12200 16348
rect 12200 16292 12256 16348
rect 12256 16292 12260 16348
rect 12196 16288 12260 16292
rect 12276 16348 12340 16352
rect 12276 16292 12280 16348
rect 12280 16292 12336 16348
rect 12336 16292 12340 16348
rect 12276 16288 12340 16292
rect 12356 16348 12420 16352
rect 12356 16292 12360 16348
rect 12360 16292 12416 16348
rect 12416 16292 12420 16348
rect 12356 16288 12420 16292
rect 12436 16348 12500 16352
rect 12436 16292 12440 16348
rect 12440 16292 12496 16348
rect 12496 16292 12500 16348
rect 12436 16288 12500 16292
rect 2826 15804 2890 15808
rect 2826 15748 2830 15804
rect 2830 15748 2886 15804
rect 2886 15748 2890 15804
rect 2826 15744 2890 15748
rect 2906 15804 2970 15808
rect 2906 15748 2910 15804
rect 2910 15748 2966 15804
rect 2966 15748 2970 15804
rect 2906 15744 2970 15748
rect 2986 15804 3050 15808
rect 2986 15748 2990 15804
rect 2990 15748 3046 15804
rect 3046 15748 3050 15804
rect 2986 15744 3050 15748
rect 3066 15804 3130 15808
rect 3066 15748 3070 15804
rect 3070 15748 3126 15804
rect 3126 15748 3130 15804
rect 3066 15744 3130 15748
rect 6574 15804 6638 15808
rect 6574 15748 6578 15804
rect 6578 15748 6634 15804
rect 6634 15748 6638 15804
rect 6574 15744 6638 15748
rect 6654 15804 6718 15808
rect 6654 15748 6658 15804
rect 6658 15748 6714 15804
rect 6714 15748 6718 15804
rect 6654 15744 6718 15748
rect 6734 15804 6798 15808
rect 6734 15748 6738 15804
rect 6738 15748 6794 15804
rect 6794 15748 6798 15804
rect 6734 15744 6798 15748
rect 6814 15804 6878 15808
rect 6814 15748 6818 15804
rect 6818 15748 6874 15804
rect 6874 15748 6878 15804
rect 6814 15744 6878 15748
rect 10322 15804 10386 15808
rect 10322 15748 10326 15804
rect 10326 15748 10382 15804
rect 10382 15748 10386 15804
rect 10322 15744 10386 15748
rect 10402 15804 10466 15808
rect 10402 15748 10406 15804
rect 10406 15748 10462 15804
rect 10462 15748 10466 15804
rect 10402 15744 10466 15748
rect 10482 15804 10546 15808
rect 10482 15748 10486 15804
rect 10486 15748 10542 15804
rect 10542 15748 10546 15804
rect 10482 15744 10546 15748
rect 10562 15804 10626 15808
rect 10562 15748 10566 15804
rect 10566 15748 10622 15804
rect 10622 15748 10626 15804
rect 10562 15744 10626 15748
rect 14070 15804 14134 15808
rect 14070 15748 14074 15804
rect 14074 15748 14130 15804
rect 14130 15748 14134 15804
rect 14070 15744 14134 15748
rect 14150 15804 14214 15808
rect 14150 15748 14154 15804
rect 14154 15748 14210 15804
rect 14210 15748 14214 15804
rect 14150 15744 14214 15748
rect 14230 15804 14294 15808
rect 14230 15748 14234 15804
rect 14234 15748 14290 15804
rect 14290 15748 14294 15804
rect 14230 15744 14294 15748
rect 14310 15804 14374 15808
rect 14310 15748 14314 15804
rect 14314 15748 14370 15804
rect 14370 15748 14374 15804
rect 14310 15744 14374 15748
rect 4700 15260 4764 15264
rect 4700 15204 4704 15260
rect 4704 15204 4760 15260
rect 4760 15204 4764 15260
rect 4700 15200 4764 15204
rect 4780 15260 4844 15264
rect 4780 15204 4784 15260
rect 4784 15204 4840 15260
rect 4840 15204 4844 15260
rect 4780 15200 4844 15204
rect 4860 15260 4924 15264
rect 4860 15204 4864 15260
rect 4864 15204 4920 15260
rect 4920 15204 4924 15260
rect 4860 15200 4924 15204
rect 4940 15260 5004 15264
rect 4940 15204 4944 15260
rect 4944 15204 5000 15260
rect 5000 15204 5004 15260
rect 4940 15200 5004 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 12196 15260 12260 15264
rect 12196 15204 12200 15260
rect 12200 15204 12256 15260
rect 12256 15204 12260 15260
rect 12196 15200 12260 15204
rect 12276 15260 12340 15264
rect 12276 15204 12280 15260
rect 12280 15204 12336 15260
rect 12336 15204 12340 15260
rect 12276 15200 12340 15204
rect 12356 15260 12420 15264
rect 12356 15204 12360 15260
rect 12360 15204 12416 15260
rect 12416 15204 12420 15260
rect 12356 15200 12420 15204
rect 12436 15260 12500 15264
rect 12436 15204 12440 15260
rect 12440 15204 12496 15260
rect 12496 15204 12500 15260
rect 12436 15200 12500 15204
rect 2826 14716 2890 14720
rect 2826 14660 2830 14716
rect 2830 14660 2886 14716
rect 2886 14660 2890 14716
rect 2826 14656 2890 14660
rect 2906 14716 2970 14720
rect 2906 14660 2910 14716
rect 2910 14660 2966 14716
rect 2966 14660 2970 14716
rect 2906 14656 2970 14660
rect 2986 14716 3050 14720
rect 2986 14660 2990 14716
rect 2990 14660 3046 14716
rect 3046 14660 3050 14716
rect 2986 14656 3050 14660
rect 3066 14716 3130 14720
rect 3066 14660 3070 14716
rect 3070 14660 3126 14716
rect 3126 14660 3130 14716
rect 3066 14656 3130 14660
rect 6574 14716 6638 14720
rect 6574 14660 6578 14716
rect 6578 14660 6634 14716
rect 6634 14660 6638 14716
rect 6574 14656 6638 14660
rect 6654 14716 6718 14720
rect 6654 14660 6658 14716
rect 6658 14660 6714 14716
rect 6714 14660 6718 14716
rect 6654 14656 6718 14660
rect 6734 14716 6798 14720
rect 6734 14660 6738 14716
rect 6738 14660 6794 14716
rect 6794 14660 6798 14716
rect 6734 14656 6798 14660
rect 6814 14716 6878 14720
rect 6814 14660 6818 14716
rect 6818 14660 6874 14716
rect 6874 14660 6878 14716
rect 6814 14656 6878 14660
rect 10322 14716 10386 14720
rect 10322 14660 10326 14716
rect 10326 14660 10382 14716
rect 10382 14660 10386 14716
rect 10322 14656 10386 14660
rect 10402 14716 10466 14720
rect 10402 14660 10406 14716
rect 10406 14660 10462 14716
rect 10462 14660 10466 14716
rect 10402 14656 10466 14660
rect 10482 14716 10546 14720
rect 10482 14660 10486 14716
rect 10486 14660 10542 14716
rect 10542 14660 10546 14716
rect 10482 14656 10546 14660
rect 10562 14716 10626 14720
rect 10562 14660 10566 14716
rect 10566 14660 10622 14716
rect 10622 14660 10626 14716
rect 10562 14656 10626 14660
rect 14070 14716 14134 14720
rect 14070 14660 14074 14716
rect 14074 14660 14130 14716
rect 14130 14660 14134 14716
rect 14070 14656 14134 14660
rect 14150 14716 14214 14720
rect 14150 14660 14154 14716
rect 14154 14660 14210 14716
rect 14210 14660 14214 14716
rect 14150 14656 14214 14660
rect 14230 14716 14294 14720
rect 14230 14660 14234 14716
rect 14234 14660 14290 14716
rect 14290 14660 14294 14716
rect 14230 14656 14294 14660
rect 14310 14716 14374 14720
rect 14310 14660 14314 14716
rect 14314 14660 14370 14716
rect 14370 14660 14374 14716
rect 14310 14656 14374 14660
rect 4700 14172 4764 14176
rect 4700 14116 4704 14172
rect 4704 14116 4760 14172
rect 4760 14116 4764 14172
rect 4700 14112 4764 14116
rect 4780 14172 4844 14176
rect 4780 14116 4784 14172
rect 4784 14116 4840 14172
rect 4840 14116 4844 14172
rect 4780 14112 4844 14116
rect 4860 14172 4924 14176
rect 4860 14116 4864 14172
rect 4864 14116 4920 14172
rect 4920 14116 4924 14172
rect 4860 14112 4924 14116
rect 4940 14172 5004 14176
rect 4940 14116 4944 14172
rect 4944 14116 5000 14172
rect 5000 14116 5004 14172
rect 4940 14112 5004 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 12196 14172 12260 14176
rect 12196 14116 12200 14172
rect 12200 14116 12256 14172
rect 12256 14116 12260 14172
rect 12196 14112 12260 14116
rect 12276 14172 12340 14176
rect 12276 14116 12280 14172
rect 12280 14116 12336 14172
rect 12336 14116 12340 14172
rect 12276 14112 12340 14116
rect 12356 14172 12420 14176
rect 12356 14116 12360 14172
rect 12360 14116 12416 14172
rect 12416 14116 12420 14172
rect 12356 14112 12420 14116
rect 12436 14172 12500 14176
rect 12436 14116 12440 14172
rect 12440 14116 12496 14172
rect 12496 14116 12500 14172
rect 12436 14112 12500 14116
rect 2826 13628 2890 13632
rect 2826 13572 2830 13628
rect 2830 13572 2886 13628
rect 2886 13572 2890 13628
rect 2826 13568 2890 13572
rect 2906 13628 2970 13632
rect 2906 13572 2910 13628
rect 2910 13572 2966 13628
rect 2966 13572 2970 13628
rect 2906 13568 2970 13572
rect 2986 13628 3050 13632
rect 2986 13572 2990 13628
rect 2990 13572 3046 13628
rect 3046 13572 3050 13628
rect 2986 13568 3050 13572
rect 3066 13628 3130 13632
rect 3066 13572 3070 13628
rect 3070 13572 3126 13628
rect 3126 13572 3130 13628
rect 3066 13568 3130 13572
rect 6574 13628 6638 13632
rect 6574 13572 6578 13628
rect 6578 13572 6634 13628
rect 6634 13572 6638 13628
rect 6574 13568 6638 13572
rect 6654 13628 6718 13632
rect 6654 13572 6658 13628
rect 6658 13572 6714 13628
rect 6714 13572 6718 13628
rect 6654 13568 6718 13572
rect 6734 13628 6798 13632
rect 6734 13572 6738 13628
rect 6738 13572 6794 13628
rect 6794 13572 6798 13628
rect 6734 13568 6798 13572
rect 6814 13628 6878 13632
rect 6814 13572 6818 13628
rect 6818 13572 6874 13628
rect 6874 13572 6878 13628
rect 6814 13568 6878 13572
rect 10322 13628 10386 13632
rect 10322 13572 10326 13628
rect 10326 13572 10382 13628
rect 10382 13572 10386 13628
rect 10322 13568 10386 13572
rect 10402 13628 10466 13632
rect 10402 13572 10406 13628
rect 10406 13572 10462 13628
rect 10462 13572 10466 13628
rect 10402 13568 10466 13572
rect 10482 13628 10546 13632
rect 10482 13572 10486 13628
rect 10486 13572 10542 13628
rect 10542 13572 10546 13628
rect 10482 13568 10546 13572
rect 10562 13628 10626 13632
rect 10562 13572 10566 13628
rect 10566 13572 10622 13628
rect 10622 13572 10626 13628
rect 10562 13568 10626 13572
rect 14070 13628 14134 13632
rect 14070 13572 14074 13628
rect 14074 13572 14130 13628
rect 14130 13572 14134 13628
rect 14070 13568 14134 13572
rect 14150 13628 14214 13632
rect 14150 13572 14154 13628
rect 14154 13572 14210 13628
rect 14210 13572 14214 13628
rect 14150 13568 14214 13572
rect 14230 13628 14294 13632
rect 14230 13572 14234 13628
rect 14234 13572 14290 13628
rect 14290 13572 14294 13628
rect 14230 13568 14294 13572
rect 14310 13628 14374 13632
rect 14310 13572 14314 13628
rect 14314 13572 14370 13628
rect 14370 13572 14374 13628
rect 14310 13568 14374 13572
rect 4700 13084 4764 13088
rect 4700 13028 4704 13084
rect 4704 13028 4760 13084
rect 4760 13028 4764 13084
rect 4700 13024 4764 13028
rect 4780 13084 4844 13088
rect 4780 13028 4784 13084
rect 4784 13028 4840 13084
rect 4840 13028 4844 13084
rect 4780 13024 4844 13028
rect 4860 13084 4924 13088
rect 4860 13028 4864 13084
rect 4864 13028 4920 13084
rect 4920 13028 4924 13084
rect 4860 13024 4924 13028
rect 4940 13084 5004 13088
rect 4940 13028 4944 13084
rect 4944 13028 5000 13084
rect 5000 13028 5004 13084
rect 4940 13024 5004 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 12196 13084 12260 13088
rect 12196 13028 12200 13084
rect 12200 13028 12256 13084
rect 12256 13028 12260 13084
rect 12196 13024 12260 13028
rect 12276 13084 12340 13088
rect 12276 13028 12280 13084
rect 12280 13028 12336 13084
rect 12336 13028 12340 13084
rect 12276 13024 12340 13028
rect 12356 13084 12420 13088
rect 12356 13028 12360 13084
rect 12360 13028 12416 13084
rect 12416 13028 12420 13084
rect 12356 13024 12420 13028
rect 12436 13084 12500 13088
rect 12436 13028 12440 13084
rect 12440 13028 12496 13084
rect 12496 13028 12500 13084
rect 12436 13024 12500 13028
rect 2826 12540 2890 12544
rect 2826 12484 2830 12540
rect 2830 12484 2886 12540
rect 2886 12484 2890 12540
rect 2826 12480 2890 12484
rect 2906 12540 2970 12544
rect 2906 12484 2910 12540
rect 2910 12484 2966 12540
rect 2966 12484 2970 12540
rect 2906 12480 2970 12484
rect 2986 12540 3050 12544
rect 2986 12484 2990 12540
rect 2990 12484 3046 12540
rect 3046 12484 3050 12540
rect 2986 12480 3050 12484
rect 3066 12540 3130 12544
rect 3066 12484 3070 12540
rect 3070 12484 3126 12540
rect 3126 12484 3130 12540
rect 3066 12480 3130 12484
rect 6574 12540 6638 12544
rect 6574 12484 6578 12540
rect 6578 12484 6634 12540
rect 6634 12484 6638 12540
rect 6574 12480 6638 12484
rect 6654 12540 6718 12544
rect 6654 12484 6658 12540
rect 6658 12484 6714 12540
rect 6714 12484 6718 12540
rect 6654 12480 6718 12484
rect 6734 12540 6798 12544
rect 6734 12484 6738 12540
rect 6738 12484 6794 12540
rect 6794 12484 6798 12540
rect 6734 12480 6798 12484
rect 6814 12540 6878 12544
rect 6814 12484 6818 12540
rect 6818 12484 6874 12540
rect 6874 12484 6878 12540
rect 6814 12480 6878 12484
rect 10322 12540 10386 12544
rect 10322 12484 10326 12540
rect 10326 12484 10382 12540
rect 10382 12484 10386 12540
rect 10322 12480 10386 12484
rect 10402 12540 10466 12544
rect 10402 12484 10406 12540
rect 10406 12484 10462 12540
rect 10462 12484 10466 12540
rect 10402 12480 10466 12484
rect 10482 12540 10546 12544
rect 10482 12484 10486 12540
rect 10486 12484 10542 12540
rect 10542 12484 10546 12540
rect 10482 12480 10546 12484
rect 10562 12540 10626 12544
rect 10562 12484 10566 12540
rect 10566 12484 10622 12540
rect 10622 12484 10626 12540
rect 10562 12480 10626 12484
rect 14070 12540 14134 12544
rect 14070 12484 14074 12540
rect 14074 12484 14130 12540
rect 14130 12484 14134 12540
rect 14070 12480 14134 12484
rect 14150 12540 14214 12544
rect 14150 12484 14154 12540
rect 14154 12484 14210 12540
rect 14210 12484 14214 12540
rect 14150 12480 14214 12484
rect 14230 12540 14294 12544
rect 14230 12484 14234 12540
rect 14234 12484 14290 12540
rect 14290 12484 14294 12540
rect 14230 12480 14294 12484
rect 14310 12540 14374 12544
rect 14310 12484 14314 12540
rect 14314 12484 14370 12540
rect 14370 12484 14374 12540
rect 14310 12480 14374 12484
rect 4700 11996 4764 12000
rect 4700 11940 4704 11996
rect 4704 11940 4760 11996
rect 4760 11940 4764 11996
rect 4700 11936 4764 11940
rect 4780 11996 4844 12000
rect 4780 11940 4784 11996
rect 4784 11940 4840 11996
rect 4840 11940 4844 11996
rect 4780 11936 4844 11940
rect 4860 11996 4924 12000
rect 4860 11940 4864 11996
rect 4864 11940 4920 11996
rect 4920 11940 4924 11996
rect 4860 11936 4924 11940
rect 4940 11996 5004 12000
rect 4940 11940 4944 11996
rect 4944 11940 5000 11996
rect 5000 11940 5004 11996
rect 4940 11936 5004 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 12196 11996 12260 12000
rect 12196 11940 12200 11996
rect 12200 11940 12256 11996
rect 12256 11940 12260 11996
rect 12196 11936 12260 11940
rect 12276 11996 12340 12000
rect 12276 11940 12280 11996
rect 12280 11940 12336 11996
rect 12336 11940 12340 11996
rect 12276 11936 12340 11940
rect 12356 11996 12420 12000
rect 12356 11940 12360 11996
rect 12360 11940 12416 11996
rect 12416 11940 12420 11996
rect 12356 11936 12420 11940
rect 12436 11996 12500 12000
rect 12436 11940 12440 11996
rect 12440 11940 12496 11996
rect 12496 11940 12500 11996
rect 12436 11936 12500 11940
rect 2826 11452 2890 11456
rect 2826 11396 2830 11452
rect 2830 11396 2886 11452
rect 2886 11396 2890 11452
rect 2826 11392 2890 11396
rect 2906 11452 2970 11456
rect 2906 11396 2910 11452
rect 2910 11396 2966 11452
rect 2966 11396 2970 11452
rect 2906 11392 2970 11396
rect 2986 11452 3050 11456
rect 2986 11396 2990 11452
rect 2990 11396 3046 11452
rect 3046 11396 3050 11452
rect 2986 11392 3050 11396
rect 3066 11452 3130 11456
rect 3066 11396 3070 11452
rect 3070 11396 3126 11452
rect 3126 11396 3130 11452
rect 3066 11392 3130 11396
rect 6574 11452 6638 11456
rect 6574 11396 6578 11452
rect 6578 11396 6634 11452
rect 6634 11396 6638 11452
rect 6574 11392 6638 11396
rect 6654 11452 6718 11456
rect 6654 11396 6658 11452
rect 6658 11396 6714 11452
rect 6714 11396 6718 11452
rect 6654 11392 6718 11396
rect 6734 11452 6798 11456
rect 6734 11396 6738 11452
rect 6738 11396 6794 11452
rect 6794 11396 6798 11452
rect 6734 11392 6798 11396
rect 6814 11452 6878 11456
rect 6814 11396 6818 11452
rect 6818 11396 6874 11452
rect 6874 11396 6878 11452
rect 6814 11392 6878 11396
rect 10322 11452 10386 11456
rect 10322 11396 10326 11452
rect 10326 11396 10382 11452
rect 10382 11396 10386 11452
rect 10322 11392 10386 11396
rect 10402 11452 10466 11456
rect 10402 11396 10406 11452
rect 10406 11396 10462 11452
rect 10462 11396 10466 11452
rect 10402 11392 10466 11396
rect 10482 11452 10546 11456
rect 10482 11396 10486 11452
rect 10486 11396 10542 11452
rect 10542 11396 10546 11452
rect 10482 11392 10546 11396
rect 10562 11452 10626 11456
rect 10562 11396 10566 11452
rect 10566 11396 10622 11452
rect 10622 11396 10626 11452
rect 10562 11392 10626 11396
rect 14070 11452 14134 11456
rect 14070 11396 14074 11452
rect 14074 11396 14130 11452
rect 14130 11396 14134 11452
rect 14070 11392 14134 11396
rect 14150 11452 14214 11456
rect 14150 11396 14154 11452
rect 14154 11396 14210 11452
rect 14210 11396 14214 11452
rect 14150 11392 14214 11396
rect 14230 11452 14294 11456
rect 14230 11396 14234 11452
rect 14234 11396 14290 11452
rect 14290 11396 14294 11452
rect 14230 11392 14294 11396
rect 14310 11452 14374 11456
rect 14310 11396 14314 11452
rect 14314 11396 14370 11452
rect 14370 11396 14374 11452
rect 14310 11392 14374 11396
rect 8892 11188 8956 11252
rect 4700 10908 4764 10912
rect 4700 10852 4704 10908
rect 4704 10852 4760 10908
rect 4760 10852 4764 10908
rect 4700 10848 4764 10852
rect 4780 10908 4844 10912
rect 4780 10852 4784 10908
rect 4784 10852 4840 10908
rect 4840 10852 4844 10908
rect 4780 10848 4844 10852
rect 4860 10908 4924 10912
rect 4860 10852 4864 10908
rect 4864 10852 4920 10908
rect 4920 10852 4924 10908
rect 4860 10848 4924 10852
rect 4940 10908 5004 10912
rect 4940 10852 4944 10908
rect 4944 10852 5000 10908
rect 5000 10852 5004 10908
rect 4940 10848 5004 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 12196 10908 12260 10912
rect 12196 10852 12200 10908
rect 12200 10852 12256 10908
rect 12256 10852 12260 10908
rect 12196 10848 12260 10852
rect 12276 10908 12340 10912
rect 12276 10852 12280 10908
rect 12280 10852 12336 10908
rect 12336 10852 12340 10908
rect 12276 10848 12340 10852
rect 12356 10908 12420 10912
rect 12356 10852 12360 10908
rect 12360 10852 12416 10908
rect 12416 10852 12420 10908
rect 12356 10848 12420 10852
rect 12436 10908 12500 10912
rect 12436 10852 12440 10908
rect 12440 10852 12496 10908
rect 12496 10852 12500 10908
rect 12436 10848 12500 10852
rect 2826 10364 2890 10368
rect 2826 10308 2830 10364
rect 2830 10308 2886 10364
rect 2886 10308 2890 10364
rect 2826 10304 2890 10308
rect 2906 10364 2970 10368
rect 2906 10308 2910 10364
rect 2910 10308 2966 10364
rect 2966 10308 2970 10364
rect 2906 10304 2970 10308
rect 2986 10364 3050 10368
rect 2986 10308 2990 10364
rect 2990 10308 3046 10364
rect 3046 10308 3050 10364
rect 2986 10304 3050 10308
rect 3066 10364 3130 10368
rect 3066 10308 3070 10364
rect 3070 10308 3126 10364
rect 3126 10308 3130 10364
rect 3066 10304 3130 10308
rect 6574 10364 6638 10368
rect 6574 10308 6578 10364
rect 6578 10308 6634 10364
rect 6634 10308 6638 10364
rect 6574 10304 6638 10308
rect 6654 10364 6718 10368
rect 6654 10308 6658 10364
rect 6658 10308 6714 10364
rect 6714 10308 6718 10364
rect 6654 10304 6718 10308
rect 6734 10364 6798 10368
rect 6734 10308 6738 10364
rect 6738 10308 6794 10364
rect 6794 10308 6798 10364
rect 6734 10304 6798 10308
rect 6814 10364 6878 10368
rect 6814 10308 6818 10364
rect 6818 10308 6874 10364
rect 6874 10308 6878 10364
rect 6814 10304 6878 10308
rect 10322 10364 10386 10368
rect 10322 10308 10326 10364
rect 10326 10308 10382 10364
rect 10382 10308 10386 10364
rect 10322 10304 10386 10308
rect 10402 10364 10466 10368
rect 10402 10308 10406 10364
rect 10406 10308 10462 10364
rect 10462 10308 10466 10364
rect 10402 10304 10466 10308
rect 10482 10364 10546 10368
rect 10482 10308 10486 10364
rect 10486 10308 10542 10364
rect 10542 10308 10546 10364
rect 10482 10304 10546 10308
rect 10562 10364 10626 10368
rect 10562 10308 10566 10364
rect 10566 10308 10622 10364
rect 10622 10308 10626 10364
rect 10562 10304 10626 10308
rect 14070 10364 14134 10368
rect 14070 10308 14074 10364
rect 14074 10308 14130 10364
rect 14130 10308 14134 10364
rect 14070 10304 14134 10308
rect 14150 10364 14214 10368
rect 14150 10308 14154 10364
rect 14154 10308 14210 10364
rect 14210 10308 14214 10364
rect 14150 10304 14214 10308
rect 14230 10364 14294 10368
rect 14230 10308 14234 10364
rect 14234 10308 14290 10364
rect 14290 10308 14294 10364
rect 14230 10304 14294 10308
rect 14310 10364 14374 10368
rect 14310 10308 14314 10364
rect 14314 10308 14370 10364
rect 14370 10308 14374 10364
rect 14310 10304 14374 10308
rect 4700 9820 4764 9824
rect 4700 9764 4704 9820
rect 4704 9764 4760 9820
rect 4760 9764 4764 9820
rect 4700 9760 4764 9764
rect 4780 9820 4844 9824
rect 4780 9764 4784 9820
rect 4784 9764 4840 9820
rect 4840 9764 4844 9820
rect 4780 9760 4844 9764
rect 4860 9820 4924 9824
rect 4860 9764 4864 9820
rect 4864 9764 4920 9820
rect 4920 9764 4924 9820
rect 4860 9760 4924 9764
rect 4940 9820 5004 9824
rect 4940 9764 4944 9820
rect 4944 9764 5000 9820
rect 5000 9764 5004 9820
rect 4940 9760 5004 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 12196 9820 12260 9824
rect 12196 9764 12200 9820
rect 12200 9764 12256 9820
rect 12256 9764 12260 9820
rect 12196 9760 12260 9764
rect 12276 9820 12340 9824
rect 12276 9764 12280 9820
rect 12280 9764 12336 9820
rect 12336 9764 12340 9820
rect 12276 9760 12340 9764
rect 12356 9820 12420 9824
rect 12356 9764 12360 9820
rect 12360 9764 12416 9820
rect 12416 9764 12420 9820
rect 12356 9760 12420 9764
rect 12436 9820 12500 9824
rect 12436 9764 12440 9820
rect 12440 9764 12496 9820
rect 12496 9764 12500 9820
rect 12436 9760 12500 9764
rect 8892 9752 8956 9756
rect 8892 9696 8906 9752
rect 8906 9696 8956 9752
rect 8892 9692 8956 9696
rect 2826 9276 2890 9280
rect 2826 9220 2830 9276
rect 2830 9220 2886 9276
rect 2886 9220 2890 9276
rect 2826 9216 2890 9220
rect 2906 9276 2970 9280
rect 2906 9220 2910 9276
rect 2910 9220 2966 9276
rect 2966 9220 2970 9276
rect 2906 9216 2970 9220
rect 2986 9276 3050 9280
rect 2986 9220 2990 9276
rect 2990 9220 3046 9276
rect 3046 9220 3050 9276
rect 2986 9216 3050 9220
rect 3066 9276 3130 9280
rect 3066 9220 3070 9276
rect 3070 9220 3126 9276
rect 3126 9220 3130 9276
rect 3066 9216 3130 9220
rect 6574 9276 6638 9280
rect 6574 9220 6578 9276
rect 6578 9220 6634 9276
rect 6634 9220 6638 9276
rect 6574 9216 6638 9220
rect 6654 9276 6718 9280
rect 6654 9220 6658 9276
rect 6658 9220 6714 9276
rect 6714 9220 6718 9276
rect 6654 9216 6718 9220
rect 6734 9276 6798 9280
rect 6734 9220 6738 9276
rect 6738 9220 6794 9276
rect 6794 9220 6798 9276
rect 6734 9216 6798 9220
rect 6814 9276 6878 9280
rect 6814 9220 6818 9276
rect 6818 9220 6874 9276
rect 6874 9220 6878 9276
rect 6814 9216 6878 9220
rect 10322 9276 10386 9280
rect 10322 9220 10326 9276
rect 10326 9220 10382 9276
rect 10382 9220 10386 9276
rect 10322 9216 10386 9220
rect 10402 9276 10466 9280
rect 10402 9220 10406 9276
rect 10406 9220 10462 9276
rect 10462 9220 10466 9276
rect 10402 9216 10466 9220
rect 10482 9276 10546 9280
rect 10482 9220 10486 9276
rect 10486 9220 10542 9276
rect 10542 9220 10546 9276
rect 10482 9216 10546 9220
rect 10562 9276 10626 9280
rect 10562 9220 10566 9276
rect 10566 9220 10622 9276
rect 10622 9220 10626 9276
rect 10562 9216 10626 9220
rect 14070 9276 14134 9280
rect 14070 9220 14074 9276
rect 14074 9220 14130 9276
rect 14130 9220 14134 9276
rect 14070 9216 14134 9220
rect 14150 9276 14214 9280
rect 14150 9220 14154 9276
rect 14154 9220 14210 9276
rect 14210 9220 14214 9276
rect 14150 9216 14214 9220
rect 14230 9276 14294 9280
rect 14230 9220 14234 9276
rect 14234 9220 14290 9276
rect 14290 9220 14294 9276
rect 14230 9216 14294 9220
rect 14310 9276 14374 9280
rect 14310 9220 14314 9276
rect 14314 9220 14370 9276
rect 14370 9220 14374 9276
rect 14310 9216 14374 9220
rect 4700 8732 4764 8736
rect 4700 8676 4704 8732
rect 4704 8676 4760 8732
rect 4760 8676 4764 8732
rect 4700 8672 4764 8676
rect 4780 8732 4844 8736
rect 4780 8676 4784 8732
rect 4784 8676 4840 8732
rect 4840 8676 4844 8732
rect 4780 8672 4844 8676
rect 4860 8732 4924 8736
rect 4860 8676 4864 8732
rect 4864 8676 4920 8732
rect 4920 8676 4924 8732
rect 4860 8672 4924 8676
rect 4940 8732 5004 8736
rect 4940 8676 4944 8732
rect 4944 8676 5000 8732
rect 5000 8676 5004 8732
rect 4940 8672 5004 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 12196 8732 12260 8736
rect 12196 8676 12200 8732
rect 12200 8676 12256 8732
rect 12256 8676 12260 8732
rect 12196 8672 12260 8676
rect 12276 8732 12340 8736
rect 12276 8676 12280 8732
rect 12280 8676 12336 8732
rect 12336 8676 12340 8732
rect 12276 8672 12340 8676
rect 12356 8732 12420 8736
rect 12356 8676 12360 8732
rect 12360 8676 12416 8732
rect 12416 8676 12420 8732
rect 12356 8672 12420 8676
rect 12436 8732 12500 8736
rect 12436 8676 12440 8732
rect 12440 8676 12496 8732
rect 12496 8676 12500 8732
rect 12436 8672 12500 8676
rect 2826 8188 2890 8192
rect 2826 8132 2830 8188
rect 2830 8132 2886 8188
rect 2886 8132 2890 8188
rect 2826 8128 2890 8132
rect 2906 8188 2970 8192
rect 2906 8132 2910 8188
rect 2910 8132 2966 8188
rect 2966 8132 2970 8188
rect 2906 8128 2970 8132
rect 2986 8188 3050 8192
rect 2986 8132 2990 8188
rect 2990 8132 3046 8188
rect 3046 8132 3050 8188
rect 2986 8128 3050 8132
rect 3066 8188 3130 8192
rect 3066 8132 3070 8188
rect 3070 8132 3126 8188
rect 3126 8132 3130 8188
rect 3066 8128 3130 8132
rect 6574 8188 6638 8192
rect 6574 8132 6578 8188
rect 6578 8132 6634 8188
rect 6634 8132 6638 8188
rect 6574 8128 6638 8132
rect 6654 8188 6718 8192
rect 6654 8132 6658 8188
rect 6658 8132 6714 8188
rect 6714 8132 6718 8188
rect 6654 8128 6718 8132
rect 6734 8188 6798 8192
rect 6734 8132 6738 8188
rect 6738 8132 6794 8188
rect 6794 8132 6798 8188
rect 6734 8128 6798 8132
rect 6814 8188 6878 8192
rect 6814 8132 6818 8188
rect 6818 8132 6874 8188
rect 6874 8132 6878 8188
rect 6814 8128 6878 8132
rect 10322 8188 10386 8192
rect 10322 8132 10326 8188
rect 10326 8132 10382 8188
rect 10382 8132 10386 8188
rect 10322 8128 10386 8132
rect 10402 8188 10466 8192
rect 10402 8132 10406 8188
rect 10406 8132 10462 8188
rect 10462 8132 10466 8188
rect 10402 8128 10466 8132
rect 10482 8188 10546 8192
rect 10482 8132 10486 8188
rect 10486 8132 10542 8188
rect 10542 8132 10546 8188
rect 10482 8128 10546 8132
rect 10562 8188 10626 8192
rect 10562 8132 10566 8188
rect 10566 8132 10622 8188
rect 10622 8132 10626 8188
rect 10562 8128 10626 8132
rect 14070 8188 14134 8192
rect 14070 8132 14074 8188
rect 14074 8132 14130 8188
rect 14130 8132 14134 8188
rect 14070 8128 14134 8132
rect 14150 8188 14214 8192
rect 14150 8132 14154 8188
rect 14154 8132 14210 8188
rect 14210 8132 14214 8188
rect 14150 8128 14214 8132
rect 14230 8188 14294 8192
rect 14230 8132 14234 8188
rect 14234 8132 14290 8188
rect 14290 8132 14294 8188
rect 14230 8128 14294 8132
rect 14310 8188 14374 8192
rect 14310 8132 14314 8188
rect 14314 8132 14370 8188
rect 14370 8132 14374 8188
rect 14310 8128 14374 8132
rect 4700 7644 4764 7648
rect 4700 7588 4704 7644
rect 4704 7588 4760 7644
rect 4760 7588 4764 7644
rect 4700 7584 4764 7588
rect 4780 7644 4844 7648
rect 4780 7588 4784 7644
rect 4784 7588 4840 7644
rect 4840 7588 4844 7644
rect 4780 7584 4844 7588
rect 4860 7644 4924 7648
rect 4860 7588 4864 7644
rect 4864 7588 4920 7644
rect 4920 7588 4924 7644
rect 4860 7584 4924 7588
rect 4940 7644 5004 7648
rect 4940 7588 4944 7644
rect 4944 7588 5000 7644
rect 5000 7588 5004 7644
rect 4940 7584 5004 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 12196 7644 12260 7648
rect 12196 7588 12200 7644
rect 12200 7588 12256 7644
rect 12256 7588 12260 7644
rect 12196 7584 12260 7588
rect 12276 7644 12340 7648
rect 12276 7588 12280 7644
rect 12280 7588 12336 7644
rect 12336 7588 12340 7644
rect 12276 7584 12340 7588
rect 12356 7644 12420 7648
rect 12356 7588 12360 7644
rect 12360 7588 12416 7644
rect 12416 7588 12420 7644
rect 12356 7584 12420 7588
rect 12436 7644 12500 7648
rect 12436 7588 12440 7644
rect 12440 7588 12496 7644
rect 12496 7588 12500 7644
rect 12436 7584 12500 7588
rect 2826 7100 2890 7104
rect 2826 7044 2830 7100
rect 2830 7044 2886 7100
rect 2886 7044 2890 7100
rect 2826 7040 2890 7044
rect 2906 7100 2970 7104
rect 2906 7044 2910 7100
rect 2910 7044 2966 7100
rect 2966 7044 2970 7100
rect 2906 7040 2970 7044
rect 2986 7100 3050 7104
rect 2986 7044 2990 7100
rect 2990 7044 3046 7100
rect 3046 7044 3050 7100
rect 2986 7040 3050 7044
rect 3066 7100 3130 7104
rect 3066 7044 3070 7100
rect 3070 7044 3126 7100
rect 3126 7044 3130 7100
rect 3066 7040 3130 7044
rect 6574 7100 6638 7104
rect 6574 7044 6578 7100
rect 6578 7044 6634 7100
rect 6634 7044 6638 7100
rect 6574 7040 6638 7044
rect 6654 7100 6718 7104
rect 6654 7044 6658 7100
rect 6658 7044 6714 7100
rect 6714 7044 6718 7100
rect 6654 7040 6718 7044
rect 6734 7100 6798 7104
rect 6734 7044 6738 7100
rect 6738 7044 6794 7100
rect 6794 7044 6798 7100
rect 6734 7040 6798 7044
rect 6814 7100 6878 7104
rect 6814 7044 6818 7100
rect 6818 7044 6874 7100
rect 6874 7044 6878 7100
rect 6814 7040 6878 7044
rect 10322 7100 10386 7104
rect 10322 7044 10326 7100
rect 10326 7044 10382 7100
rect 10382 7044 10386 7100
rect 10322 7040 10386 7044
rect 10402 7100 10466 7104
rect 10402 7044 10406 7100
rect 10406 7044 10462 7100
rect 10462 7044 10466 7100
rect 10402 7040 10466 7044
rect 10482 7100 10546 7104
rect 10482 7044 10486 7100
rect 10486 7044 10542 7100
rect 10542 7044 10546 7100
rect 10482 7040 10546 7044
rect 10562 7100 10626 7104
rect 10562 7044 10566 7100
rect 10566 7044 10622 7100
rect 10622 7044 10626 7100
rect 10562 7040 10626 7044
rect 14070 7100 14134 7104
rect 14070 7044 14074 7100
rect 14074 7044 14130 7100
rect 14130 7044 14134 7100
rect 14070 7040 14134 7044
rect 14150 7100 14214 7104
rect 14150 7044 14154 7100
rect 14154 7044 14210 7100
rect 14210 7044 14214 7100
rect 14150 7040 14214 7044
rect 14230 7100 14294 7104
rect 14230 7044 14234 7100
rect 14234 7044 14290 7100
rect 14290 7044 14294 7100
rect 14230 7040 14294 7044
rect 14310 7100 14374 7104
rect 14310 7044 14314 7100
rect 14314 7044 14370 7100
rect 14370 7044 14374 7100
rect 14310 7040 14374 7044
rect 4700 6556 4764 6560
rect 4700 6500 4704 6556
rect 4704 6500 4760 6556
rect 4760 6500 4764 6556
rect 4700 6496 4764 6500
rect 4780 6556 4844 6560
rect 4780 6500 4784 6556
rect 4784 6500 4840 6556
rect 4840 6500 4844 6556
rect 4780 6496 4844 6500
rect 4860 6556 4924 6560
rect 4860 6500 4864 6556
rect 4864 6500 4920 6556
rect 4920 6500 4924 6556
rect 4860 6496 4924 6500
rect 4940 6556 5004 6560
rect 4940 6500 4944 6556
rect 4944 6500 5000 6556
rect 5000 6500 5004 6556
rect 4940 6496 5004 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 12196 6556 12260 6560
rect 12196 6500 12200 6556
rect 12200 6500 12256 6556
rect 12256 6500 12260 6556
rect 12196 6496 12260 6500
rect 12276 6556 12340 6560
rect 12276 6500 12280 6556
rect 12280 6500 12336 6556
rect 12336 6500 12340 6556
rect 12276 6496 12340 6500
rect 12356 6556 12420 6560
rect 12356 6500 12360 6556
rect 12360 6500 12416 6556
rect 12416 6500 12420 6556
rect 12356 6496 12420 6500
rect 12436 6556 12500 6560
rect 12436 6500 12440 6556
rect 12440 6500 12496 6556
rect 12496 6500 12500 6556
rect 12436 6496 12500 6500
rect 2826 6012 2890 6016
rect 2826 5956 2830 6012
rect 2830 5956 2886 6012
rect 2886 5956 2890 6012
rect 2826 5952 2890 5956
rect 2906 6012 2970 6016
rect 2906 5956 2910 6012
rect 2910 5956 2966 6012
rect 2966 5956 2970 6012
rect 2906 5952 2970 5956
rect 2986 6012 3050 6016
rect 2986 5956 2990 6012
rect 2990 5956 3046 6012
rect 3046 5956 3050 6012
rect 2986 5952 3050 5956
rect 3066 6012 3130 6016
rect 3066 5956 3070 6012
rect 3070 5956 3126 6012
rect 3126 5956 3130 6012
rect 3066 5952 3130 5956
rect 6574 6012 6638 6016
rect 6574 5956 6578 6012
rect 6578 5956 6634 6012
rect 6634 5956 6638 6012
rect 6574 5952 6638 5956
rect 6654 6012 6718 6016
rect 6654 5956 6658 6012
rect 6658 5956 6714 6012
rect 6714 5956 6718 6012
rect 6654 5952 6718 5956
rect 6734 6012 6798 6016
rect 6734 5956 6738 6012
rect 6738 5956 6794 6012
rect 6794 5956 6798 6012
rect 6734 5952 6798 5956
rect 6814 6012 6878 6016
rect 6814 5956 6818 6012
rect 6818 5956 6874 6012
rect 6874 5956 6878 6012
rect 6814 5952 6878 5956
rect 10322 6012 10386 6016
rect 10322 5956 10326 6012
rect 10326 5956 10382 6012
rect 10382 5956 10386 6012
rect 10322 5952 10386 5956
rect 10402 6012 10466 6016
rect 10402 5956 10406 6012
rect 10406 5956 10462 6012
rect 10462 5956 10466 6012
rect 10402 5952 10466 5956
rect 10482 6012 10546 6016
rect 10482 5956 10486 6012
rect 10486 5956 10542 6012
rect 10542 5956 10546 6012
rect 10482 5952 10546 5956
rect 10562 6012 10626 6016
rect 10562 5956 10566 6012
rect 10566 5956 10622 6012
rect 10622 5956 10626 6012
rect 10562 5952 10626 5956
rect 14070 6012 14134 6016
rect 14070 5956 14074 6012
rect 14074 5956 14130 6012
rect 14130 5956 14134 6012
rect 14070 5952 14134 5956
rect 14150 6012 14214 6016
rect 14150 5956 14154 6012
rect 14154 5956 14210 6012
rect 14210 5956 14214 6012
rect 14150 5952 14214 5956
rect 14230 6012 14294 6016
rect 14230 5956 14234 6012
rect 14234 5956 14290 6012
rect 14290 5956 14294 6012
rect 14230 5952 14294 5956
rect 14310 6012 14374 6016
rect 14310 5956 14314 6012
rect 14314 5956 14370 6012
rect 14370 5956 14374 6012
rect 14310 5952 14374 5956
rect 4700 5468 4764 5472
rect 4700 5412 4704 5468
rect 4704 5412 4760 5468
rect 4760 5412 4764 5468
rect 4700 5408 4764 5412
rect 4780 5468 4844 5472
rect 4780 5412 4784 5468
rect 4784 5412 4840 5468
rect 4840 5412 4844 5468
rect 4780 5408 4844 5412
rect 4860 5468 4924 5472
rect 4860 5412 4864 5468
rect 4864 5412 4920 5468
rect 4920 5412 4924 5468
rect 4860 5408 4924 5412
rect 4940 5468 5004 5472
rect 4940 5412 4944 5468
rect 4944 5412 5000 5468
rect 5000 5412 5004 5468
rect 4940 5408 5004 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 12196 5468 12260 5472
rect 12196 5412 12200 5468
rect 12200 5412 12256 5468
rect 12256 5412 12260 5468
rect 12196 5408 12260 5412
rect 12276 5468 12340 5472
rect 12276 5412 12280 5468
rect 12280 5412 12336 5468
rect 12336 5412 12340 5468
rect 12276 5408 12340 5412
rect 12356 5468 12420 5472
rect 12356 5412 12360 5468
rect 12360 5412 12416 5468
rect 12416 5412 12420 5468
rect 12356 5408 12420 5412
rect 12436 5468 12500 5472
rect 12436 5412 12440 5468
rect 12440 5412 12496 5468
rect 12496 5412 12500 5468
rect 12436 5408 12500 5412
rect 2826 4924 2890 4928
rect 2826 4868 2830 4924
rect 2830 4868 2886 4924
rect 2886 4868 2890 4924
rect 2826 4864 2890 4868
rect 2906 4924 2970 4928
rect 2906 4868 2910 4924
rect 2910 4868 2966 4924
rect 2966 4868 2970 4924
rect 2906 4864 2970 4868
rect 2986 4924 3050 4928
rect 2986 4868 2990 4924
rect 2990 4868 3046 4924
rect 3046 4868 3050 4924
rect 2986 4864 3050 4868
rect 3066 4924 3130 4928
rect 3066 4868 3070 4924
rect 3070 4868 3126 4924
rect 3126 4868 3130 4924
rect 3066 4864 3130 4868
rect 6574 4924 6638 4928
rect 6574 4868 6578 4924
rect 6578 4868 6634 4924
rect 6634 4868 6638 4924
rect 6574 4864 6638 4868
rect 6654 4924 6718 4928
rect 6654 4868 6658 4924
rect 6658 4868 6714 4924
rect 6714 4868 6718 4924
rect 6654 4864 6718 4868
rect 6734 4924 6798 4928
rect 6734 4868 6738 4924
rect 6738 4868 6794 4924
rect 6794 4868 6798 4924
rect 6734 4864 6798 4868
rect 6814 4924 6878 4928
rect 6814 4868 6818 4924
rect 6818 4868 6874 4924
rect 6874 4868 6878 4924
rect 6814 4864 6878 4868
rect 10322 4924 10386 4928
rect 10322 4868 10326 4924
rect 10326 4868 10382 4924
rect 10382 4868 10386 4924
rect 10322 4864 10386 4868
rect 10402 4924 10466 4928
rect 10402 4868 10406 4924
rect 10406 4868 10462 4924
rect 10462 4868 10466 4924
rect 10402 4864 10466 4868
rect 10482 4924 10546 4928
rect 10482 4868 10486 4924
rect 10486 4868 10542 4924
rect 10542 4868 10546 4924
rect 10482 4864 10546 4868
rect 10562 4924 10626 4928
rect 10562 4868 10566 4924
rect 10566 4868 10622 4924
rect 10622 4868 10626 4924
rect 10562 4864 10626 4868
rect 14070 4924 14134 4928
rect 14070 4868 14074 4924
rect 14074 4868 14130 4924
rect 14130 4868 14134 4924
rect 14070 4864 14134 4868
rect 14150 4924 14214 4928
rect 14150 4868 14154 4924
rect 14154 4868 14210 4924
rect 14210 4868 14214 4924
rect 14150 4864 14214 4868
rect 14230 4924 14294 4928
rect 14230 4868 14234 4924
rect 14234 4868 14290 4924
rect 14290 4868 14294 4924
rect 14230 4864 14294 4868
rect 14310 4924 14374 4928
rect 14310 4868 14314 4924
rect 14314 4868 14370 4924
rect 14370 4868 14374 4924
rect 14310 4864 14374 4868
rect 4700 4380 4764 4384
rect 4700 4324 4704 4380
rect 4704 4324 4760 4380
rect 4760 4324 4764 4380
rect 4700 4320 4764 4324
rect 4780 4380 4844 4384
rect 4780 4324 4784 4380
rect 4784 4324 4840 4380
rect 4840 4324 4844 4380
rect 4780 4320 4844 4324
rect 4860 4380 4924 4384
rect 4860 4324 4864 4380
rect 4864 4324 4920 4380
rect 4920 4324 4924 4380
rect 4860 4320 4924 4324
rect 4940 4380 5004 4384
rect 4940 4324 4944 4380
rect 4944 4324 5000 4380
rect 5000 4324 5004 4380
rect 4940 4320 5004 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 12196 4380 12260 4384
rect 12196 4324 12200 4380
rect 12200 4324 12256 4380
rect 12256 4324 12260 4380
rect 12196 4320 12260 4324
rect 12276 4380 12340 4384
rect 12276 4324 12280 4380
rect 12280 4324 12336 4380
rect 12336 4324 12340 4380
rect 12276 4320 12340 4324
rect 12356 4380 12420 4384
rect 12356 4324 12360 4380
rect 12360 4324 12416 4380
rect 12416 4324 12420 4380
rect 12356 4320 12420 4324
rect 12436 4380 12500 4384
rect 12436 4324 12440 4380
rect 12440 4324 12496 4380
rect 12496 4324 12500 4380
rect 12436 4320 12500 4324
rect 2826 3836 2890 3840
rect 2826 3780 2830 3836
rect 2830 3780 2886 3836
rect 2886 3780 2890 3836
rect 2826 3776 2890 3780
rect 2906 3836 2970 3840
rect 2906 3780 2910 3836
rect 2910 3780 2966 3836
rect 2966 3780 2970 3836
rect 2906 3776 2970 3780
rect 2986 3836 3050 3840
rect 2986 3780 2990 3836
rect 2990 3780 3046 3836
rect 3046 3780 3050 3836
rect 2986 3776 3050 3780
rect 3066 3836 3130 3840
rect 3066 3780 3070 3836
rect 3070 3780 3126 3836
rect 3126 3780 3130 3836
rect 3066 3776 3130 3780
rect 6574 3836 6638 3840
rect 6574 3780 6578 3836
rect 6578 3780 6634 3836
rect 6634 3780 6638 3836
rect 6574 3776 6638 3780
rect 6654 3836 6718 3840
rect 6654 3780 6658 3836
rect 6658 3780 6714 3836
rect 6714 3780 6718 3836
rect 6654 3776 6718 3780
rect 6734 3836 6798 3840
rect 6734 3780 6738 3836
rect 6738 3780 6794 3836
rect 6794 3780 6798 3836
rect 6734 3776 6798 3780
rect 6814 3836 6878 3840
rect 6814 3780 6818 3836
rect 6818 3780 6874 3836
rect 6874 3780 6878 3836
rect 6814 3776 6878 3780
rect 10322 3836 10386 3840
rect 10322 3780 10326 3836
rect 10326 3780 10382 3836
rect 10382 3780 10386 3836
rect 10322 3776 10386 3780
rect 10402 3836 10466 3840
rect 10402 3780 10406 3836
rect 10406 3780 10462 3836
rect 10462 3780 10466 3836
rect 10402 3776 10466 3780
rect 10482 3836 10546 3840
rect 10482 3780 10486 3836
rect 10486 3780 10542 3836
rect 10542 3780 10546 3836
rect 10482 3776 10546 3780
rect 10562 3836 10626 3840
rect 10562 3780 10566 3836
rect 10566 3780 10622 3836
rect 10622 3780 10626 3836
rect 10562 3776 10626 3780
rect 14070 3836 14134 3840
rect 14070 3780 14074 3836
rect 14074 3780 14130 3836
rect 14130 3780 14134 3836
rect 14070 3776 14134 3780
rect 14150 3836 14214 3840
rect 14150 3780 14154 3836
rect 14154 3780 14210 3836
rect 14210 3780 14214 3836
rect 14150 3776 14214 3780
rect 14230 3836 14294 3840
rect 14230 3780 14234 3836
rect 14234 3780 14290 3836
rect 14290 3780 14294 3836
rect 14230 3776 14294 3780
rect 14310 3836 14374 3840
rect 14310 3780 14314 3836
rect 14314 3780 14370 3836
rect 14370 3780 14374 3836
rect 14310 3776 14374 3780
rect 4700 3292 4764 3296
rect 4700 3236 4704 3292
rect 4704 3236 4760 3292
rect 4760 3236 4764 3292
rect 4700 3232 4764 3236
rect 4780 3292 4844 3296
rect 4780 3236 4784 3292
rect 4784 3236 4840 3292
rect 4840 3236 4844 3292
rect 4780 3232 4844 3236
rect 4860 3292 4924 3296
rect 4860 3236 4864 3292
rect 4864 3236 4920 3292
rect 4920 3236 4924 3292
rect 4860 3232 4924 3236
rect 4940 3292 5004 3296
rect 4940 3236 4944 3292
rect 4944 3236 5000 3292
rect 5000 3236 5004 3292
rect 4940 3232 5004 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 12196 3292 12260 3296
rect 12196 3236 12200 3292
rect 12200 3236 12256 3292
rect 12256 3236 12260 3292
rect 12196 3232 12260 3236
rect 12276 3292 12340 3296
rect 12276 3236 12280 3292
rect 12280 3236 12336 3292
rect 12336 3236 12340 3292
rect 12276 3232 12340 3236
rect 12356 3292 12420 3296
rect 12356 3236 12360 3292
rect 12360 3236 12416 3292
rect 12416 3236 12420 3292
rect 12356 3232 12420 3236
rect 12436 3292 12500 3296
rect 12436 3236 12440 3292
rect 12440 3236 12496 3292
rect 12496 3236 12500 3292
rect 12436 3232 12500 3236
rect 2826 2748 2890 2752
rect 2826 2692 2830 2748
rect 2830 2692 2886 2748
rect 2886 2692 2890 2748
rect 2826 2688 2890 2692
rect 2906 2748 2970 2752
rect 2906 2692 2910 2748
rect 2910 2692 2966 2748
rect 2966 2692 2970 2748
rect 2906 2688 2970 2692
rect 2986 2748 3050 2752
rect 2986 2692 2990 2748
rect 2990 2692 3046 2748
rect 3046 2692 3050 2748
rect 2986 2688 3050 2692
rect 3066 2748 3130 2752
rect 3066 2692 3070 2748
rect 3070 2692 3126 2748
rect 3126 2692 3130 2748
rect 3066 2688 3130 2692
rect 6574 2748 6638 2752
rect 6574 2692 6578 2748
rect 6578 2692 6634 2748
rect 6634 2692 6638 2748
rect 6574 2688 6638 2692
rect 6654 2748 6718 2752
rect 6654 2692 6658 2748
rect 6658 2692 6714 2748
rect 6714 2692 6718 2748
rect 6654 2688 6718 2692
rect 6734 2748 6798 2752
rect 6734 2692 6738 2748
rect 6738 2692 6794 2748
rect 6794 2692 6798 2748
rect 6734 2688 6798 2692
rect 6814 2748 6878 2752
rect 6814 2692 6818 2748
rect 6818 2692 6874 2748
rect 6874 2692 6878 2748
rect 6814 2688 6878 2692
rect 10322 2748 10386 2752
rect 10322 2692 10326 2748
rect 10326 2692 10382 2748
rect 10382 2692 10386 2748
rect 10322 2688 10386 2692
rect 10402 2748 10466 2752
rect 10402 2692 10406 2748
rect 10406 2692 10462 2748
rect 10462 2692 10466 2748
rect 10402 2688 10466 2692
rect 10482 2748 10546 2752
rect 10482 2692 10486 2748
rect 10486 2692 10542 2748
rect 10542 2692 10546 2748
rect 10482 2688 10546 2692
rect 10562 2748 10626 2752
rect 10562 2692 10566 2748
rect 10566 2692 10622 2748
rect 10622 2692 10626 2748
rect 10562 2688 10626 2692
rect 14070 2748 14134 2752
rect 14070 2692 14074 2748
rect 14074 2692 14130 2748
rect 14130 2692 14134 2748
rect 14070 2688 14134 2692
rect 14150 2748 14214 2752
rect 14150 2692 14154 2748
rect 14154 2692 14210 2748
rect 14210 2692 14214 2748
rect 14150 2688 14214 2692
rect 14230 2748 14294 2752
rect 14230 2692 14234 2748
rect 14234 2692 14290 2748
rect 14290 2692 14294 2748
rect 14230 2688 14294 2692
rect 14310 2748 14374 2752
rect 14310 2692 14314 2748
rect 14314 2692 14370 2748
rect 14370 2692 14374 2748
rect 14310 2688 14374 2692
rect 4700 2204 4764 2208
rect 4700 2148 4704 2204
rect 4704 2148 4760 2204
rect 4760 2148 4764 2204
rect 4700 2144 4764 2148
rect 4780 2204 4844 2208
rect 4780 2148 4784 2204
rect 4784 2148 4840 2204
rect 4840 2148 4844 2204
rect 4780 2144 4844 2148
rect 4860 2204 4924 2208
rect 4860 2148 4864 2204
rect 4864 2148 4920 2204
rect 4920 2148 4924 2204
rect 4860 2144 4924 2148
rect 4940 2204 5004 2208
rect 4940 2148 4944 2204
rect 4944 2148 5000 2204
rect 5000 2148 5004 2204
rect 4940 2144 5004 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 12196 2204 12260 2208
rect 12196 2148 12200 2204
rect 12200 2148 12256 2204
rect 12256 2148 12260 2204
rect 12196 2144 12260 2148
rect 12276 2204 12340 2208
rect 12276 2148 12280 2204
rect 12280 2148 12336 2204
rect 12336 2148 12340 2204
rect 12276 2144 12340 2148
rect 12356 2204 12420 2208
rect 12356 2148 12360 2204
rect 12360 2148 12416 2204
rect 12416 2148 12420 2204
rect 12356 2144 12420 2148
rect 12436 2204 12500 2208
rect 12436 2148 12440 2204
rect 12440 2148 12496 2204
rect 12496 2148 12500 2204
rect 12436 2144 12500 2148
<< metal4 >>
rect 2818 16896 3138 17456
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 15808 3138 16832
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 2818 14720 3138 15744
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 2818 13632 3138 14656
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 12544 3138 13568
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2818 11456 3138 12480
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 10368 3138 11392
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 2818 9280 3138 10304
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 8192 3138 9216
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 7104 3138 8128
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2818 6016 3138 7040
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2818 4928 3138 5952
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 2818 3840 3138 4864
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2818 2752 3138 3776
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 2818 2128 3138 2688
rect 4692 17440 5012 17456
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 4692 16352 5012 17376
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4692 15264 5012 16288
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4692 14176 5012 15200
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 4692 13088 5012 14112
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 4692 12000 5012 13024
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4692 10912 5012 11936
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 4692 9824 5012 10848
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 4692 8736 5012 9760
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 4692 7648 5012 8672
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4692 6560 5012 7584
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 4692 5472 5012 6496
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4692 4384 5012 5408
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 4692 3296 5012 4320
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 4692 2208 5012 3232
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2128 5012 2144
rect 6566 16896 6886 17456
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 6566 15808 6886 16832
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 6566 14720 6886 15744
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 13632 6886 14656
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6566 12544 6886 13568
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 6566 11456 6886 12480
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6566 10368 6886 11392
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 6566 9280 6886 10304
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6566 8192 6886 9216
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 7104 6886 8128
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 6566 6016 6886 7040
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 6566 4928 6886 5952
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 6566 3840 6886 4864
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 6566 2752 6886 3776
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 6566 2128 6886 2688
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 10314 16896 10634 17456
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 10314 15808 10634 16832
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 10314 14720 10634 15744
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 10314 13632 10634 14656
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 10314 12544 10634 13568
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10314 11456 10634 12480
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 8891 11252 8957 11253
rect 8891 11188 8892 11252
rect 8956 11188 8957 11252
rect 8891 11187 8957 11188
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 8894 9757 8954 11187
rect 10314 10368 10634 11392
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 8891 9756 8957 9757
rect 8891 9692 8892 9756
rect 8956 9692 8957 9756
rect 8891 9691 8957 9692
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 2208 8760 3232
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 10314 9280 10634 10304
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 10314 8192 10634 9216
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10314 7104 10634 8128
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 10314 6016 10634 7040
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 10314 4928 10634 5952
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 10314 3840 10634 4864
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 10314 2752 10634 3776
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 10314 2128 10634 2688
rect 12188 17440 12508 17456
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 12188 16352 12508 17376
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 12188 15264 12508 16288
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12188 14176 12508 15200
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 12188 13088 12508 14112
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12188 12000 12508 13024
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 10912 12508 11936
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12188 9824 12508 10848
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 12188 8736 12508 9760
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 12188 7648 12508 8672
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12188 6560 12508 7584
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 12188 5472 12508 6496
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 12188 4384 12508 5408
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12188 3296 12508 4320
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 12188 2208 12508 3232
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2128 12508 2144
rect 14062 16896 14382 17456
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 14062 15808 14382 16832
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 14062 14720 14382 15744
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 14062 13632 14382 14656
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 14062 12544 14382 13568
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 14062 11456 14382 12480
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 14062 10368 14382 11392
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 14062 9280 14382 10304
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 14062 8192 14382 9216
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 14062 7104 14382 8128
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 14062 6016 14382 7040
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 14062 4928 14382 5952
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 3840 14382 4864
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 14062 2752 14382 3776
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 14062 2128 14382 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__02__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5520 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__03__A
timestamp 1649977179
transform -1 0 5612 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__04__A
timestamp 1649977179
transform -1 0 6072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__05__A
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__06__A
timestamp 1649977179
transform -1 0 6440 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__07__A
timestamp 1649977179
transform -1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__08__A
timestamp 1649977179
transform -1 0 8096 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__09__A
timestamp 1649977179
transform -1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__10__A
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__11__A
timestamp 1649977179
transform -1 0 7912 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__12__A
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__13__A
timestamp 1649977179
transform 1 0 9936 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__14__A
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__15__A
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__16__A
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__17__A
timestamp 1649977179
transform -1 0 9844 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1649977179
transform -1 0 13432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1649977179
transform 1 0 12696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1649977179
transform 1 0 12880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1649977179
transform 1 0 14076 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1649977179
transform -1 0 5060 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1649977179
transform -1 0 5612 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1649977179
transform -1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1649977179
transform -1 0 6164 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1649977179
transform -1 0 6440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1649977179
transform -1 0 6808 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1649977179
transform -1 0 6624 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1649977179
transform -1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1649977179
transform 1 0 10120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1649977179
transform -1 0 7912 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1649977179
transform -1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1649977179
transform -1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform 1 0 11776 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform -1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform 1 0 12144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform -1 0 5060 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform 1 0 5336 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 4324 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 9016 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 9752 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10488 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_153 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_149 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_157 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15548 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_157
timestamp 1649977179
transform 1 0 15548 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp 1649977179
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1649977179
transform 1 0 4324 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_65
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_74
timestamp 1649977179
transform 1 0 7912 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_86
timestamp 1649977179
transform 1 0 9016 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_94
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_157
timestamp 1649977179
transform 1 0 15548 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_88
timestamp 1649977179
transform 1 0 9200 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_100
timestamp 1649977179
transform 1 0 10304 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_127
timestamp 1649977179
transform 1 0 12788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_139
timestamp 1649977179
transform 1 0 13892 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_151
timestamp 1649977179
transform 1 0 14996 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_5
timestamp 1649977179
transform 1 0 1564 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_17
timestamp 1649977179
transform 1 0 2668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1649977179
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_47
timestamp 1649977179
transform 1 0 5428 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_50
timestamp 1649977179
transform 1 0 5704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_54
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1649977179
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_78
timestamp 1649977179
transform 1 0 8280 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_100
timestamp 1649977179
transform 1 0 10304 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_112
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_124
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_16
timestamp 1649977179
transform 1 0 2576 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_28
timestamp 1649977179
transform 1 0 3680 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_40
timestamp 1649977179
transform 1 0 4784 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_96
timestamp 1649977179
transform 1 0 9936 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 1649977179
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_130
timestamp 1649977179
transform 1 0 13064 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_142
timestamp 1649977179
transform 1 0 14168 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_154
timestamp 1649977179
transform 1 0 15272 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_158
timestamp 1649977179
transform 1 0 15640 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_37
timestamp 1649977179
transform 1 0 4508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_23
timestamp 1649977179
transform 1 0 3220 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_28
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_40
timestamp 1649977179
transform 1 0 4784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_45
timestamp 1649977179
transform 1 0 5244 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_104
timestamp 1649977179
transform 1 0 10672 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_115
timestamp 1649977179
transform 1 0 11684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1649977179
transform 1 0 11960 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_122
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_134
timestamp 1649977179
transform 1 0 13432 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_146
timestamp 1649977179
transform 1 0 14536 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_49
timestamp 1649977179
transform 1 0 5612 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_54
timestamp 1649977179
transform 1 0 6072 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_96
timestamp 1649977179
transform 1 0 9936 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_108
timestamp 1649977179
transform 1 0 11040 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_120
timestamp 1649977179
transform 1 0 12144 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_132
timestamp 1649977179
transform 1 0 13248 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_63
timestamp 1649977179
transform 1 0 6900 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_74
timestamp 1649977179
transform 1 0 7912 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_100
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_49
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_61
timestamp 1649977179
transform 1 0 6716 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_67
timestamp 1649977179
transform 1 0 7268 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_76
timestamp 1649977179
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_95
timestamp 1649977179
transform 1 0 9844 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_107
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_119
timestamp 1649977179
transform 1 0 12052 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp 1649977179
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_59
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_71
timestamp 1649977179
transform 1 0 7636 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_83
timestamp 1649977179
transform 1 0 8740 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_95
timestamp 1649977179
transform 1 0 9844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1649977179
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_147
timestamp 1649977179
transform 1 0 14628 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1649977179
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_157
timestamp 1649977179
transform 1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_29
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_41
timestamp 1649977179
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1649977179
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1649977179
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1649977179
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_141
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_153
timestamp 1649977179
transform 1 0 15180 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _01_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8648 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _02_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5520 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _03_
timestamp 1649977179
transform -1 0 5428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _04_
timestamp 1649977179
transform -1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1649977179
transform -1 0 6164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _06_
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _07_
timestamp 1649977179
transform -1 0 7544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1649977179
transform -1 0 7912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _09_
timestamp 1649977179
transform -1 0 6900 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1649977179
transform -1 0 8740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1649977179
transform -1 0 7728 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1649977179
transform -1 0 9568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1649977179
transform -1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1649977179
transform -1 0 10396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1649977179
transform -1 0 10764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1649977179
transform -1 0 11132 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1649977179
transform -1 0 9660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1649977179
transform -1 0 12512 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1649977179
transform -1 0 12328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1649977179
transform -1 0 12696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1649977179
transform 1 0 14260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1649977179
transform -1 0 4876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1649977179
transform -1 0 5060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1649977179
transform -1 0 5428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1649977179
transform -1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1649977179
transform -1 0 5980 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1649977179
transform -1 0 6256 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1649977179
transform -1 0 7176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1649977179
transform -1 0 6900 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1649977179
transform -1 0 8372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1649977179
transform -1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1649977179
transform -1 0 7728 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1649977179
transform -1 0 9568 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1649977179
transform -1 0 9936 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1649977179
transform -1 0 11040 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1649977179
transform -1 0 11408 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1649977179
transform -1 0 11776 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1649977179
transform -1 0 9568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1649977179
transform -1 0 12144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1649977179
transform -1 0 12880 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1649977179
transform -1 0 13248 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1649977179
transform -1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5888 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7728 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7176 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8372 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6808 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7728 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8832 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8372 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9844 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8004 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9016 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 7176 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5060 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12604 0 -1 8704
box -38 -48 1142 592
<< labels >>
flabel metal2 s 1214 19200 1270 20000 0 FreeSans 224 90 0 0 IO_ISOL_N
port 0 nsew signal input
flabel metal4 s 4692 2128 5012 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 8440 2128 8760 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 12188 2128 12508 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 2818 2128 3138 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 6566 2128 6886 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 10314 2128 10634 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 14062 2128 14382 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal3 s 0 18096 800 18216 0 FreeSans 480 0 0 0 ccff_head
port 3 nsew signal input
flabel metal3 s 16400 12384 17200 12504 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 5 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 6 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 7 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 8 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 9 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 10 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 11 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 12 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 13 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 14 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 15 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 16 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 17 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 18 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 19 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 20 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 21 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 22 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 23 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 24 nsew signal input
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 25 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 26 nsew signal tristate
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 27 nsew signal tristate
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 28 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 29 nsew signal tristate
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 30 nsew signal tristate
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 31 nsew signal tristate
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 32 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 33 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 34 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 35 nsew signal tristate
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 36 nsew signal tristate
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 37 nsew signal tristate
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 38 nsew signal tristate
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 39 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 40 nsew signal tristate
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 41 nsew signal tristate
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 42 nsew signal tristate
flabel metal2 s 4342 0 4398 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 43 nsew signal tristate
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 44 nsew signal tristate
flabel metal2 s 8942 19200 8998 20000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 45 nsew signal input
flabel metal2 s 12622 19200 12678 20000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 46 nsew signal input
flabel metal2 s 12990 19200 13046 20000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 47 nsew signal input
flabel metal2 s 13358 19200 13414 20000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 48 nsew signal input
flabel metal2 s 13726 19200 13782 20000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 49 nsew signal input
flabel metal2 s 14094 19200 14150 20000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 50 nsew signal input
flabel metal2 s 14462 19200 14518 20000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 51 nsew signal input
flabel metal2 s 14830 19200 14886 20000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 52 nsew signal input
flabel metal2 s 15198 19200 15254 20000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 53 nsew signal input
flabel metal2 s 15566 19200 15622 20000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 54 nsew signal input
flabel metal2 s 15934 19200 15990 20000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 55 nsew signal input
flabel metal2 s 9310 19200 9366 20000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 56 nsew signal input
flabel metal2 s 9678 19200 9734 20000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 57 nsew signal input
flabel metal2 s 10046 19200 10102 20000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 58 nsew signal input
flabel metal2 s 10414 19200 10470 20000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 59 nsew signal input
flabel metal2 s 10782 19200 10838 20000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 60 nsew signal input
flabel metal2 s 11150 19200 11206 20000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 61 nsew signal input
flabel metal2 s 11518 19200 11574 20000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 62 nsew signal input
flabel metal2 s 11886 19200 11942 20000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 63 nsew signal input
flabel metal2 s 12254 19200 12310 20000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 64 nsew signal input
flabel metal2 s 1582 19200 1638 20000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 65 nsew signal tristate
flabel metal2 s 5262 19200 5318 20000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 66 nsew signal tristate
flabel metal2 s 5630 19200 5686 20000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 67 nsew signal tristate
flabel metal2 s 5998 19200 6054 20000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 68 nsew signal tristate
flabel metal2 s 6366 19200 6422 20000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 69 nsew signal tristate
flabel metal2 s 6734 19200 6790 20000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 70 nsew signal tristate
flabel metal2 s 7102 19200 7158 20000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 71 nsew signal tristate
flabel metal2 s 7470 19200 7526 20000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 72 nsew signal tristate
flabel metal2 s 7838 19200 7894 20000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 73 nsew signal tristate
flabel metal2 s 8206 19200 8262 20000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 74 nsew signal tristate
flabel metal2 s 8574 19200 8630 20000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 75 nsew signal tristate
flabel metal2 s 1950 19200 2006 20000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 76 nsew signal tristate
flabel metal2 s 2318 19200 2374 20000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 77 nsew signal tristate
flabel metal2 s 2686 19200 2742 20000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 78 nsew signal tristate
flabel metal2 s 3054 19200 3110 20000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 79 nsew signal tristate
flabel metal2 s 3422 19200 3478 20000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 80 nsew signal tristate
flabel metal2 s 3790 19200 3846 20000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 81 nsew signal tristate
flabel metal2 s 4158 19200 4214 20000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 82 nsew signal tristate
flabel metal2 s 4526 19200 4582 20000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 83 nsew signal tristate
flabel metal2 s 4894 19200 4950 20000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 84 nsew signal tristate
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 85 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 86 nsew signal input
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 87 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 left_grid_pin_0_
port 88 nsew signal tristate
flabel metal3 s 16400 7488 17200 7608 0 FreeSans 480 0 0 0 prog_clk_0_E_in
port 89 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_0_
port 90 nsew signal input
flabel metal3 s 16400 2592 17200 2712 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_1_lower
port 91 nsew signal tristate
flabel metal3 s 16400 17280 17200 17400 0 FreeSans 480 0 0 0 right_width_0_height_0__pin_1_upper
port 92 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
