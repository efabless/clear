magic
tech sky130A
magscale 1 2
timestamp 1679357742
<< viali >>
rect 9137 24361 9171 24395
rect 25789 24361 25823 24395
rect 32321 24361 32355 24395
rect 33425 24361 33459 24395
rect 34161 24361 34195 24395
rect 35081 24361 35115 24395
rect 35817 24361 35851 24395
rect 39313 24361 39347 24395
rect 11713 24293 11747 24327
rect 19441 24293 19475 24327
rect 46857 24293 46891 24327
rect 3249 24225 3283 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 13553 24225 13587 24259
rect 16865 24225 16899 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25237 24225 25271 24259
rect 26341 24225 26375 24259
rect 27721 24225 27755 24259
rect 29745 24225 29779 24259
rect 30021 24225 30055 24259
rect 40049 24225 40083 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 6745 24157 6779 24191
rect 7205 24157 7239 24191
rect 9321 24157 9355 24191
rect 9965 24157 9999 24191
rect 10885 24157 10919 24191
rect 11897 24157 11931 24191
rect 12541 24157 12575 24191
rect 14473 24157 14507 24191
rect 14933 24157 14967 24191
rect 19625 24157 19659 24191
rect 20085 24157 20119 24191
rect 22109 24157 22143 24191
rect 24041 24157 24075 24191
rect 28549 24157 28583 24191
rect 29193 24157 29227 24191
rect 31493 24157 31527 24191
rect 32505 24157 32539 24191
rect 33333 24157 33367 24191
rect 34069 24157 34103 24191
rect 34989 24157 35023 24191
rect 35725 24157 35759 24191
rect 36553 24157 36587 24191
rect 37657 24157 37691 24191
rect 38485 24157 38519 24191
rect 38669 24157 38703 24191
rect 39221 24157 39255 24191
rect 40325 24157 40359 24191
rect 41521 24157 41555 24191
rect 42625 24157 42659 24191
rect 45201 24157 45235 24191
rect 45937 24157 45971 24191
rect 46673 24157 46707 24191
rect 47777 24157 47811 24191
rect 48513 24157 48547 24191
rect 16129 24089 16163 24123
rect 17141 24089 17175 24123
rect 27629 24089 27663 24123
rect 6561 24021 6595 24055
rect 14289 24021 14323 24055
rect 18613 24021 18647 24055
rect 23857 24021 23891 24055
rect 24593 24021 24627 24055
rect 24961 24021 24995 24055
rect 25053 24021 25087 24055
rect 26157 24021 26191 24055
rect 26249 24021 26283 24055
rect 27169 24021 27203 24055
rect 27537 24021 27571 24055
rect 28365 24021 28399 24055
rect 29009 24021 29043 24055
rect 31309 24021 31343 24055
rect 36369 24021 36403 24055
rect 37473 24021 37507 24055
rect 41337 24021 41371 24055
rect 43913 24021 43947 24055
rect 45385 24021 45419 24055
rect 46121 24021 46155 24055
rect 47961 24021 47995 24055
rect 48697 24021 48731 24055
rect 11897 23817 11931 23851
rect 12265 23817 12299 23851
rect 12357 23817 12391 23851
rect 32321 23817 32355 23851
rect 35173 23817 35207 23851
rect 2145 23749 2179 23783
rect 3985 23749 4019 23783
rect 9137 23749 9171 23783
rect 10977 23749 11011 23783
rect 14289 23749 14323 23783
rect 18153 23749 18187 23783
rect 27445 23749 27479 23783
rect 34529 23749 34563 23783
rect 36001 23749 36035 23783
rect 43637 23749 43671 23783
rect 2789 23681 2823 23715
rect 4629 23681 4663 23715
rect 6653 23681 6687 23715
rect 7481 23681 7515 23715
rect 8125 23681 8159 23715
rect 9965 23681 9999 23715
rect 13277 23681 13311 23715
rect 15117 23681 15151 23715
rect 16957 23681 16991 23715
rect 21097 23681 21131 23715
rect 24409 23681 24443 23715
rect 27169 23681 27203 23715
rect 29561 23681 29595 23715
rect 30021 23681 30055 23715
rect 31493 23681 31527 23715
rect 32505 23681 32539 23715
rect 33149 23681 33183 23715
rect 33793 23681 33827 23715
rect 34345 23681 34379 23715
rect 35081 23681 35115 23715
rect 35817 23681 35851 23715
rect 36645 23681 36679 23715
rect 37933 23681 37967 23715
rect 41521 23681 41555 23715
rect 44281 23681 44315 23715
rect 46765 23681 46799 23715
rect 48329 23681 48363 23715
rect 49065 23681 49099 23715
rect 5457 23613 5491 23647
rect 12541 23613 12575 23647
rect 16129 23613 16163 23647
rect 18797 23613 18831 23647
rect 19073 23613 19107 23647
rect 22017 23613 22051 23647
rect 22293 23613 22327 23647
rect 24869 23613 24903 23647
rect 25145 23613 25179 23647
rect 30297 23613 30331 23647
rect 2329 23545 2363 23579
rect 21281 23545 21315 23579
rect 29377 23545 29411 23579
rect 33609 23545 33643 23579
rect 43821 23545 43855 23579
rect 44465 23545 44499 23579
rect 6745 23477 6779 23511
rect 7297 23477 7331 23511
rect 20545 23477 20579 23511
rect 23765 23477 23799 23511
rect 26617 23477 26651 23511
rect 28917 23477 28951 23511
rect 31309 23477 31343 23511
rect 32965 23477 32999 23511
rect 36461 23477 36495 23511
rect 37749 23477 37783 23511
rect 41337 23477 41371 23511
rect 46949 23477 46983 23511
rect 48513 23477 48547 23511
rect 49249 23477 49283 23511
rect 14473 23273 14507 23307
rect 19441 23273 19475 23307
rect 32137 23273 32171 23307
rect 5365 23205 5399 23239
rect 18889 23205 18923 23239
rect 29101 23205 29135 23239
rect 3985 23137 4019 23171
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 11437 23137 11471 23171
rect 16497 23137 16531 23171
rect 20085 23137 20119 23171
rect 22569 23137 22603 23171
rect 25145 23137 25179 23171
rect 26341 23137 26375 23171
rect 27353 23137 27387 23171
rect 29745 23137 29779 23171
rect 1777 23069 1811 23103
rect 4261 23069 4295 23103
rect 5457 23069 5491 23103
rect 7297 23069 7331 23103
rect 9229 23069 9263 23103
rect 15485 23069 15519 23103
rect 17141 23069 17175 23103
rect 19625 23069 19659 23103
rect 22293 23069 22327 23103
rect 26157 23069 26191 23103
rect 33425 23069 33459 23103
rect 48605 23069 48639 23103
rect 49065 23069 49099 23103
rect 2789 23001 2823 23035
rect 9505 23001 9539 23035
rect 11713 23001 11747 23035
rect 14381 23001 14415 23035
rect 17417 23001 17451 23035
rect 20361 23001 20395 23035
rect 25053 23001 25087 23035
rect 27629 23001 27663 23035
rect 30021 23001 30055 23035
rect 32689 23001 32723 23035
rect 34161 23001 34195 23035
rect 10977 22933 11011 22967
rect 13185 22933 13219 22967
rect 21833 22933 21867 22967
rect 24041 22933 24075 22967
rect 24593 22933 24627 22967
rect 24961 22933 24995 22967
rect 25789 22933 25823 22967
rect 26249 22933 26283 22967
rect 31493 22933 31527 22967
rect 32781 22933 32815 22967
rect 33517 22933 33551 22967
rect 34253 22933 34287 22967
rect 48421 22933 48455 22967
rect 49249 22933 49283 22967
rect 21465 22729 21499 22763
rect 25789 22729 25823 22763
rect 27629 22729 27663 22763
rect 32505 22729 32539 22763
rect 3801 22661 3835 22695
rect 7113 22661 7147 22695
rect 7941 22661 7975 22695
rect 10701 22661 10735 22695
rect 16129 22661 16163 22695
rect 19993 22661 20027 22695
rect 28641 22661 28675 22695
rect 31033 22661 31067 22695
rect 1685 22593 1719 22627
rect 4721 22593 4755 22627
rect 7205 22593 7239 22627
rect 8125 22593 8159 22627
rect 9965 22593 9999 22627
rect 11805 22593 11839 22627
rect 15117 22593 15151 22627
rect 16865 22593 16899 22627
rect 19257 22593 19291 22627
rect 19717 22593 19751 22627
rect 22661 22593 22695 22627
rect 25697 22593 25731 22627
rect 27537 22593 27571 22627
rect 28365 22593 28399 22627
rect 30941 22593 30975 22627
rect 32413 22593 32447 22627
rect 33149 22593 33183 22627
rect 34253 22593 34287 22627
rect 37933 22593 37967 22627
rect 2789 22525 2823 22559
rect 3893 22525 3927 22559
rect 4077 22525 4111 22559
rect 5089 22525 5123 22559
rect 7389 22525 7423 22559
rect 8677 22525 8711 22559
rect 12449 22525 12483 22559
rect 17141 22525 17175 22559
rect 18613 22525 18647 22559
rect 23121 22525 23155 22559
rect 23397 22525 23431 22559
rect 25881 22525 25915 22559
rect 27721 22525 27755 22559
rect 31125 22525 31159 22559
rect 38209 22525 38243 22559
rect 27169 22457 27203 22491
rect 30573 22457 30607 22491
rect 33977 22457 34011 22491
rect 34713 22457 34747 22491
rect 3433 22389 3467 22423
rect 6745 22389 6779 22423
rect 11897 22389 11931 22423
rect 12706 22389 12740 22423
rect 14197 22389 14231 22423
rect 19073 22389 19107 22423
rect 24869 22389 24903 22423
rect 25329 22389 25363 22423
rect 30113 22389 30147 22423
rect 33241 22389 33275 22423
rect 34345 22389 34379 22423
rect 39681 22389 39715 22423
rect 14473 22185 14507 22219
rect 22845 22117 22879 22151
rect 28181 22117 28215 22151
rect 2053 22049 2087 22083
rect 4445 22049 4479 22083
rect 7297 22049 7331 22083
rect 9965 22049 9999 22083
rect 10609 22049 10643 22083
rect 13369 22049 13403 22083
rect 15669 22049 15703 22083
rect 17141 22049 17175 22083
rect 20821 22049 20855 22083
rect 23949 22049 23983 22083
rect 25145 22049 25179 22083
rect 27537 22049 27571 22083
rect 30757 22049 30791 22083
rect 1777 21981 1811 22015
rect 3985 21981 4019 22015
rect 7021 21981 7055 22015
rect 9689 21981 9723 22015
rect 10885 21981 10919 22015
rect 11621 21981 11655 22015
rect 12541 21981 12575 22015
rect 15393 21981 15427 22015
rect 20361 21981 20395 22015
rect 25789 21981 25823 22015
rect 28825 21981 28859 22015
rect 30573 21981 30607 22015
rect 32597 21981 32631 22015
rect 32873 21981 32907 22015
rect 49065 21981 49099 22015
rect 6193 21913 6227 21947
rect 9781 21913 9815 21947
rect 14381 21913 14415 21947
rect 17417 21913 17451 21947
rect 19497 21913 19531 21947
rect 23673 21913 23707 21947
rect 23765 21913 23799 21947
rect 24961 21913 24995 21947
rect 26065 21913 26099 21947
rect 31401 21913 31435 21947
rect 6285 21845 6319 21879
rect 9321 21845 9355 21879
rect 15025 21845 15059 21879
rect 18889 21845 18923 21879
rect 19625 21845 19659 21879
rect 23305 21845 23339 21879
rect 24593 21845 24627 21879
rect 25053 21845 25087 21879
rect 28641 21845 28675 21879
rect 30113 21845 30147 21879
rect 30481 21845 30515 21879
rect 31493 21845 31527 21879
rect 49249 21845 49283 21879
rect 11897 21641 11931 21675
rect 12357 21641 12391 21675
rect 25973 21641 26007 21675
rect 27721 21641 27755 21675
rect 32505 21641 32539 21675
rect 33057 21641 33091 21675
rect 5733 21573 5767 21607
rect 7389 21573 7423 21607
rect 12265 21573 12299 21607
rect 23673 21573 23707 21607
rect 31125 21573 31159 21607
rect 1777 21505 1811 21539
rect 3617 21505 3651 21539
rect 5641 21505 5675 21539
rect 6837 21505 6871 21539
rect 10241 21505 10275 21539
rect 10333 21505 10367 21539
rect 12817 21505 12851 21539
rect 15945 21505 15979 21539
rect 17233 21505 17267 21539
rect 21465 21505 21499 21539
rect 22385 21505 22419 21539
rect 22477 21505 22511 21539
rect 23397 21505 23431 21539
rect 26065 21505 26099 21539
rect 27629 21505 27663 21539
rect 31033 21505 31067 21539
rect 32413 21505 32447 21539
rect 33241 21505 33275 21539
rect 47961 21505 47995 21539
rect 2053 21437 2087 21471
rect 4169 21437 4203 21471
rect 5825 21437 5859 21471
rect 7113 21437 7147 21471
rect 10425 21437 10459 21471
rect 12449 21437 12483 21471
rect 13093 21437 13127 21471
rect 16037 21437 16071 21471
rect 16221 21437 16255 21471
rect 17693 21437 17727 21471
rect 18705 21437 18739 21471
rect 18981 21437 19015 21471
rect 22661 21437 22695 21471
rect 25145 21437 25179 21471
rect 26249 21437 26283 21471
rect 27813 21437 27847 21471
rect 28457 21437 28491 21471
rect 28733 21437 28767 21471
rect 31217 21437 31251 21471
rect 49157 21437 49191 21471
rect 8861 21369 8895 21403
rect 20453 21369 20487 21403
rect 22017 21369 22051 21403
rect 25605 21369 25639 21403
rect 5273 21301 5307 21335
rect 6929 21301 6963 21335
rect 9321 21301 9355 21335
rect 9873 21301 9907 21335
rect 14565 21301 14599 21335
rect 15393 21301 15427 21335
rect 15577 21301 15611 21335
rect 17049 21301 17083 21335
rect 27261 21301 27295 21335
rect 30205 21301 30239 21335
rect 30665 21301 30699 21335
rect 11437 21097 11471 21131
rect 14381 21097 14415 21131
rect 19704 21097 19738 21131
rect 21189 21097 21223 21131
rect 24685 21097 24719 21131
rect 32505 21097 32539 21131
rect 5365 21029 5399 21063
rect 7665 21029 7699 21063
rect 23305 21029 23339 21063
rect 4721 20961 4755 20995
rect 5825 20961 5859 20995
rect 8217 20961 8251 20995
rect 9597 20961 9631 20995
rect 12633 20961 12667 20995
rect 14841 20961 14875 20995
rect 15025 20961 15059 20995
rect 15669 20961 15703 20995
rect 15853 20961 15887 20995
rect 17601 20961 17635 20995
rect 18613 20961 18647 20995
rect 18797 20961 18831 20995
rect 19441 20961 19475 20995
rect 22109 20961 22143 20995
rect 23857 20961 23891 20995
rect 25145 20961 25179 20995
rect 25329 20961 25363 20995
rect 26065 20961 26099 20995
rect 30021 20961 30055 20995
rect 1777 20893 1811 20927
rect 5549 20893 5583 20927
rect 9321 20893 9355 20927
rect 12173 20893 12207 20927
rect 17325 20893 17359 20927
rect 22753 20893 22787 20927
rect 28273 20893 28307 20927
rect 28549 20893 28583 20927
rect 29745 20893 29779 20927
rect 31033 20893 31067 20927
rect 31309 20893 31343 20927
rect 2789 20825 2823 20859
rect 4537 20825 4571 20859
rect 8125 20825 8159 20859
rect 11345 20825 11379 20859
rect 21373 20825 21407 20859
rect 23765 20825 23799 20859
rect 25053 20825 25087 20859
rect 26341 20825 26375 20859
rect 32413 20825 32447 20859
rect 4169 20757 4203 20791
rect 4629 20757 4663 20791
rect 7297 20757 7331 20791
rect 8033 20757 8067 20791
rect 14749 20757 14783 20791
rect 15209 20757 15243 20791
rect 15577 20757 15611 20791
rect 16405 20757 16439 20791
rect 16957 20757 16991 20791
rect 17417 20757 17451 20791
rect 18153 20757 18187 20791
rect 18521 20757 18555 20791
rect 23673 20757 23707 20791
rect 27813 20757 27847 20791
rect 5641 20553 5675 20587
rect 11897 20553 11931 20587
rect 13001 20553 13035 20587
rect 17325 20553 17359 20587
rect 17417 20553 17451 20587
rect 21465 20553 21499 20587
rect 23489 20553 23523 20587
rect 23581 20553 23615 20587
rect 27629 20553 27663 20587
rect 30113 20553 30147 20587
rect 31033 20553 31067 20587
rect 12909 20485 12943 20519
rect 18613 20485 18647 20519
rect 22109 20485 22143 20519
rect 1777 20417 1811 20451
rect 3617 20417 3651 20451
rect 6561 20417 6595 20451
rect 8401 20417 8435 20451
rect 10701 20417 10735 20451
rect 11805 20417 11839 20451
rect 16037 20417 16071 20451
rect 18521 20417 18555 20451
rect 19717 20417 19751 20451
rect 24317 20417 24351 20451
rect 27537 20417 27571 20451
rect 28365 20417 28399 20451
rect 30941 20417 30975 20451
rect 2789 20349 2823 20383
rect 3893 20349 3927 20383
rect 5733 20349 5767 20383
rect 5825 20349 5859 20383
rect 7021 20349 7055 20383
rect 8677 20349 8711 20383
rect 13185 20349 13219 20383
rect 13737 20349 13771 20383
rect 14013 20349 14047 20383
rect 17601 20349 17635 20383
rect 18797 20349 18831 20383
rect 19993 20349 20027 20383
rect 23765 20349 23799 20383
rect 24593 20349 24627 20383
rect 27721 20349 27755 20383
rect 28641 20349 28675 20383
rect 31125 20349 31159 20383
rect 5273 20281 5307 20315
rect 10885 20281 10919 20315
rect 12541 20281 12575 20315
rect 23121 20281 23155 20315
rect 26065 20281 26099 20315
rect 10149 20213 10183 20247
rect 15485 20213 15519 20247
rect 16129 20213 16163 20247
rect 16957 20213 16991 20247
rect 18153 20213 18187 20247
rect 22201 20213 22235 20247
rect 27169 20213 27203 20247
rect 30573 20213 30607 20247
rect 6285 20009 6319 20043
rect 7008 20009 7042 20043
rect 11713 20009 11747 20043
rect 16313 20009 16347 20043
rect 16957 20009 16991 20043
rect 23305 20009 23339 20043
rect 27629 20009 27663 20043
rect 22017 19941 22051 19975
rect 22845 19941 22879 19975
rect 24685 19941 24719 19975
rect 2053 19873 2087 19907
rect 4537 19873 4571 19907
rect 6745 19873 6779 19907
rect 9965 19873 9999 19907
rect 13645 19873 13679 19907
rect 14841 19873 14875 19907
rect 17417 19873 17451 19907
rect 17601 19873 17635 19907
rect 18705 19873 18739 19907
rect 20269 19873 20303 19907
rect 20545 19873 20579 19907
rect 23857 19873 23891 19907
rect 25329 19873 25363 19907
rect 28365 19873 28399 19907
rect 29745 19873 29779 19907
rect 31585 19873 31619 19907
rect 1777 19805 1811 19839
rect 14565 19805 14599 19839
rect 17325 19805 17359 19839
rect 19625 19805 19659 19839
rect 23765 19805 23799 19839
rect 25881 19805 25915 19839
rect 30021 19805 30055 19839
rect 4813 19737 4847 19771
rect 9321 19737 9355 19771
rect 10241 19737 10275 19771
rect 12265 19737 12299 19771
rect 13369 19737 13403 19771
rect 25053 19737 25087 19771
rect 26157 19737 26191 19771
rect 31493 19737 31527 19771
rect 8493 19669 8527 19703
rect 9413 19669 9447 19703
rect 12357 19669 12391 19703
rect 13001 19669 13035 19703
rect 13461 19669 13495 19703
rect 18153 19669 18187 19703
rect 18521 19669 18555 19703
rect 18613 19669 18647 19703
rect 19717 19669 19751 19703
rect 23673 19669 23707 19703
rect 25145 19669 25179 19703
rect 28595 19669 28629 19703
rect 31033 19669 31067 19703
rect 31401 19669 31435 19703
rect 5733 19465 5767 19499
rect 8769 19465 8803 19499
rect 21465 19465 21499 19499
rect 22477 19465 22511 19499
rect 22845 19465 22879 19499
rect 22937 19465 22971 19499
rect 23673 19465 23707 19499
rect 24041 19465 24075 19499
rect 27629 19465 27663 19499
rect 4537 19397 4571 19431
rect 10149 19397 10183 19431
rect 14657 19397 14691 19431
rect 15761 19397 15795 19431
rect 1777 19329 1811 19363
rect 3617 19329 3651 19363
rect 5641 19329 5675 19363
rect 7028 19329 7062 19363
rect 9229 19329 9263 19363
rect 11713 19329 11747 19363
rect 13921 19329 13955 19363
rect 15669 19329 15703 19363
rect 17233 19329 17267 19363
rect 17325 19329 17359 19363
rect 18521 19329 18555 19363
rect 24133 19329 24167 19363
rect 25053 19329 25087 19363
rect 27813 19329 27847 19363
rect 2053 19261 2087 19295
rect 5825 19261 5859 19295
rect 7297 19261 7331 19295
rect 11989 19261 12023 19295
rect 15853 19261 15887 19295
rect 17509 19261 17543 19295
rect 18613 19261 18647 19295
rect 18797 19261 18831 19295
rect 19717 19261 19751 19295
rect 19993 19261 20027 19295
rect 23121 19261 23155 19295
rect 24317 19261 24351 19295
rect 25881 19261 25915 19295
rect 26617 19261 26651 19295
rect 28365 19261 28399 19295
rect 28641 19261 28675 19295
rect 5273 19125 5307 19159
rect 13461 19125 13495 19159
rect 15301 19125 15335 19159
rect 16865 19125 16899 19159
rect 18153 19125 18187 19159
rect 30113 19125 30147 19159
rect 12081 18921 12115 18955
rect 22937 18921 22971 18955
rect 24777 18921 24811 18955
rect 27169 18921 27203 18955
rect 28825 18921 28859 18955
rect 14657 18853 14691 18887
rect 17877 18853 17911 18887
rect 23397 18853 23431 18887
rect 29745 18853 29779 18887
rect 31033 18853 31067 18887
rect 6561 18785 6595 18819
rect 7481 18785 7515 18819
rect 9689 18785 9723 18819
rect 11437 18785 11471 18819
rect 12633 18785 12667 18819
rect 15117 18785 15151 18819
rect 18429 18785 18463 18819
rect 20453 18785 20487 18819
rect 21189 18785 21223 18819
rect 21465 18785 21499 18819
rect 25421 18785 25455 18819
rect 28181 18785 28215 18819
rect 30297 18785 30331 18819
rect 1777 18717 1811 18751
rect 4353 18717 4387 18751
rect 4813 18717 4847 18751
rect 7205 18717 7239 18751
rect 9505 18717 9539 18751
rect 13369 18717 13403 18751
rect 14473 18717 14507 18751
rect 18245 18717 18279 18751
rect 23581 18717 23615 18751
rect 29009 18717 29043 18751
rect 30113 18717 30147 18751
rect 2513 18649 2547 18683
rect 5089 18649 5123 18683
rect 10425 18649 10459 18683
rect 11253 18649 11287 18683
rect 13553 18649 13587 18683
rect 15393 18649 15427 18683
rect 19717 18649 19751 18683
rect 25697 18649 25731 18683
rect 28089 18649 28123 18683
rect 4169 18581 4203 18615
rect 9137 18581 9171 18615
rect 9597 18581 9631 18615
rect 10885 18581 10919 18615
rect 11345 18581 11379 18615
rect 12449 18581 12483 18615
rect 12541 18581 12575 18615
rect 16865 18581 16899 18615
rect 18337 18581 18371 18615
rect 27629 18581 27663 18615
rect 27997 18581 28031 18615
rect 30205 18581 30239 18615
rect 5733 18377 5767 18411
rect 10885 18377 10919 18411
rect 15117 18377 15151 18411
rect 15577 18377 15611 18411
rect 19717 18377 19751 18411
rect 20085 18377 20119 18411
rect 24869 18377 24903 18411
rect 30297 18377 30331 18411
rect 30757 18377 30791 18411
rect 8585 18309 8619 18343
rect 13737 18309 13771 18343
rect 14565 18309 14599 18343
rect 17417 18309 17451 18343
rect 22477 18309 22511 18343
rect 25329 18309 25363 18343
rect 26065 18309 26099 18343
rect 30665 18309 30699 18343
rect 1777 18241 1811 18275
rect 3433 18241 3467 18275
rect 5641 18241 5675 18275
rect 6561 18241 6595 18275
rect 10793 18241 10827 18275
rect 12449 18241 12483 18275
rect 12541 18241 12575 18275
rect 15485 18241 15519 18275
rect 17233 18241 17267 18275
rect 18705 18241 18739 18275
rect 22017 18241 22051 18275
rect 22569 18241 22603 18275
rect 27353 18241 27387 18275
rect 28089 18241 28123 18275
rect 2789 18173 2823 18207
rect 3893 18173 3927 18207
rect 5917 18173 5951 18207
rect 7021 18173 7055 18207
rect 9321 18173 9355 18207
rect 10977 18173 11011 18207
rect 12725 18173 12759 18207
rect 15761 18173 15795 18207
rect 18429 18173 18463 18207
rect 20177 18173 20211 18207
rect 20269 18173 20303 18207
rect 22661 18173 22695 18207
rect 23121 18173 23155 18207
rect 23397 18173 23431 18207
rect 28365 18173 28399 18207
rect 30849 18173 30883 18207
rect 10425 18105 10459 18139
rect 13277 18105 13311 18139
rect 5273 18037 5307 18071
rect 12081 18037 12115 18071
rect 21465 18037 21499 18071
rect 22109 18037 22143 18071
rect 29837 18037 29871 18071
rect 4353 17833 4387 17867
rect 6653 17833 6687 17867
rect 7297 17833 7331 17867
rect 14473 17833 14507 17867
rect 15025 17833 15059 17867
rect 19441 17833 19475 17867
rect 26617 17833 26651 17867
rect 26972 17833 27006 17867
rect 29745 17833 29779 17867
rect 7849 17765 7883 17799
rect 10609 17765 10643 17799
rect 13737 17765 13771 17799
rect 20729 17765 20763 17799
rect 2053 17697 2087 17731
rect 8493 17697 8527 17731
rect 9873 17697 9907 17731
rect 11161 17697 11195 17731
rect 12265 17697 12299 17731
rect 16313 17697 16347 17731
rect 16589 17697 16623 17731
rect 21281 17697 21315 17731
rect 22569 17697 22603 17731
rect 24869 17697 24903 17731
rect 26709 17697 26743 17731
rect 30297 17697 30331 17731
rect 1777 17629 1811 17663
rect 4905 17629 4939 17663
rect 8217 17629 8251 17663
rect 9137 17629 9171 17663
rect 11989 17629 12023 17663
rect 15209 17629 15243 17663
rect 15853 17629 15887 17663
rect 18889 17629 18923 17663
rect 19625 17629 19659 17663
rect 20545 17629 20579 17663
rect 22293 17629 22327 17663
rect 29009 17629 29043 17663
rect 30113 17629 30147 17663
rect 4261 17561 4295 17595
rect 5181 17561 5215 17595
rect 7205 17561 7239 17595
rect 10977 17561 11011 17595
rect 14381 17561 14415 17595
rect 25145 17561 25179 17595
rect 8309 17493 8343 17527
rect 11069 17493 11103 17527
rect 15669 17493 15703 17527
rect 18061 17493 18095 17527
rect 18705 17493 18739 17527
rect 20177 17493 20211 17527
rect 21097 17493 21131 17527
rect 21189 17493 21223 17527
rect 24041 17493 24075 17527
rect 28457 17493 28491 17527
rect 30205 17493 30239 17527
rect 30941 17493 30975 17527
rect 6837 17289 6871 17323
rect 7205 17289 7239 17323
rect 7297 17289 7331 17323
rect 8033 17289 8067 17323
rect 9689 17289 9723 17323
rect 10793 17289 10827 17323
rect 12541 17289 12575 17323
rect 13001 17289 13035 17323
rect 20729 17289 20763 17323
rect 21097 17289 21131 17323
rect 21925 17289 21959 17323
rect 26525 17289 26559 17323
rect 5733 17221 5767 17255
rect 8493 17221 8527 17255
rect 9597 17221 9631 17255
rect 14749 17221 14783 17255
rect 21189 17221 21223 17255
rect 1777 17153 1811 17187
rect 3433 17153 3467 17187
rect 5641 17153 5675 17187
rect 8401 17153 8435 17187
rect 11805 17153 11839 17187
rect 12909 17153 12943 17187
rect 14657 17153 14691 17187
rect 17233 17153 17267 17187
rect 22293 17153 22327 17187
rect 22385 17153 22419 17187
rect 23673 17153 23707 17187
rect 24501 17153 24535 17187
rect 24777 17153 24811 17187
rect 27905 17153 27939 17187
rect 2053 17085 2087 17119
rect 3893 17085 3927 17119
rect 5917 17085 5951 17119
rect 7481 17085 7515 17119
rect 8585 17085 8619 17119
rect 9781 17085 9815 17119
rect 10885 17085 10919 17119
rect 10977 17085 11011 17119
rect 13185 17085 13219 17119
rect 14841 17085 14875 17119
rect 17325 17085 17359 17119
rect 17509 17085 17543 17119
rect 18153 17085 18187 17119
rect 18429 17085 18463 17119
rect 19901 17085 19935 17119
rect 21281 17085 21315 17119
rect 22477 17085 22511 17119
rect 23765 17085 23799 17119
rect 23857 17085 23891 17119
rect 25053 17085 25087 17119
rect 28181 17085 28215 17119
rect 11989 17017 12023 17051
rect 23305 17017 23339 17051
rect 5273 16949 5307 16983
rect 9229 16949 9263 16983
rect 10425 16949 10459 16983
rect 14289 16949 14323 16983
rect 15853 16949 15887 16983
rect 16865 16949 16899 16983
rect 23121 16949 23155 16983
rect 27445 16949 27479 16983
rect 29653 16949 29687 16983
rect 16865 16745 16899 16779
rect 18797 16745 18831 16779
rect 10057 16677 10091 16711
rect 10149 16677 10183 16711
rect 13001 16677 13035 16711
rect 22661 16677 22695 16711
rect 7113 16609 7147 16643
rect 7205 16609 7239 16643
rect 8401 16609 8435 16643
rect 10701 16609 10735 16643
rect 12265 16609 12299 16643
rect 12449 16609 12483 16643
rect 13461 16609 13495 16643
rect 13645 16609 13679 16643
rect 14565 16609 14599 16643
rect 15669 16609 15703 16643
rect 19717 16609 19751 16643
rect 23765 16609 23799 16643
rect 25145 16609 25179 16643
rect 25329 16609 25363 16643
rect 27077 16609 27111 16643
rect 27261 16609 27295 16643
rect 28457 16609 28491 16643
rect 1777 16541 1811 16575
rect 4077 16541 4111 16575
rect 6101 16541 6135 16575
rect 8217 16541 8251 16575
rect 9689 16541 9723 16575
rect 9873 16541 9907 16575
rect 10609 16541 10643 16575
rect 17509 16541 17543 16575
rect 18153 16541 18187 16575
rect 19441 16541 19475 16575
rect 23581 16541 23615 16575
rect 26985 16541 27019 16575
rect 28181 16541 28215 16575
rect 2513 16473 2547 16507
rect 4905 16473 4939 16507
rect 5917 16473 5951 16507
rect 8309 16473 8343 16507
rect 21465 16473 21499 16507
rect 25053 16473 25087 16507
rect 28273 16473 28307 16507
rect 6653 16405 6687 16439
rect 7021 16405 7055 16439
rect 7849 16405 7883 16439
rect 10517 16405 10551 16439
rect 11805 16405 11839 16439
rect 12173 16405 12207 16439
rect 13369 16405 13403 16439
rect 15025 16405 15059 16439
rect 15393 16405 15427 16439
rect 15485 16405 15519 16439
rect 17325 16405 17359 16439
rect 17969 16405 18003 16439
rect 23213 16405 23247 16439
rect 23673 16405 23707 16439
rect 24685 16405 24719 16439
rect 26617 16405 26651 16439
rect 27813 16405 27847 16439
rect 5641 16201 5675 16235
rect 7297 16201 7331 16235
rect 13829 16201 13863 16235
rect 14841 16201 14875 16235
rect 17785 16201 17819 16235
rect 17877 16201 17911 16235
rect 21097 16201 21131 16235
rect 22201 16201 22235 16235
rect 22845 16201 22879 16235
rect 23673 16201 23707 16235
rect 23765 16201 23799 16235
rect 26617 16201 26651 16235
rect 4353 16133 4387 16167
rect 6837 16133 6871 16167
rect 8769 16133 8803 16167
rect 1777 16065 1811 16099
rect 3617 16065 3651 16099
rect 5733 16065 5767 16099
rect 6653 16065 6687 16099
rect 7665 16065 7699 16099
rect 8493 16065 8527 16099
rect 11161 16065 11195 16099
rect 12081 16065 12115 16099
rect 16313 16065 16347 16099
rect 18797 16065 18831 16099
rect 19165 16065 19199 16099
rect 20177 16065 20211 16099
rect 21189 16065 21223 16099
rect 24869 16065 24903 16099
rect 2053 15997 2087 16031
rect 5917 15997 5951 16031
rect 7757 15997 7791 16031
rect 7849 15997 7883 16031
rect 10241 15997 10275 16031
rect 12357 15997 12391 16031
rect 14933 15997 14967 16031
rect 15025 15997 15059 16031
rect 17969 15997 18003 16031
rect 18889 15997 18923 16031
rect 21373 15997 21407 16031
rect 23857 15997 23891 16031
rect 25145 15997 25179 16031
rect 23305 15929 23339 15963
rect 5273 15861 5307 15895
rect 10977 15861 11011 15895
rect 14473 15861 14507 15895
rect 16129 15861 16163 15895
rect 17417 15861 17451 15895
rect 20729 15861 20763 15895
rect 3985 15657 4019 15691
rect 7849 15657 7883 15691
rect 9321 15657 9355 15691
rect 12081 15657 12115 15691
rect 19441 15657 19475 15691
rect 10241 15589 10275 15623
rect 10885 15589 10919 15623
rect 13553 15589 13587 15623
rect 14749 15589 14783 15623
rect 15945 15589 15979 15623
rect 23029 15589 23063 15623
rect 2053 15521 2087 15555
rect 4445 15521 4479 15555
rect 4629 15521 4663 15555
rect 5733 15521 5767 15555
rect 7021 15521 7055 15555
rect 8493 15521 8527 15555
rect 11437 15521 11471 15555
rect 12725 15521 12759 15555
rect 15301 15521 15335 15555
rect 16405 15521 16439 15555
rect 16589 15521 16623 15555
rect 17417 15521 17451 15555
rect 19717 15521 19751 15555
rect 22477 15521 22511 15555
rect 22661 15521 22695 15555
rect 25789 15521 25823 15555
rect 1777 15453 1811 15487
rect 8309 15453 8343 15487
rect 10425 15453 10459 15487
rect 11253 15453 11287 15487
rect 12541 15453 12575 15487
rect 13737 15453 13771 15487
rect 17141 15453 17175 15487
rect 19625 15453 19659 15487
rect 22385 15453 22419 15487
rect 23121 15453 23155 15487
rect 25605 15453 25639 15487
rect 5641 15385 5675 15419
rect 6837 15385 6871 15419
rect 9229 15385 9263 15419
rect 11345 15385 11379 15419
rect 15209 15385 15243 15419
rect 19993 15385 20027 15419
rect 23949 15385 23983 15419
rect 25697 15385 25731 15419
rect 4353 15317 4387 15351
rect 5181 15317 5215 15351
rect 5549 15317 5583 15351
rect 6377 15317 6411 15351
rect 6745 15317 6779 15351
rect 8217 15317 8251 15351
rect 12449 15317 12483 15351
rect 15117 15317 15151 15351
rect 16313 15317 16347 15351
rect 18889 15317 18923 15351
rect 21465 15317 21499 15351
rect 22017 15317 22051 15351
rect 25237 15317 25271 15351
rect 6745 15113 6779 15147
rect 7757 15113 7791 15147
rect 9229 15113 9263 15147
rect 13001 15113 13035 15147
rect 19441 15113 19475 15147
rect 4445 15045 4479 15079
rect 10793 15045 10827 15079
rect 10885 15045 10919 15079
rect 13369 15045 13403 15079
rect 19809 15045 19843 15079
rect 19901 15045 19935 15079
rect 25145 15045 25179 15079
rect 1777 14977 1811 15011
rect 4169 14977 4203 15011
rect 6653 14977 6687 15011
rect 9597 14977 9631 15011
rect 11989 14977 12023 15011
rect 17141 14977 17175 15011
rect 20637 14977 20671 15011
rect 20913 14977 20947 15011
rect 22017 14977 22051 15011
rect 24869 14977 24903 15011
rect 2053 14909 2087 14943
rect 7849 14909 7883 14943
rect 7941 14909 7975 14943
rect 8769 14909 8803 14943
rect 9689 14909 9723 14943
rect 9781 14909 9815 14943
rect 10977 14909 11011 14943
rect 11713 14909 11747 14943
rect 13461 14909 13495 14943
rect 13553 14909 13587 14943
rect 14565 14909 14599 14943
rect 14841 14909 14875 14943
rect 16313 14909 16347 14943
rect 18889 14909 18923 14943
rect 20085 14909 20119 14943
rect 23765 14909 23799 14943
rect 5917 14841 5951 14875
rect 10425 14841 10459 14875
rect 3709 14773 3743 14807
rect 7389 14773 7423 14807
rect 22280 14773 22314 14807
rect 26617 14773 26651 14807
rect 3985 14569 4019 14603
rect 9413 14569 9447 14603
rect 18613 14569 18647 14603
rect 13737 14501 13771 14535
rect 2053 14433 2087 14467
rect 4537 14433 4571 14467
rect 5549 14433 5583 14467
rect 8401 14433 8435 14467
rect 10057 14433 10091 14467
rect 11161 14433 11195 14467
rect 12265 14433 12299 14467
rect 14933 14433 14967 14467
rect 19717 14433 19751 14467
rect 21281 14433 21315 14467
rect 22293 14433 22327 14467
rect 25145 14433 25179 14467
rect 26341 14433 26375 14467
rect 1777 14365 1811 14399
rect 5273 14365 5307 14399
rect 7297 14365 7331 14399
rect 8217 14365 8251 14399
rect 8309 14365 8343 14399
rect 9873 14365 9907 14399
rect 10977 14365 11011 14399
rect 11989 14365 12023 14399
rect 14657 14365 14691 14399
rect 16865 14365 16899 14399
rect 19441 14365 19475 14399
rect 21097 14365 21131 14399
rect 24961 14365 24995 14399
rect 26249 14365 26283 14399
rect 4445 14297 4479 14331
rect 17141 14297 17175 14331
rect 22569 14297 22603 14331
rect 26157 14297 26191 14331
rect 4353 14229 4387 14263
rect 7849 14229 7883 14263
rect 9781 14229 9815 14263
rect 10609 14229 10643 14263
rect 11069 14229 11103 14263
rect 16405 14229 16439 14263
rect 20729 14229 20763 14263
rect 21189 14229 21223 14263
rect 24041 14229 24075 14263
rect 24593 14229 24627 14263
rect 25053 14229 25087 14263
rect 25789 14229 25823 14263
rect 5273 14025 5307 14059
rect 5641 14025 5675 14059
rect 6929 14025 6963 14059
rect 7297 14025 7331 14059
rect 8585 14025 8619 14059
rect 11989 14025 12023 14059
rect 14749 14025 14783 14059
rect 14841 14025 14875 14059
rect 15577 14025 15611 14059
rect 18889 14025 18923 14059
rect 20177 14025 20211 14059
rect 23397 14025 23431 14059
rect 24593 14025 24627 14059
rect 24961 14025 24995 14059
rect 8493 13957 8527 13991
rect 9597 13957 9631 13991
rect 12357 13957 12391 13991
rect 13645 13957 13679 13991
rect 17417 13957 17451 13991
rect 22569 13957 22603 13991
rect 22661 13957 22695 13991
rect 25053 13957 25087 13991
rect 2973 13889 3007 13923
rect 3433 13889 3467 13923
rect 3709 13889 3743 13923
rect 7389 13889 7423 13923
rect 12449 13889 12483 13923
rect 13553 13889 13587 13923
rect 15945 13889 15979 13923
rect 19625 13889 19659 13923
rect 20545 13889 20579 13923
rect 20637 13889 20671 13923
rect 23765 13889 23799 13923
rect 23857 13889 23891 13923
rect 5733 13821 5767 13855
rect 5825 13821 5859 13855
rect 7573 13821 7607 13855
rect 8677 13821 8711 13855
rect 9321 13821 9355 13855
rect 11069 13821 11103 13855
rect 12633 13821 12667 13855
rect 13829 13821 13863 13855
rect 15025 13821 15059 13855
rect 16037 13821 16071 13855
rect 16129 13821 16163 13855
rect 17141 13821 17175 13855
rect 20821 13821 20855 13855
rect 22753 13821 22787 13855
rect 23949 13821 23983 13855
rect 25145 13821 25179 13855
rect 13185 13753 13219 13787
rect 14381 13753 14415 13787
rect 19441 13753 19475 13787
rect 8125 13685 8159 13719
rect 22201 13685 22235 13719
rect 13737 13481 13771 13515
rect 18889 13481 18923 13515
rect 22845 13481 22879 13515
rect 8493 13413 8527 13447
rect 16037 13413 16071 13447
rect 22109 13413 22143 13447
rect 2789 13345 2823 13379
rect 4169 13345 4203 13379
rect 6745 13345 6779 13379
rect 10793 13345 10827 13379
rect 11989 13345 12023 13379
rect 14289 13345 14323 13379
rect 17141 13345 17175 13379
rect 20361 13345 20395 13379
rect 23305 13345 23339 13379
rect 23489 13345 23523 13379
rect 1777 13277 1811 13311
rect 9781 13277 9815 13311
rect 16681 13277 16715 13311
rect 19625 13277 19659 13311
rect 4445 13209 4479 13243
rect 7021 13209 7055 13243
rect 10609 13209 10643 13243
rect 12265 13209 12299 13243
rect 14565 13209 14599 13243
rect 17417 13209 17451 13243
rect 20637 13209 20671 13243
rect 23213 13209 23247 13243
rect 24593 13209 24627 13243
rect 25421 13209 25455 13243
rect 5917 13141 5951 13175
rect 9597 13141 9631 13175
rect 10241 13141 10275 13175
rect 10701 13141 10735 13175
rect 16497 13141 16531 13175
rect 19441 13141 19475 13175
rect 3525 12937 3559 12971
rect 4077 12937 4111 12971
rect 7389 12937 7423 12971
rect 7481 12937 7515 12971
rect 12633 12937 12667 12971
rect 13001 12937 13035 12971
rect 13093 12937 13127 12971
rect 17969 12937 18003 12971
rect 18337 12937 18371 12971
rect 24777 12937 24811 12971
rect 2789 12869 2823 12903
rect 3433 12869 3467 12903
rect 4445 12869 4479 12903
rect 8493 12869 8527 12903
rect 10241 12869 10275 12903
rect 14289 12869 14323 12903
rect 15025 12869 15059 12903
rect 19165 12869 19199 12903
rect 21097 12869 21131 12903
rect 1777 12801 1811 12835
rect 5641 12801 5675 12835
rect 5733 12801 5767 12835
rect 8217 12801 8251 12835
rect 11161 12801 11195 12835
rect 14197 12801 14231 12835
rect 18429 12801 18463 12835
rect 23029 12801 23063 12835
rect 4537 12733 4571 12767
rect 4721 12733 4755 12767
rect 5917 12733 5951 12767
rect 7665 12733 7699 12767
rect 13277 12733 13311 12767
rect 14473 12733 14507 12767
rect 15853 12733 15887 12767
rect 18613 12733 18647 12767
rect 19993 12733 20027 12767
rect 21189 12733 21223 12767
rect 21373 12733 21407 12767
rect 23305 12733 23339 12767
rect 7021 12665 7055 12699
rect 12173 12665 12207 12699
rect 5273 12597 5307 12631
rect 13829 12597 13863 12631
rect 17049 12597 17083 12631
rect 20729 12597 20763 12631
rect 4077 12393 4111 12427
rect 7849 12393 7883 12427
rect 11805 12393 11839 12427
rect 13001 12393 13035 12427
rect 18061 12393 18095 12427
rect 21833 12393 21867 12427
rect 3433 12325 3467 12359
rect 1593 12257 1627 12291
rect 1869 12257 1903 12291
rect 4721 12257 4755 12291
rect 7389 12257 7423 12291
rect 8309 12257 8343 12291
rect 8493 12257 8527 12291
rect 9873 12257 9907 12291
rect 10793 12257 10827 12291
rect 12357 12257 12391 12291
rect 13645 12257 13679 12291
rect 16313 12257 16347 12291
rect 20085 12257 20119 12291
rect 22569 12257 22603 12291
rect 2605 12189 2639 12223
rect 3249 12189 3283 12223
rect 4445 12189 4479 12223
rect 5365 12189 5399 12223
rect 8217 12189 8251 12223
rect 9137 12189 9171 12223
rect 10517 12189 10551 12223
rect 12265 12189 12299 12223
rect 22293 12189 22327 12223
rect 2789 12121 2823 12155
rect 4537 12121 4571 12155
rect 5641 12121 5675 12155
rect 14381 12121 14415 12155
rect 15117 12121 15151 12155
rect 16589 12121 16623 12155
rect 20361 12121 20395 12155
rect 12173 12053 12207 12087
rect 13369 12053 13403 12087
rect 13461 12053 13495 12087
rect 24041 12053 24075 12087
rect 1777 11849 1811 11883
rect 4445 11849 4479 11883
rect 6561 11849 6595 11883
rect 9137 11849 9171 11883
rect 11989 11849 12023 11883
rect 14933 11849 14967 11883
rect 15577 11849 15611 11883
rect 17417 11849 17451 11883
rect 18153 11849 18187 11883
rect 18521 11849 18555 11883
rect 18613 11849 18647 11883
rect 24133 11849 24167 11883
rect 7665 11781 7699 11815
rect 9597 11781 9631 11815
rect 16037 11781 16071 11815
rect 22661 11781 22695 11815
rect 1961 11713 1995 11747
rect 2145 11713 2179 11747
rect 2421 11713 2455 11747
rect 4353 11713 4387 11747
rect 5457 11713 5491 11747
rect 6745 11713 6779 11747
rect 11161 11713 11195 11747
rect 12357 11713 12391 11747
rect 15945 11713 15979 11747
rect 17325 11713 17359 11747
rect 4629 11645 4663 11679
rect 5181 11645 5215 11679
rect 7297 11645 7331 11679
rect 7389 11645 7423 11679
rect 10333 11645 10367 11679
rect 12449 11645 12483 11679
rect 12541 11645 12575 11679
rect 13185 11645 13219 11679
rect 13461 11645 13495 11679
rect 16221 11645 16255 11679
rect 17509 11645 17543 11679
rect 18705 11645 18739 11679
rect 19717 11645 19751 11679
rect 19993 11645 20027 11679
rect 22385 11645 22419 11679
rect 16957 11577 16991 11611
rect 3985 11509 4019 11543
rect 21465 11509 21499 11543
rect 2145 11305 2179 11339
rect 2605 11305 2639 11339
rect 6561 11305 6595 11339
rect 7389 11305 7423 11339
rect 7849 11305 7883 11339
rect 10333 11305 10367 11339
rect 13277 11305 13311 11339
rect 16497 11305 16531 11339
rect 17398 11305 17432 11339
rect 18889 11305 18923 11339
rect 3985 11237 4019 11271
rect 9137 11237 9171 11271
rect 2789 11169 2823 11203
rect 4813 11169 4847 11203
rect 5089 11169 5123 11203
rect 8309 11169 8343 11203
rect 8493 11169 8527 11203
rect 9689 11169 9723 11203
rect 10977 11169 11011 11203
rect 11529 11169 11563 11203
rect 11805 11169 11839 11203
rect 14749 11169 14783 11203
rect 22661 11169 22695 11203
rect 29745 11169 29779 11203
rect 3065 11101 3099 11135
rect 4169 11101 4203 11135
rect 8217 11101 8251 11135
rect 9505 11101 9539 11135
rect 9597 11101 9631 11135
rect 17141 11101 17175 11135
rect 19533 11101 19567 11135
rect 20913 11101 20947 11135
rect 10701 11033 10735 11067
rect 10793 11033 10827 11067
rect 15025 11033 15059 11067
rect 20269 11033 20303 11067
rect 21189 11033 21223 11067
rect 30021 11033 30055 11067
rect 31769 11033 31803 11067
rect 3893 10761 3927 10795
rect 5273 10761 5307 10795
rect 10333 10761 10367 10795
rect 13829 10761 13863 10795
rect 14381 10761 14415 10795
rect 15945 10761 15979 10795
rect 19257 10761 19291 10795
rect 4721 10693 4755 10727
rect 9413 10693 9447 10727
rect 14749 10693 14783 10727
rect 2053 10625 2087 10659
rect 2329 10625 2363 10659
rect 3801 10625 3835 10659
rect 4537 10625 4571 10659
rect 5641 10625 5675 10659
rect 6929 10625 6963 10659
rect 10701 10625 10735 10659
rect 12081 10625 12115 10659
rect 17049 10625 17083 10659
rect 17509 10625 17543 10659
rect 5733 10557 5767 10591
rect 5917 10557 5951 10591
rect 7389 10557 7423 10591
rect 7665 10557 7699 10591
rect 10793 10557 10827 10591
rect 10977 10557 11011 10591
rect 14841 10557 14875 10591
rect 14933 10557 14967 10591
rect 16037 10557 16071 10591
rect 16221 10557 16255 10591
rect 17785 10557 17819 10591
rect 19717 10557 19751 10591
rect 19993 10557 20027 10591
rect 15577 10489 15611 10523
rect 6745 10421 6779 10455
rect 12338 10421 12372 10455
rect 21465 10421 21499 10455
rect 6009 10217 6043 10251
rect 9597 10217 9631 10251
rect 13645 10217 13679 10251
rect 16313 10217 16347 10251
rect 18889 10217 18923 10251
rect 1593 10081 1627 10115
rect 1869 10081 1903 10115
rect 4813 10081 4847 10115
rect 6837 10081 6871 10115
rect 10517 10081 10551 10115
rect 10609 10081 10643 10115
rect 11253 10081 11287 10115
rect 11529 10081 11563 10115
rect 13001 10081 13035 10115
rect 14565 10081 14599 10115
rect 14841 10081 14875 10115
rect 19441 10081 19475 10115
rect 3065 10013 3099 10047
rect 4537 10013 4571 10047
rect 10425 10013 10459 10047
rect 17141 10013 17175 10047
rect 7113 9945 7147 9979
rect 17417 9945 17451 9979
rect 19717 9945 19751 9979
rect 21649 9945 21683 9979
rect 2881 9877 2915 9911
rect 8585 9877 8619 9911
rect 10057 9877 10091 9911
rect 21189 9877 21223 9911
rect 6929 9673 6963 9707
rect 10333 9673 10367 9707
rect 13461 9673 13495 9707
rect 4905 9605 4939 9639
rect 8401 9605 8435 9639
rect 10793 9605 10827 9639
rect 19533 9605 19567 9639
rect 1593 9537 1627 9571
rect 3341 9537 3375 9571
rect 4353 9537 4387 9571
rect 5365 9537 5399 9571
rect 6009 9537 6043 9571
rect 7297 9537 7331 9571
rect 10701 9537 10735 9571
rect 11713 9537 11747 9571
rect 14473 9537 14507 9571
rect 19441 9537 19475 9571
rect 27537 9537 27571 9571
rect 1869 9469 1903 9503
rect 7389 9469 7423 9503
rect 7481 9469 7515 9503
rect 8125 9469 8159 9503
rect 10977 9469 11011 9503
rect 11989 9469 12023 9503
rect 14749 9469 14783 9503
rect 16221 9469 16255 9503
rect 16865 9469 16899 9503
rect 17141 9469 17175 9503
rect 19717 9469 19751 9503
rect 27997 9469 28031 9503
rect 3157 9401 3191 9435
rect 19073 9401 19107 9435
rect 3065 9333 3099 9367
rect 3709 9333 3743 9367
rect 9873 9333 9907 9367
rect 18613 9333 18647 9367
rect 27813 9333 27847 9367
rect 3985 9129 4019 9163
rect 4997 9129 5031 9163
rect 5181 9129 5215 9163
rect 6837 9129 6871 9163
rect 6193 9061 6227 9095
rect 10425 9061 10459 9095
rect 12817 9061 12851 9095
rect 17785 9061 17819 9095
rect 1869 8993 1903 9027
rect 5733 8993 5767 9027
rect 7757 8993 7791 9027
rect 9137 8993 9171 9027
rect 9413 8993 9447 9027
rect 10977 8993 11011 9027
rect 12265 8993 12299 9027
rect 14749 8993 14783 9027
rect 14933 8993 14967 9027
rect 16037 8993 16071 9027
rect 1593 8925 1627 8959
rect 3065 8925 3099 8959
rect 4169 8925 4203 8959
rect 5365 8925 5399 8959
rect 6377 8925 6411 8959
rect 7021 8925 7055 8959
rect 7481 8925 7515 8959
rect 10885 8925 10919 8959
rect 13001 8925 13035 8959
rect 13737 8925 13771 8959
rect 14657 8925 14691 8959
rect 16313 8857 16347 8891
rect 2881 8789 2915 8823
rect 10793 8789 10827 8823
rect 11621 8789 11655 8823
rect 11989 8789 12023 8823
rect 12081 8789 12115 8823
rect 14289 8789 14323 8823
rect 5825 8585 5859 8619
rect 11897 8585 11931 8619
rect 13093 8585 13127 8619
rect 14749 8585 14783 8619
rect 6653 8517 6687 8551
rect 6837 8517 6871 8551
rect 13461 8517 13495 8551
rect 1777 8449 1811 8483
rect 2421 8449 2455 8483
rect 3065 8449 3099 8483
rect 6009 8449 6043 8483
rect 7757 8449 7791 8483
rect 8953 8449 8987 8483
rect 9413 8449 9447 8483
rect 9689 8449 9723 8483
rect 12265 8449 12299 8483
rect 14657 8449 14691 8483
rect 15669 8449 15703 8483
rect 17049 8449 17083 8483
rect 7481 8381 7515 8415
rect 12357 8381 12391 8415
rect 12449 8381 12483 8415
rect 13553 8381 13587 8415
rect 13737 8381 13771 8415
rect 14933 8381 14967 8415
rect 1593 8313 1627 8347
rect 2237 8313 2271 8347
rect 2881 8313 2915 8347
rect 8769 8313 8803 8347
rect 14289 8313 14323 8347
rect 10885 8245 10919 8279
rect 1593 8041 1627 8075
rect 2881 8041 2915 8075
rect 9597 8041 9631 8075
rect 12081 8041 12115 8075
rect 12725 8041 12759 8075
rect 13369 8041 13403 8075
rect 23949 8041 23983 8075
rect 7941 7973 7975 8007
rect 8585 7973 8619 8007
rect 15209 7973 15243 8007
rect 10517 7905 10551 7939
rect 10977 7905 11011 7939
rect 14841 7905 14875 7939
rect 22201 7905 22235 7939
rect 1777 7837 1811 7871
rect 2421 7837 2455 7871
rect 3065 7837 3099 7871
rect 10241 7837 10275 7871
rect 10701 7837 10735 7871
rect 15025 7837 15059 7871
rect 22477 7769 22511 7803
rect 2237 7701 2271 7735
rect 9873 7701 9907 7735
rect 10333 7701 10367 7735
rect 2237 7497 2271 7531
rect 9597 7497 9631 7531
rect 9965 7497 9999 7531
rect 1777 7361 1811 7395
rect 2421 7361 2455 7395
rect 10057 7361 10091 7395
rect 10977 7361 11011 7395
rect 12081 7361 12115 7395
rect 13829 7361 13863 7395
rect 10149 7293 10183 7327
rect 1593 7225 1627 7259
rect 11897 7225 11931 7259
rect 13645 7157 13679 7191
rect 23305 6953 23339 6987
rect 1777 6749 1811 6783
rect 2421 6749 2455 6783
rect 3065 6749 3099 6783
rect 23029 6749 23063 6783
rect 1593 6613 1627 6647
rect 2237 6613 2271 6647
rect 2881 6613 2915 6647
rect 23489 6613 23523 6647
rect 22452 6273 22486 6307
rect 1593 6205 1627 6239
rect 1869 6205 1903 6239
rect 22523 6069 22557 6103
rect 18889 5865 18923 5899
rect 21005 5865 21039 5899
rect 15577 5729 15611 5763
rect 15761 5729 15795 5763
rect 17141 5729 17175 5763
rect 24777 5729 24811 5763
rect 26893 5729 26927 5763
rect 1593 5661 1627 5695
rect 1869 5661 1903 5695
rect 20913 5661 20947 5695
rect 24593 5661 24627 5695
rect 17417 5593 17451 5627
rect 26433 5593 26467 5627
rect 27077 5593 27111 5627
rect 28733 5593 28767 5627
rect 16221 5525 16255 5559
rect 21373 5525 21407 5559
rect 22891 5321 22925 5355
rect 1593 5185 1627 5219
rect 1869 5185 1903 5219
rect 15577 5185 15611 5219
rect 17509 5185 17543 5219
rect 22144 5185 22178 5219
rect 22788 5185 22822 5219
rect 15761 5117 15795 5151
rect 17693 5117 17727 5151
rect 28641 5117 28675 5151
rect 28825 5117 28859 5151
rect 30297 5117 30331 5151
rect 16221 4981 16255 5015
rect 18153 4981 18187 5015
rect 22247 4981 22281 5015
rect 19533 4777 19567 4811
rect 24731 4777 24765 4811
rect 1593 4641 1627 4675
rect 25789 4641 25823 4675
rect 1869 4573 1903 4607
rect 19441 4573 19475 4607
rect 24628 4573 24662 4607
rect 25973 4505 26007 4539
rect 27629 4505 27663 4539
rect 19901 4437 19935 4471
rect 3065 4097 3099 4131
rect 15209 4097 15243 4131
rect 1593 4029 1627 4063
rect 1869 4029 1903 4063
rect 2881 3961 2915 3995
rect 15025 3893 15059 3927
rect 2237 3689 2271 3723
rect 2881 3689 2915 3723
rect 1593 3621 1627 3655
rect 1777 3485 1811 3519
rect 2421 3485 2455 3519
rect 3065 3485 3099 3519
rect 11529 3485 11563 3519
rect 11621 3349 11655 3383
rect 2881 3145 2915 3179
rect 14013 3145 14047 3179
rect 12633 3077 12667 3111
rect 13921 3077 13955 3111
rect 15577 3077 15611 3111
rect 1869 3009 1903 3043
rect 3065 3009 3099 3043
rect 8861 3009 8895 3043
rect 17049 3009 17083 3043
rect 18337 3009 18371 3043
rect 20545 3009 20579 3043
rect 1593 2941 1627 2975
rect 9137 2941 9171 2975
rect 10609 2941 10643 2975
rect 15761 2873 15795 2907
rect 12725 2805 12759 2839
rect 16865 2805 16899 2839
rect 18153 2805 18187 2839
rect 20361 2805 20395 2839
rect 25513 2601 25547 2635
rect 28181 2601 28215 2635
rect 30849 2601 30883 2635
rect 33517 2601 33551 2635
rect 1869 2465 1903 2499
rect 4629 2465 4663 2499
rect 7297 2465 7331 2499
rect 9965 2465 9999 2499
rect 12633 2465 12667 2499
rect 15301 2465 15335 2499
rect 17969 2465 18003 2499
rect 20545 2465 20579 2499
rect 23121 2465 23155 2499
rect 36369 2465 36403 2499
rect 1593 2397 1627 2431
rect 3065 2397 3099 2431
rect 4353 2397 4387 2431
rect 7021 2397 7055 2431
rect 9597 2397 9631 2431
rect 12357 2397 12391 2431
rect 15025 2397 15059 2431
rect 17509 2397 17543 2431
rect 20085 2397 20119 2431
rect 22661 2397 22695 2431
rect 25697 2397 25731 2431
rect 28365 2397 28399 2431
rect 31033 2397 31067 2431
rect 33701 2397 33735 2431
rect 36093 2397 36127 2431
rect 2881 2261 2915 2295
<< metal1 >>
rect 20806 25508 20812 25560
rect 20864 25548 20870 25560
rect 24118 25548 24124 25560
rect 20864 25520 24124 25548
rect 20864 25508 20870 25520
rect 24118 25508 24124 25520
rect 24176 25508 24182 25560
rect 13446 25440 13452 25492
rect 13504 25480 13510 25492
rect 31754 25480 31760 25492
rect 13504 25452 31760 25480
rect 13504 25440 13510 25452
rect 31754 25440 31760 25452
rect 31812 25440 31818 25492
rect 10870 25372 10876 25424
rect 10928 25412 10934 25424
rect 34514 25412 34520 25424
rect 10928 25384 34520 25412
rect 10928 25372 10934 25384
rect 34514 25372 34520 25384
rect 34572 25372 34578 25424
rect 12250 25304 12256 25356
rect 12308 25344 12314 25356
rect 32122 25344 32128 25356
rect 12308 25316 32128 25344
rect 12308 25304 12314 25316
rect 32122 25304 32128 25316
rect 32180 25304 32186 25356
rect 11054 25236 11060 25288
rect 11112 25276 11118 25288
rect 33410 25276 33416 25288
rect 11112 25248 33416 25276
rect 11112 25236 11118 25248
rect 33410 25236 33416 25248
rect 33468 25236 33474 25288
rect 12158 25168 12164 25220
rect 12216 25208 12222 25220
rect 34146 25208 34152 25220
rect 12216 25180 34152 25208
rect 12216 25168 12222 25180
rect 34146 25168 34152 25180
rect 34204 25168 34210 25220
rect 9950 25100 9956 25152
rect 10008 25140 10014 25152
rect 32030 25140 32036 25152
rect 10008 25112 32036 25140
rect 10008 25100 10014 25112
rect 32030 25100 32036 25112
rect 32088 25100 32094 25152
rect 15838 25032 15844 25084
rect 15896 25072 15902 25084
rect 39298 25072 39304 25084
rect 15896 25044 39304 25072
rect 15896 25032 15902 25044
rect 39298 25032 39304 25044
rect 39356 25032 39362 25084
rect 11422 24964 11428 25016
rect 11480 25004 11486 25016
rect 35894 25004 35900 25016
rect 11480 24976 35900 25004
rect 11480 24964 11486 24976
rect 35894 24964 35900 24976
rect 35952 24964 35958 25016
rect 13906 24896 13912 24948
rect 13964 24936 13970 24948
rect 38654 24936 38660 24948
rect 13964 24908 38660 24936
rect 13964 24896 13970 24908
rect 38654 24896 38660 24908
rect 38712 24896 38718 24948
rect 3326 24828 3332 24880
rect 3384 24868 3390 24880
rect 8570 24868 8576 24880
rect 3384 24840 8576 24868
rect 3384 24828 3390 24840
rect 8570 24828 8576 24840
rect 8628 24828 8634 24880
rect 22554 24868 22560 24880
rect 22204 24840 22560 24868
rect 17218 24760 17224 24812
rect 17276 24800 17282 24812
rect 18598 24800 18604 24812
rect 17276 24772 18604 24800
rect 17276 24760 17282 24772
rect 18598 24760 18604 24772
rect 18656 24800 18662 24812
rect 22204 24800 22232 24840
rect 22554 24828 22560 24840
rect 22612 24828 22618 24880
rect 18656 24772 22232 24800
rect 18656 24760 18662 24772
rect 22278 24760 22284 24812
rect 22336 24800 22342 24812
rect 25958 24800 25964 24812
rect 22336 24772 25964 24800
rect 22336 24760 22342 24772
rect 25958 24760 25964 24772
rect 26016 24760 26022 24812
rect 26050 24760 26056 24812
rect 26108 24800 26114 24812
rect 28626 24800 28632 24812
rect 26108 24772 28632 24800
rect 26108 24760 26114 24772
rect 28626 24760 28632 24772
rect 28684 24760 28690 24812
rect 9582 24692 9588 24744
rect 9640 24732 9646 24744
rect 23474 24732 23480 24744
rect 9640 24704 23480 24732
rect 9640 24692 9646 24704
rect 23474 24692 23480 24704
rect 23532 24692 23538 24744
rect 25222 24692 25228 24744
rect 25280 24732 25286 24744
rect 29086 24732 29092 24744
rect 25280 24704 29092 24732
rect 25280 24692 25286 24704
rect 29086 24692 29092 24704
rect 29144 24692 29150 24744
rect 9122 24624 9128 24676
rect 9180 24664 9186 24676
rect 18782 24664 18788 24676
rect 9180 24636 18788 24664
rect 9180 24624 9186 24636
rect 18782 24624 18788 24636
rect 18840 24624 18846 24676
rect 19058 24624 19064 24676
rect 19116 24664 19122 24676
rect 25866 24664 25872 24676
rect 19116 24636 25872 24664
rect 19116 24624 19122 24636
rect 25866 24624 25872 24636
rect 25924 24624 25930 24676
rect 25958 24624 25964 24676
rect 26016 24664 26022 24676
rect 32306 24664 32312 24676
rect 26016 24636 32312 24664
rect 26016 24624 26022 24636
rect 32306 24624 32312 24636
rect 32364 24624 32370 24676
rect 12342 24556 12348 24608
rect 12400 24596 12406 24608
rect 25774 24596 25780 24608
rect 12400 24568 25780 24596
rect 12400 24556 12406 24568
rect 25774 24556 25780 24568
rect 25832 24556 25838 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 9122 24352 9128 24404
rect 9180 24352 9186 24404
rect 9232 24364 18736 24392
rect 7466 24284 7472 24336
rect 7524 24324 7530 24336
rect 9232 24324 9260 24364
rect 7524 24296 9260 24324
rect 7524 24284 7530 24296
rect 9306 24284 9312 24336
rect 9364 24284 9370 24336
rect 11701 24327 11759 24333
rect 11701 24293 11713 24327
rect 11747 24293 11759 24327
rect 11701 24287 11759 24293
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3510 24256 3516 24268
rect 3283 24228 3516 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 7374 24256 7380 24268
rect 5859 24228 7380 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 7374 24216 7380 24228
rect 7432 24216 7438 24268
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9324 24256 9352 24284
rect 8251 24228 9352 24256
rect 11716 24256 11744 24287
rect 11790 24284 11796 24336
rect 11848 24324 11854 24336
rect 13814 24324 13820 24336
rect 11848 24296 13820 24324
rect 11848 24284 11854 24296
rect 13814 24284 13820 24296
rect 13872 24284 13878 24336
rect 13541 24259 13599 24265
rect 11716 24228 13400 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2406 24188 2412 24200
rect 2271 24160 2412 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2406 24148 2412 24160
rect 2464 24148 2470 24200
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24157 4215 24191
rect 4157 24151 4215 24157
rect 4172 24120 4200 24151
rect 4798 24148 4804 24200
rect 4856 24148 4862 24200
rect 6638 24148 6644 24200
rect 6696 24188 6702 24200
rect 6733 24191 6791 24197
rect 6733 24188 6745 24191
rect 6696 24160 6745 24188
rect 6696 24148 6702 24160
rect 6733 24157 6745 24160
rect 6779 24157 6791 24191
rect 6733 24151 6791 24157
rect 6822 24148 6828 24200
rect 6880 24188 6886 24200
rect 7193 24191 7251 24197
rect 7193 24188 7205 24191
rect 6880 24160 7205 24188
rect 6880 24148 6886 24160
rect 7193 24157 7205 24160
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24188 9367 24191
rect 9582 24188 9588 24200
rect 9355 24160 9588 24188
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 9950 24148 9956 24200
rect 10008 24148 10014 24200
rect 10873 24191 10931 24197
rect 10873 24157 10885 24191
rect 10919 24188 10931 24191
rect 11790 24188 11796 24200
rect 10919 24160 11796 24188
rect 10919 24157 10931 24160
rect 10873 24151 10931 24157
rect 11790 24148 11796 24160
rect 11848 24148 11854 24200
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 11974 24188 11980 24200
rect 11931 24160 11980 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 11974 24148 11980 24160
rect 12032 24148 12038 24200
rect 12526 24148 12532 24200
rect 12584 24148 12590 24200
rect 13372 24188 13400 24228
rect 13541 24225 13553 24259
rect 13587 24256 13599 24259
rect 14274 24256 14280 24268
rect 13587 24228 14280 24256
rect 13587 24225 13599 24228
rect 13541 24219 13599 24225
rect 14274 24216 14280 24228
rect 14332 24216 14338 24268
rect 16853 24259 16911 24265
rect 14384 24228 14964 24256
rect 14384 24188 14412 24228
rect 13372 24160 14412 24188
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 14936 24197 14964 24228
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 17126 24256 17132 24268
rect 16899 24228 17132 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 17126 24216 17132 24228
rect 17184 24216 17190 24268
rect 14921 24191 14979 24197
rect 14921 24157 14933 24191
rect 14967 24157 14979 24191
rect 14921 24151 14979 24157
rect 10042 24120 10048 24132
rect 4172 24092 10048 24120
rect 10042 24080 10048 24092
rect 10100 24080 10106 24132
rect 16117 24123 16175 24129
rect 16117 24089 16129 24123
rect 16163 24120 16175 24123
rect 16206 24120 16212 24132
rect 16163 24092 16212 24120
rect 16163 24089 16175 24092
rect 16117 24083 16175 24089
rect 16206 24080 16212 24092
rect 16264 24080 16270 24132
rect 17129 24123 17187 24129
rect 17129 24089 17141 24123
rect 17175 24120 17187 24123
rect 17218 24120 17224 24132
rect 17175 24092 17224 24120
rect 17175 24089 17187 24092
rect 17129 24083 17187 24089
rect 17218 24080 17224 24092
rect 17276 24080 17282 24132
rect 18506 24120 18512 24132
rect 18354 24092 18512 24120
rect 18506 24080 18512 24092
rect 18564 24080 18570 24132
rect 4706 24012 4712 24064
rect 4764 24052 4770 24064
rect 6549 24055 6607 24061
rect 6549 24052 6561 24055
rect 4764 24024 6561 24052
rect 4764 24012 4770 24024
rect 6549 24021 6561 24024
rect 6595 24021 6607 24055
rect 6549 24015 6607 24021
rect 10134 24012 10140 24064
rect 10192 24052 10198 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 10192 24024 14289 24052
rect 10192 24012 10198 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 14277 24015 14335 24021
rect 17494 24012 17500 24064
rect 17552 24052 17558 24064
rect 18601 24055 18659 24061
rect 18601 24052 18613 24055
rect 17552 24024 18613 24052
rect 17552 24012 17558 24024
rect 18601 24021 18613 24024
rect 18647 24021 18659 24055
rect 18708 24052 18736 24364
rect 21542 24352 21548 24404
rect 21600 24392 21606 24404
rect 21600 24364 22508 24392
rect 21600 24352 21606 24364
rect 19429 24327 19487 24333
rect 19429 24293 19441 24327
rect 19475 24324 19487 24327
rect 19475 24296 22140 24324
rect 19475 24293 19487 24296
rect 19429 24287 19487 24293
rect 19306 24228 20852 24256
rect 18782 24148 18788 24200
rect 18840 24188 18846 24200
rect 19306 24188 19334 24228
rect 18840 24160 19334 24188
rect 19613 24191 19671 24197
rect 18840 24148 18846 24160
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 19628 24120 19656 24151
rect 19794 24148 19800 24200
rect 19852 24188 19858 24200
rect 20073 24191 20131 24197
rect 20073 24188 20085 24191
rect 19852 24160 20085 24188
rect 19852 24148 19858 24160
rect 20073 24157 20085 24160
rect 20119 24157 20131 24191
rect 20824 24188 20852 24228
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 21542 24188 21548 24200
rect 20824 24160 21548 24188
rect 20073 24151 20131 24157
rect 21542 24148 21548 24160
rect 21600 24148 21606 24200
rect 21910 24188 21916 24200
rect 21744 24160 21916 24188
rect 21744 24120 21772 24160
rect 21910 24148 21916 24160
rect 21968 24148 21974 24200
rect 22112 24197 22140 24296
rect 22480 24265 22508 24364
rect 22554 24352 22560 24404
rect 22612 24392 22618 24404
rect 22612 24364 25636 24392
rect 22612 24352 22618 24364
rect 22465 24259 22523 24265
rect 22465 24225 22477 24259
rect 22511 24225 22523 24259
rect 22465 24219 22523 24225
rect 25222 24216 25228 24268
rect 25280 24216 25286 24268
rect 25608 24256 25636 24364
rect 25774 24352 25780 24404
rect 25832 24352 25838 24404
rect 25866 24352 25872 24404
rect 25924 24392 25930 24404
rect 25924 24364 27016 24392
rect 25924 24352 25930 24364
rect 26329 24259 26387 24265
rect 26329 24256 26341 24259
rect 25608 24228 26341 24256
rect 26329 24225 26341 24228
rect 26375 24225 26387 24259
rect 26988 24256 27016 24364
rect 27246 24352 27252 24404
rect 27304 24392 27310 24404
rect 30374 24392 30380 24404
rect 27304 24364 30380 24392
rect 27304 24352 27310 24364
rect 30374 24352 30380 24364
rect 30432 24352 30438 24404
rect 32306 24352 32312 24404
rect 32364 24352 32370 24404
rect 33410 24352 33416 24404
rect 33468 24352 33474 24404
rect 34146 24352 34152 24404
rect 34204 24352 34210 24404
rect 34514 24352 34520 24404
rect 34572 24392 34578 24404
rect 35069 24395 35127 24401
rect 35069 24392 35081 24395
rect 34572 24364 35081 24392
rect 34572 24352 34578 24364
rect 35069 24361 35081 24364
rect 35115 24361 35127 24395
rect 35069 24355 35127 24361
rect 35805 24395 35863 24401
rect 35805 24361 35817 24395
rect 35851 24392 35863 24395
rect 35894 24392 35900 24404
rect 35851 24364 35900 24392
rect 35851 24361 35863 24364
rect 35805 24355 35863 24361
rect 35894 24352 35900 24364
rect 35952 24352 35958 24404
rect 39298 24352 39304 24404
rect 39356 24352 39362 24404
rect 28074 24284 28080 24336
rect 28132 24324 28138 24336
rect 46845 24327 46903 24333
rect 46845 24324 46857 24327
rect 28132 24296 30052 24324
rect 28132 24284 28138 24296
rect 27709 24259 27767 24265
rect 27709 24256 27721 24259
rect 26988 24228 27721 24256
rect 26329 24219 26387 24225
rect 27709 24225 27721 24228
rect 27755 24225 27767 24259
rect 27709 24219 27767 24225
rect 28350 24216 28356 24268
rect 28408 24256 28414 24268
rect 28408 24228 29316 24256
rect 28408 24216 28414 24228
rect 22097 24191 22155 24197
rect 22097 24157 22109 24191
rect 22143 24157 22155 24191
rect 22097 24151 22155 24157
rect 24029 24191 24087 24197
rect 24029 24157 24041 24191
rect 24075 24188 24087 24191
rect 25406 24188 25412 24200
rect 24075 24160 25412 24188
rect 24075 24157 24087 24160
rect 24029 24151 24087 24157
rect 25406 24148 25412 24160
rect 25464 24148 25470 24200
rect 26694 24148 26700 24200
rect 26752 24188 26758 24200
rect 28537 24191 28595 24197
rect 28537 24188 28549 24191
rect 26752 24160 28549 24188
rect 26752 24148 26758 24160
rect 28537 24157 28549 24160
rect 28583 24157 28595 24191
rect 28537 24151 28595 24157
rect 28626 24148 28632 24200
rect 28684 24188 28690 24200
rect 29181 24191 29239 24197
rect 29181 24188 29193 24191
rect 28684 24160 29193 24188
rect 28684 24148 28690 24160
rect 29181 24157 29193 24160
rect 29227 24157 29239 24191
rect 29288 24188 29316 24228
rect 29546 24216 29552 24268
rect 29604 24256 29610 24268
rect 30024 24265 30052 24296
rect 30208 24296 46857 24324
rect 29733 24259 29791 24265
rect 29733 24256 29745 24259
rect 29604 24228 29745 24256
rect 29604 24216 29610 24228
rect 29733 24225 29745 24228
rect 29779 24225 29791 24259
rect 29733 24219 29791 24225
rect 30009 24259 30067 24265
rect 30009 24225 30021 24259
rect 30055 24225 30067 24259
rect 30009 24219 30067 24225
rect 30208 24188 30236 24296
rect 46845 24293 46857 24296
rect 46891 24293 46903 24327
rect 46845 24287 46903 24293
rect 31938 24216 31944 24268
rect 31996 24256 32002 24268
rect 31996 24228 39344 24256
rect 31996 24216 32002 24228
rect 29288 24160 30236 24188
rect 29181 24151 29239 24157
rect 30558 24148 30564 24200
rect 30616 24188 30622 24200
rect 31481 24191 31539 24197
rect 31481 24188 31493 24191
rect 30616 24160 31493 24188
rect 30616 24148 30622 24160
rect 31481 24157 31493 24160
rect 31527 24157 31539 24191
rect 31481 24151 31539 24157
rect 32493 24191 32551 24197
rect 32493 24157 32505 24191
rect 32539 24157 32551 24191
rect 32493 24151 32551 24157
rect 27617 24123 27675 24129
rect 27617 24120 27629 24123
rect 19628 24092 21772 24120
rect 23860 24092 27629 24120
rect 20806 24052 20812 24064
rect 18708 24024 20812 24052
rect 18601 24015 18659 24021
rect 20806 24012 20812 24024
rect 20864 24012 20870 24064
rect 23860 24061 23888 24092
rect 27617 24089 27629 24092
rect 27663 24089 27675 24123
rect 27617 24083 27675 24089
rect 28718 24080 28724 24132
rect 28776 24120 28782 24132
rect 32508 24120 32536 24151
rect 33318 24148 33324 24200
rect 33376 24148 33382 24200
rect 33778 24148 33784 24200
rect 33836 24188 33842 24200
rect 34057 24191 34115 24197
rect 34057 24188 34069 24191
rect 33836 24160 34069 24188
rect 33836 24148 33842 24160
rect 34057 24157 34069 24160
rect 34103 24157 34115 24191
rect 34057 24151 34115 24157
rect 34514 24148 34520 24200
rect 34572 24188 34578 24200
rect 34977 24191 35035 24197
rect 34977 24188 34989 24191
rect 34572 24160 34989 24188
rect 34572 24148 34578 24160
rect 34977 24157 34989 24160
rect 35023 24157 35035 24191
rect 34977 24151 35035 24157
rect 35066 24148 35072 24200
rect 35124 24188 35130 24200
rect 35713 24191 35771 24197
rect 35713 24188 35725 24191
rect 35124 24160 35725 24188
rect 35124 24148 35130 24160
rect 35713 24157 35725 24160
rect 35759 24157 35771 24191
rect 35713 24151 35771 24157
rect 35894 24148 35900 24200
rect 35952 24188 35958 24200
rect 36541 24191 36599 24197
rect 36541 24188 36553 24191
rect 35952 24160 36553 24188
rect 35952 24148 35958 24160
rect 36541 24157 36553 24160
rect 36587 24157 36599 24191
rect 36541 24151 36599 24157
rect 37274 24148 37280 24200
rect 37332 24188 37338 24200
rect 37645 24191 37703 24197
rect 37645 24188 37657 24191
rect 37332 24160 37657 24188
rect 37332 24148 37338 24160
rect 37645 24157 37657 24160
rect 37691 24157 37703 24191
rect 37645 24151 37703 24157
rect 38470 24148 38476 24200
rect 38528 24148 38534 24200
rect 38654 24148 38660 24200
rect 38712 24148 38718 24200
rect 39206 24148 39212 24200
rect 39264 24148 39270 24200
rect 39316 24188 39344 24228
rect 40034 24216 40040 24268
rect 40092 24216 40098 24268
rect 40313 24191 40371 24197
rect 40313 24188 40325 24191
rect 39316 24160 40325 24188
rect 40313 24157 40325 24160
rect 40359 24157 40371 24191
rect 40313 24151 40371 24157
rect 40586 24148 40592 24200
rect 40644 24188 40650 24200
rect 41509 24191 41567 24197
rect 41509 24188 41521 24191
rect 40644 24160 41521 24188
rect 40644 24148 40650 24160
rect 41509 24157 41521 24160
rect 41555 24157 41567 24191
rect 41509 24151 41567 24157
rect 41598 24148 41604 24200
rect 41656 24188 41662 24200
rect 42613 24191 42671 24197
rect 42613 24188 42625 24191
rect 41656 24160 42625 24188
rect 41656 24148 41662 24160
rect 42613 24157 42625 24160
rect 42659 24157 42671 24191
rect 42613 24151 42671 24157
rect 44726 24148 44732 24200
rect 44784 24188 44790 24200
rect 45189 24191 45247 24197
rect 45189 24188 45201 24191
rect 44784 24160 45201 24188
rect 44784 24148 44790 24160
rect 45189 24157 45201 24160
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 45554 24148 45560 24200
rect 45612 24188 45618 24200
rect 45925 24191 45983 24197
rect 45925 24188 45937 24191
rect 45612 24160 45937 24188
rect 45612 24148 45618 24160
rect 45925 24157 45937 24160
rect 45971 24157 45983 24191
rect 45925 24151 45983 24157
rect 46014 24148 46020 24200
rect 46072 24188 46078 24200
rect 46661 24191 46719 24197
rect 46661 24188 46673 24191
rect 46072 24160 46673 24188
rect 46072 24148 46078 24160
rect 46661 24157 46673 24160
rect 46707 24157 46719 24191
rect 46661 24151 46719 24157
rect 47302 24148 47308 24200
rect 47360 24188 47366 24200
rect 47765 24191 47823 24197
rect 47765 24188 47777 24191
rect 47360 24160 47777 24188
rect 47360 24148 47366 24160
rect 47765 24157 47777 24160
rect 47811 24157 47823 24191
rect 47765 24151 47823 24157
rect 47946 24148 47952 24200
rect 48004 24188 48010 24200
rect 48501 24191 48559 24197
rect 48501 24188 48513 24191
rect 48004 24160 48513 24188
rect 48004 24148 48010 24160
rect 48501 24157 48513 24160
rect 48547 24157 48559 24191
rect 48501 24151 48559 24157
rect 28776 24092 32536 24120
rect 28776 24080 28782 24092
rect 34698 24080 34704 24132
rect 34756 24120 34762 24132
rect 34756 24092 37504 24120
rect 34756 24080 34762 24092
rect 23845 24055 23903 24061
rect 23845 24021 23857 24055
rect 23891 24021 23903 24055
rect 23845 24015 23903 24021
rect 23934 24012 23940 24064
rect 23992 24052 23998 24064
rect 24581 24055 24639 24061
rect 24581 24052 24593 24055
rect 23992 24024 24593 24052
rect 23992 24012 23998 24024
rect 24581 24021 24593 24024
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 24670 24012 24676 24064
rect 24728 24052 24734 24064
rect 24949 24055 25007 24061
rect 24949 24052 24961 24055
rect 24728 24024 24961 24052
rect 24728 24012 24734 24024
rect 24949 24021 24961 24024
rect 24995 24021 25007 24055
rect 24949 24015 25007 24021
rect 25038 24012 25044 24064
rect 25096 24012 25102 24064
rect 25682 24012 25688 24064
rect 25740 24052 25746 24064
rect 26145 24055 26203 24061
rect 26145 24052 26157 24055
rect 25740 24024 26157 24052
rect 25740 24012 25746 24024
rect 26145 24021 26157 24024
rect 26191 24021 26203 24055
rect 26145 24015 26203 24021
rect 26234 24012 26240 24064
rect 26292 24012 26298 24064
rect 27154 24012 27160 24064
rect 27212 24012 27218 24064
rect 27430 24012 27436 24064
rect 27488 24052 27494 24064
rect 27525 24055 27583 24061
rect 27525 24052 27537 24055
rect 27488 24024 27537 24052
rect 27488 24012 27494 24024
rect 27525 24021 27537 24024
rect 27571 24021 27583 24055
rect 27525 24015 27583 24021
rect 27706 24012 27712 24064
rect 27764 24052 27770 24064
rect 28353 24055 28411 24061
rect 28353 24052 28365 24055
rect 27764 24024 28365 24052
rect 27764 24012 27770 24024
rect 28353 24021 28365 24024
rect 28399 24021 28411 24055
rect 28353 24015 28411 24021
rect 28994 24012 29000 24064
rect 29052 24012 29058 24064
rect 29178 24012 29184 24064
rect 29236 24052 29242 24064
rect 31297 24055 31355 24061
rect 31297 24052 31309 24055
rect 29236 24024 31309 24052
rect 29236 24012 29242 24024
rect 31297 24021 31309 24024
rect 31343 24021 31355 24055
rect 31297 24015 31355 24021
rect 34514 24012 34520 24064
rect 34572 24052 34578 24064
rect 37476 24061 37504 24092
rect 40034 24080 40040 24132
rect 40092 24120 40098 24132
rect 40092 24092 43944 24120
rect 40092 24080 40098 24092
rect 36357 24055 36415 24061
rect 36357 24052 36369 24055
rect 34572 24024 36369 24052
rect 34572 24012 34578 24024
rect 36357 24021 36369 24024
rect 36403 24021 36415 24055
rect 36357 24015 36415 24021
rect 37461 24055 37519 24061
rect 37461 24021 37473 24055
rect 37507 24021 37519 24055
rect 37461 24015 37519 24021
rect 38654 24012 38660 24064
rect 38712 24052 38718 24064
rect 43916 24061 43944 24092
rect 41325 24055 41383 24061
rect 41325 24052 41337 24055
rect 38712 24024 41337 24052
rect 38712 24012 38718 24024
rect 41325 24021 41337 24024
rect 41371 24021 41383 24055
rect 41325 24015 41383 24021
rect 43901 24055 43959 24061
rect 43901 24021 43913 24055
rect 43947 24021 43959 24055
rect 43901 24015 43959 24021
rect 45370 24012 45376 24064
rect 45428 24012 45434 24064
rect 46106 24012 46112 24064
rect 46164 24012 46170 24064
rect 46382 24012 46388 24064
rect 46440 24052 46446 24064
rect 47949 24055 48007 24061
rect 47949 24052 47961 24055
rect 46440 24024 47961 24052
rect 46440 24012 46446 24024
rect 47949 24021 47961 24024
rect 47995 24021 48007 24055
rect 47949 24015 48007 24021
rect 48685 24055 48743 24061
rect 48685 24021 48697 24055
rect 48731 24052 48743 24055
rect 48774 24052 48780 24064
rect 48731 24024 48780 24052
rect 48731 24021 48743 24024
rect 48685 24015 48743 24021
rect 48774 24012 48780 24024
rect 48832 24012 48838 24064
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 1578 23808 1584 23860
rect 1636 23848 1642 23860
rect 11885 23851 11943 23857
rect 11885 23848 11897 23851
rect 1636 23820 11897 23848
rect 1636 23808 1642 23820
rect 11885 23817 11897 23820
rect 11931 23817 11943 23851
rect 11885 23811 11943 23817
rect 12250 23808 12256 23860
rect 12308 23808 12314 23860
rect 12342 23808 12348 23860
rect 12400 23808 12406 23860
rect 14458 23808 14464 23860
rect 14516 23848 14522 23860
rect 21910 23848 21916 23860
rect 14516 23820 21916 23848
rect 14516 23808 14522 23820
rect 21910 23808 21916 23820
rect 21968 23808 21974 23860
rect 22020 23820 23612 23848
rect 2133 23783 2191 23789
rect 2133 23749 2145 23783
rect 2179 23780 2191 23783
rect 3786 23780 3792 23792
rect 2179 23752 3792 23780
rect 2179 23749 2191 23752
rect 2133 23743 2191 23749
rect 3786 23740 3792 23752
rect 3844 23740 3850 23792
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 4062 23780 4068 23792
rect 4019 23752 4068 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 4062 23740 4068 23752
rect 4120 23740 4126 23792
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9674 23780 9680 23792
rect 9171 23752 9680 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 9674 23740 9680 23752
rect 9732 23740 9738 23792
rect 10965 23783 11023 23789
rect 10965 23749 10977 23783
rect 11011 23780 11023 23783
rect 12434 23780 12440 23792
rect 11011 23752 12440 23780
rect 11011 23749 11023 23752
rect 10965 23743 11023 23749
rect 12434 23740 12440 23752
rect 12492 23740 12498 23792
rect 14277 23783 14335 23789
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 15746 23780 15752 23792
rect 14323 23752 15752 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 15746 23740 15752 23752
rect 15804 23740 15810 23792
rect 18141 23783 18199 23789
rect 18141 23749 18153 23783
rect 18187 23780 18199 23783
rect 19334 23780 19340 23792
rect 18187 23752 19340 23780
rect 18187 23749 18199 23752
rect 18141 23743 18199 23749
rect 19334 23740 19340 23752
rect 19392 23740 19398 23792
rect 21450 23780 21456 23792
rect 20286 23752 21456 23780
rect 21450 23740 21456 23752
rect 21508 23780 21514 23792
rect 22020 23780 22048 23820
rect 23584 23780 23612 23820
rect 25038 23808 25044 23860
rect 25096 23848 25102 23860
rect 27246 23848 27252 23860
rect 25096 23820 27252 23848
rect 25096 23808 25102 23820
rect 27246 23808 27252 23820
rect 27304 23808 27310 23860
rect 27338 23808 27344 23860
rect 27396 23848 27402 23860
rect 27396 23820 29592 23848
rect 27396 23808 27402 23820
rect 24486 23780 24492 23792
rect 21508 23752 22048 23780
rect 23506 23752 24492 23780
rect 21508 23740 21514 23752
rect 24486 23740 24492 23752
rect 24544 23740 24550 23792
rect 26602 23740 26608 23792
rect 26660 23780 26666 23792
rect 27433 23783 27491 23789
rect 27433 23780 27445 23783
rect 26660 23752 27445 23780
rect 26660 23740 26666 23752
rect 27433 23749 27445 23752
rect 27479 23749 27491 23783
rect 27433 23743 27491 23749
rect 28902 23740 28908 23792
rect 28960 23780 28966 23792
rect 29178 23780 29184 23792
rect 28960 23752 29184 23780
rect 28960 23740 28966 23752
rect 29178 23740 29184 23752
rect 29236 23740 29242 23792
rect 2777 23715 2835 23721
rect 2777 23681 2789 23715
rect 2823 23681 2835 23715
rect 2777 23675 2835 23681
rect 1118 23604 1124 23656
rect 1176 23644 1182 23656
rect 2792 23644 2820 23675
rect 4614 23672 4620 23724
rect 4672 23672 4678 23724
rect 4890 23672 4896 23724
rect 4948 23712 4954 23724
rect 6641 23715 6699 23721
rect 6641 23712 6653 23715
rect 4948 23684 6653 23712
rect 4948 23672 4954 23684
rect 6641 23681 6653 23684
rect 6687 23681 6699 23715
rect 6641 23675 6699 23681
rect 7466 23672 7472 23724
rect 7524 23672 7530 23724
rect 8110 23672 8116 23724
rect 8168 23672 8174 23724
rect 9950 23672 9956 23724
rect 10008 23672 10014 23724
rect 10042 23672 10048 23724
rect 10100 23712 10106 23724
rect 13265 23715 13323 23721
rect 10100 23684 13032 23712
rect 10100 23672 10106 23684
rect 1176 23616 2820 23644
rect 1176 23604 1182 23616
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 12529 23647 12587 23653
rect 12529 23613 12541 23647
rect 12575 23613 12587 23647
rect 13004 23644 13032 23684
rect 13265 23681 13277 23715
rect 13311 23712 13323 23715
rect 13446 23712 13452 23724
rect 13311 23684 13452 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 13446 23672 13452 23684
rect 13504 23672 13510 23724
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23681 15163 23715
rect 15105 23675 15163 23681
rect 13538 23644 13544 23656
rect 13004 23616 13544 23644
rect 12529 23607 12587 23613
rect 2314 23536 2320 23588
rect 2372 23536 2378 23588
rect 12544 23576 12572 23607
rect 13538 23604 13544 23616
rect 13596 23604 13602 23656
rect 15120 23644 15148 23675
rect 15194 23672 15200 23724
rect 15252 23712 15258 23724
rect 16945 23715 17003 23721
rect 16945 23712 16957 23715
rect 15252 23684 16957 23712
rect 15252 23672 15258 23684
rect 16945 23681 16957 23684
rect 16991 23681 17003 23715
rect 16945 23675 17003 23681
rect 21085 23715 21143 23721
rect 21085 23681 21097 23715
rect 21131 23712 21143 23715
rect 21726 23712 21732 23724
rect 21131 23684 21732 23712
rect 21131 23681 21143 23684
rect 21085 23675 21143 23681
rect 21726 23672 21732 23684
rect 21784 23672 21790 23724
rect 24397 23715 24455 23721
rect 24397 23681 24409 23715
rect 24443 23712 24455 23715
rect 24670 23712 24676 23724
rect 24443 23684 24676 23712
rect 24443 23681 24455 23684
rect 24397 23675 24455 23681
rect 24670 23672 24676 23684
rect 24728 23672 24734 23724
rect 26266 23684 27003 23712
rect 16117 23647 16175 23653
rect 15120 23616 15516 23644
rect 15286 23576 15292 23588
rect 12544 23548 15292 23576
rect 15286 23536 15292 23548
rect 15344 23536 15350 23588
rect 15488 23576 15516 23616
rect 16117 23613 16129 23647
rect 16163 23644 16175 23647
rect 18322 23644 18328 23656
rect 16163 23616 18328 23644
rect 16163 23613 16175 23616
rect 16117 23607 16175 23613
rect 18322 23604 18328 23616
rect 18380 23604 18386 23656
rect 18785 23647 18843 23653
rect 18785 23613 18797 23647
rect 18831 23644 18843 23647
rect 18831 23616 18920 23644
rect 18831 23613 18843 23616
rect 18785 23607 18843 23613
rect 17770 23576 17776 23588
rect 15488 23548 17776 23576
rect 17770 23536 17776 23548
rect 17828 23536 17834 23588
rect 1854 23468 1860 23520
rect 1912 23508 1918 23520
rect 6733 23511 6791 23517
rect 6733 23508 6745 23511
rect 1912 23480 6745 23508
rect 1912 23468 1918 23480
rect 6733 23477 6745 23480
rect 6779 23477 6791 23511
rect 6733 23471 6791 23477
rect 7285 23511 7343 23517
rect 7285 23477 7297 23511
rect 7331 23508 7343 23511
rect 12342 23508 12348 23520
rect 7331 23480 12348 23508
rect 7331 23477 7343 23480
rect 7285 23471 7343 23477
rect 12342 23468 12348 23480
rect 12400 23468 12406 23520
rect 18892 23508 18920 23616
rect 19058 23604 19064 23656
rect 19116 23604 19122 23656
rect 19610 23604 19616 23656
rect 19668 23644 19674 23656
rect 19668 23616 20116 23644
rect 19668 23604 19674 23616
rect 20088 23576 20116 23616
rect 20346 23604 20352 23656
rect 20404 23644 20410 23656
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 20404 23616 22017 23644
rect 20404 23604 20410 23616
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22281 23647 22339 23653
rect 22281 23644 22293 23647
rect 22005 23607 22063 23613
rect 22112 23616 22293 23644
rect 21269 23579 21327 23585
rect 21269 23576 21281 23579
rect 20088 23548 21281 23576
rect 21269 23545 21281 23548
rect 21315 23545 21327 23579
rect 21269 23539 21327 23545
rect 21818 23536 21824 23588
rect 21876 23576 21882 23588
rect 22112 23576 22140 23616
rect 22281 23613 22293 23616
rect 22327 23613 22339 23647
rect 22281 23607 22339 23613
rect 24854 23604 24860 23656
rect 24912 23604 24918 23656
rect 25133 23647 25191 23653
rect 25133 23613 25145 23647
rect 25179 23644 25191 23647
rect 25866 23644 25872 23656
rect 25179 23616 25872 23644
rect 25179 23613 25191 23616
rect 25133 23607 25191 23613
rect 25866 23604 25872 23616
rect 25924 23604 25930 23656
rect 26878 23644 26884 23656
rect 26160 23616 26884 23644
rect 21876 23548 22140 23576
rect 21876 23536 21882 23548
rect 19702 23508 19708 23520
rect 18892 23480 19708 23508
rect 19702 23468 19708 23480
rect 19760 23468 19766 23520
rect 20070 23468 20076 23520
rect 20128 23508 20134 23520
rect 20533 23511 20591 23517
rect 20533 23508 20545 23511
rect 20128 23480 20545 23508
rect 20128 23468 20134 23480
rect 20533 23477 20545 23480
rect 20579 23477 20591 23511
rect 20533 23471 20591 23477
rect 23750 23468 23756 23520
rect 23808 23468 23814 23520
rect 24854 23468 24860 23520
rect 24912 23508 24918 23520
rect 26160 23508 26188 23616
rect 26878 23604 26884 23616
rect 26936 23604 26942 23656
rect 26975 23644 27003 23684
rect 27062 23672 27068 23724
rect 27120 23712 27126 23724
rect 27157 23715 27215 23721
rect 27157 23712 27169 23715
rect 27120 23684 27169 23712
rect 27120 23672 27126 23684
rect 27157 23681 27169 23684
rect 27203 23681 27215 23715
rect 28994 23712 29000 23724
rect 28566 23698 29000 23712
rect 27157 23675 27215 23681
rect 28552 23684 29000 23698
rect 28552 23644 28580 23684
rect 28994 23672 29000 23684
rect 29052 23672 29058 23724
rect 29564 23721 29592 23820
rect 29730 23808 29736 23860
rect 29788 23848 29794 23860
rect 32309 23851 32367 23857
rect 32309 23848 32321 23851
rect 29788 23820 32321 23848
rect 29788 23808 29794 23820
rect 32309 23817 32321 23820
rect 32355 23817 32367 23851
rect 32309 23811 32367 23817
rect 32416 23820 33916 23848
rect 29638 23740 29644 23792
rect 29696 23780 29702 23792
rect 32416 23780 32444 23820
rect 29696 23752 32444 23780
rect 29696 23740 29702 23752
rect 32582 23740 32588 23792
rect 32640 23780 32646 23792
rect 32640 23752 33824 23780
rect 32640 23740 32646 23752
rect 29549 23715 29607 23721
rect 29549 23681 29561 23715
rect 29595 23681 29607 23715
rect 29549 23675 29607 23681
rect 30006 23672 30012 23724
rect 30064 23672 30070 23724
rect 31481 23715 31539 23721
rect 31481 23712 31493 23715
rect 30116 23684 31493 23712
rect 26975 23616 28580 23644
rect 28626 23604 28632 23656
rect 28684 23644 28690 23656
rect 30116 23644 30144 23684
rect 31481 23681 31493 23684
rect 31527 23681 31539 23715
rect 31481 23675 31539 23681
rect 31846 23672 31852 23724
rect 31904 23712 31910 23724
rect 33796 23721 33824 23752
rect 32493 23715 32551 23721
rect 32493 23712 32505 23715
rect 31904 23684 32505 23712
rect 31904 23672 31910 23684
rect 32493 23681 32505 23684
rect 32539 23681 32551 23715
rect 32493 23675 32551 23681
rect 33137 23715 33195 23721
rect 33137 23681 33149 23715
rect 33183 23681 33195 23715
rect 33137 23675 33195 23681
rect 33781 23715 33839 23721
rect 33781 23681 33793 23715
rect 33827 23681 33839 23715
rect 33781 23675 33839 23681
rect 28684 23616 30144 23644
rect 28684 23604 28690 23616
rect 30282 23604 30288 23656
rect 30340 23604 30346 23656
rect 31202 23604 31208 23656
rect 31260 23644 31266 23656
rect 33152 23644 33180 23675
rect 31260 23616 33180 23644
rect 33888 23644 33916 23820
rect 35158 23808 35164 23860
rect 35216 23808 35222 23860
rect 46106 23848 46112 23860
rect 35866 23820 46112 23848
rect 34517 23783 34575 23789
rect 34517 23749 34529 23783
rect 34563 23780 34575 23783
rect 34606 23780 34612 23792
rect 34563 23752 34612 23780
rect 34563 23749 34575 23752
rect 34517 23743 34575 23749
rect 34606 23740 34612 23752
rect 34664 23740 34670 23792
rect 35866 23780 35894 23820
rect 46106 23808 46112 23820
rect 46164 23808 46170 23860
rect 34716 23752 35894 23780
rect 34054 23672 34060 23724
rect 34112 23712 34118 23724
rect 34333 23715 34391 23721
rect 34333 23712 34345 23715
rect 34112 23684 34345 23712
rect 34112 23672 34118 23684
rect 34333 23681 34345 23684
rect 34379 23681 34391 23715
rect 34333 23675 34391 23681
rect 34422 23672 34428 23724
rect 34480 23712 34486 23724
rect 34716 23712 34744 23752
rect 35986 23740 35992 23792
rect 36044 23740 36050 23792
rect 43622 23740 43628 23792
rect 43680 23740 43686 23792
rect 34480 23684 34744 23712
rect 34480 23672 34486 23684
rect 35066 23672 35072 23724
rect 35124 23672 35130 23724
rect 35802 23672 35808 23724
rect 35860 23672 35866 23724
rect 36630 23672 36636 23724
rect 36688 23672 36694 23724
rect 37642 23672 37648 23724
rect 37700 23712 37706 23724
rect 37921 23715 37979 23721
rect 37921 23712 37933 23715
rect 37700 23684 37933 23712
rect 37700 23672 37706 23684
rect 37921 23681 37933 23684
rect 37967 23681 37979 23715
rect 37921 23675 37979 23681
rect 41138 23672 41144 23724
rect 41196 23712 41202 23724
rect 41509 23715 41567 23721
rect 41509 23712 41521 23715
rect 41196 23684 41521 23712
rect 41196 23672 41202 23684
rect 41509 23681 41521 23684
rect 41555 23681 41567 23715
rect 41509 23675 41567 23681
rect 44174 23672 44180 23724
rect 44232 23712 44238 23724
rect 44269 23715 44327 23721
rect 44269 23712 44281 23715
rect 44232 23684 44281 23712
rect 44232 23672 44238 23684
rect 44269 23681 44281 23684
rect 44315 23681 44327 23715
rect 44269 23675 44327 23681
rect 46658 23672 46664 23724
rect 46716 23712 46722 23724
rect 46753 23715 46811 23721
rect 46753 23712 46765 23715
rect 46716 23684 46765 23712
rect 46716 23672 46722 23684
rect 46753 23681 46765 23684
rect 46799 23681 46811 23715
rect 46753 23675 46811 23681
rect 48314 23672 48320 23724
rect 48372 23672 48378 23724
rect 49050 23672 49056 23724
rect 49108 23672 49114 23724
rect 33888 23616 35894 23644
rect 31260 23604 31266 23616
rect 26234 23536 26240 23588
rect 26292 23576 26298 23588
rect 29365 23579 29423 23585
rect 29365 23576 29377 23579
rect 26292 23548 26740 23576
rect 26292 23536 26298 23548
rect 24912 23480 26188 23508
rect 24912 23468 24918 23480
rect 26602 23468 26608 23520
rect 26660 23468 26666 23520
rect 26712 23508 26740 23548
rect 28460 23548 29377 23576
rect 28460 23508 28488 23548
rect 29365 23545 29377 23548
rect 29411 23545 29423 23579
rect 29365 23539 29423 23545
rect 31018 23536 31024 23588
rect 31076 23576 31082 23588
rect 33597 23579 33655 23585
rect 33597 23576 33609 23579
rect 31076 23548 33609 23576
rect 31076 23536 31082 23548
rect 33597 23545 33609 23548
rect 33643 23545 33655 23579
rect 35866 23576 35894 23616
rect 37182 23604 37188 23656
rect 37240 23644 37246 23656
rect 37240 23616 44496 23644
rect 37240 23604 37246 23616
rect 44468 23585 44496 23616
rect 43809 23579 43867 23585
rect 43809 23576 43821 23579
rect 35866 23548 43821 23576
rect 33597 23539 33655 23545
rect 43809 23545 43821 23548
rect 43855 23545 43867 23579
rect 43809 23539 43867 23545
rect 44453 23579 44511 23585
rect 44453 23545 44465 23579
rect 44499 23545 44511 23579
rect 44453 23539 44511 23545
rect 26712 23480 28488 23508
rect 28718 23468 28724 23520
rect 28776 23508 28782 23520
rect 28905 23511 28963 23517
rect 28905 23508 28917 23511
rect 28776 23480 28917 23508
rect 28776 23468 28782 23480
rect 28905 23477 28917 23480
rect 28951 23477 28963 23511
rect 28905 23471 28963 23477
rect 30558 23468 30564 23520
rect 30616 23508 30622 23520
rect 31297 23511 31355 23517
rect 31297 23508 31309 23511
rect 30616 23480 31309 23508
rect 30616 23468 30622 23480
rect 31297 23477 31309 23480
rect 31343 23477 31355 23511
rect 31297 23471 31355 23477
rect 31754 23468 31760 23520
rect 31812 23508 31818 23520
rect 32953 23511 33011 23517
rect 32953 23508 32965 23511
rect 31812 23480 32965 23508
rect 31812 23468 31818 23480
rect 32953 23477 32965 23480
rect 32999 23477 33011 23511
rect 32953 23471 33011 23477
rect 35250 23468 35256 23520
rect 35308 23508 35314 23520
rect 36449 23511 36507 23517
rect 36449 23508 36461 23511
rect 35308 23480 36461 23508
rect 35308 23468 35314 23480
rect 36449 23477 36461 23480
rect 36495 23477 36507 23511
rect 36449 23471 36507 23477
rect 37734 23468 37740 23520
rect 37792 23468 37798 23520
rect 41322 23468 41328 23520
rect 41380 23468 41386 23520
rect 46934 23468 46940 23520
rect 46992 23468 46998 23520
rect 48498 23468 48504 23520
rect 48556 23468 48562 23520
rect 48682 23468 48688 23520
rect 48740 23508 48746 23520
rect 49237 23511 49295 23517
rect 49237 23508 49249 23511
rect 48740 23480 49249 23508
rect 48740 23468 48746 23480
rect 49237 23477 49249 23480
rect 49283 23477 49295 23511
rect 49237 23471 49295 23477
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 1670 23264 1676 23316
rect 1728 23304 1734 23316
rect 14461 23307 14519 23313
rect 14461 23304 14473 23307
rect 1728 23276 14473 23304
rect 1728 23264 1734 23276
rect 14461 23273 14473 23276
rect 14507 23273 14519 23307
rect 14461 23267 14519 23273
rect 16206 23264 16212 23316
rect 16264 23304 16270 23316
rect 18966 23304 18972 23316
rect 16264 23276 18972 23304
rect 16264 23264 16270 23276
rect 18966 23264 18972 23276
rect 19024 23264 19030 23316
rect 19429 23307 19487 23313
rect 19429 23273 19441 23307
rect 19475 23304 19487 23307
rect 19518 23304 19524 23316
rect 19475 23276 19524 23304
rect 19475 23273 19487 23276
rect 19429 23267 19487 23273
rect 19518 23264 19524 23276
rect 19576 23264 19582 23316
rect 24762 23304 24768 23316
rect 19628 23276 24768 23304
rect 2866 23196 2872 23248
rect 2924 23236 2930 23248
rect 4154 23236 4160 23248
rect 2924 23208 4160 23236
rect 2924 23196 2930 23208
rect 4154 23196 4160 23208
rect 4212 23196 4218 23248
rect 5353 23239 5411 23245
rect 5353 23205 5365 23239
rect 5399 23236 5411 23239
rect 9030 23236 9036 23248
rect 5399 23208 9036 23236
rect 5399 23205 5411 23208
rect 5353 23199 5411 23205
rect 3973 23171 4031 23177
rect 3973 23137 3985 23171
rect 4019 23168 4031 23171
rect 5368 23168 5396 23199
rect 9030 23196 9036 23208
rect 9088 23196 9094 23248
rect 18877 23239 18935 23245
rect 18877 23205 18889 23239
rect 18923 23236 18935 23239
rect 19058 23236 19064 23248
rect 18923 23208 19064 23236
rect 18923 23205 18935 23208
rect 18877 23199 18935 23205
rect 19058 23196 19064 23208
rect 19116 23196 19122 23248
rect 4019 23140 5396 23168
rect 4019 23137 4031 23140
rect 3973 23131 4031 23137
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 11425 23171 11483 23177
rect 11425 23137 11437 23171
rect 11471 23168 11483 23171
rect 12434 23168 12440 23180
rect 11471 23140 12440 23168
rect 11471 23137 11483 23140
rect 11425 23131 11483 23137
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 12710 23128 12716 23180
rect 12768 23168 12774 23180
rect 15194 23168 15200 23180
rect 12768 23140 15200 23168
rect 12768 23128 12774 23140
rect 15194 23128 15200 23140
rect 15252 23128 15258 23180
rect 16485 23171 16543 23177
rect 16485 23137 16497 23171
rect 16531 23168 16543 23171
rect 17402 23168 17408 23180
rect 16531 23140 17408 23168
rect 16531 23137 16543 23140
rect 16485 23131 16543 23137
rect 17402 23128 17408 23140
rect 17460 23128 17466 23180
rect 1762 23060 1768 23112
rect 1820 23060 1826 23112
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23069 4307 23103
rect 4249 23063 4307 23069
rect 2774 22992 2780 23044
rect 2832 22992 2838 23044
rect 4264 23032 4292 23063
rect 5442 23060 5448 23112
rect 5500 23060 5506 23112
rect 7282 23060 7288 23112
rect 7340 23060 7346 23112
rect 8478 23060 8484 23112
rect 8536 23100 8542 23112
rect 9217 23103 9275 23109
rect 9217 23100 9229 23103
rect 8536 23072 9229 23100
rect 8536 23060 8542 23072
rect 9217 23069 9229 23072
rect 9263 23069 9275 23103
rect 9217 23063 9275 23069
rect 10962 23060 10968 23112
rect 11020 23100 11026 23112
rect 15473 23103 15531 23109
rect 11020 23072 11192 23100
rect 11020 23060 11026 23072
rect 4264 23004 8340 23032
rect 3878 22924 3884 22976
rect 3936 22964 3942 22976
rect 4798 22964 4804 22976
rect 3936 22936 4804 22964
rect 3936 22924 3942 22936
rect 4798 22924 4804 22936
rect 4856 22924 4862 22976
rect 4982 22924 4988 22976
rect 5040 22964 5046 22976
rect 8202 22964 8208 22976
rect 5040 22936 8208 22964
rect 5040 22924 5046 22936
rect 8202 22924 8208 22936
rect 8260 22924 8266 22976
rect 8312 22964 8340 23004
rect 9490 22992 9496 23044
rect 9548 22992 9554 23044
rect 10778 23032 10784 23044
rect 10718 23004 10784 23032
rect 10778 22992 10784 23004
rect 10836 22992 10842 23044
rect 11164 23032 11192 23072
rect 15473 23069 15485 23103
rect 15519 23100 15531 23103
rect 16942 23100 16948 23112
rect 15519 23072 16948 23100
rect 15519 23069 15531 23072
rect 15473 23063 15531 23069
rect 16942 23060 16948 23072
rect 17000 23060 17006 23112
rect 17126 23060 17132 23112
rect 17184 23060 17190 23112
rect 18506 23060 18512 23112
rect 18564 23060 18570 23112
rect 19628 23109 19656 23276
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 25866 23264 25872 23316
rect 25924 23304 25930 23316
rect 27430 23304 27436 23316
rect 25924 23276 27436 23304
rect 25924 23264 25930 23276
rect 27430 23264 27436 23276
rect 27488 23264 27494 23316
rect 27614 23264 27620 23316
rect 27672 23304 27678 23316
rect 29730 23304 29736 23316
rect 27672 23276 29736 23304
rect 27672 23264 27678 23276
rect 29730 23264 29736 23276
rect 29788 23264 29794 23316
rect 30006 23304 30012 23316
rect 29840 23276 30012 23304
rect 22278 23196 22284 23248
rect 22336 23196 22342 23248
rect 23750 23196 23756 23248
rect 23808 23236 23814 23248
rect 23808 23208 26234 23236
rect 23808 23196 23814 23208
rect 19702 23128 19708 23180
rect 19760 23168 19766 23180
rect 20073 23171 20131 23177
rect 20073 23168 20085 23171
rect 19760 23140 20085 23168
rect 19760 23128 19766 23140
rect 20073 23137 20085 23140
rect 20119 23168 20131 23171
rect 20346 23168 20352 23180
rect 20119 23140 20352 23168
rect 20119 23137 20131 23140
rect 20073 23131 20131 23137
rect 20346 23128 20352 23140
rect 20404 23128 20410 23180
rect 22296 23168 22324 23196
rect 21652 23140 22324 23168
rect 22557 23171 22615 23177
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23069 19671 23103
rect 19613 23063 19671 23069
rect 21450 23060 21456 23112
rect 21508 23060 21514 23112
rect 11701 23035 11759 23041
rect 11701 23032 11713 23035
rect 10888 23004 11100 23032
rect 11164 23004 11713 23032
rect 10888 22964 10916 23004
rect 8312 22936 10916 22964
rect 10962 22924 10968 22976
rect 11020 22924 11026 22976
rect 11072 22964 11100 23004
rect 11701 23001 11713 23004
rect 11747 23001 11759 23035
rect 13814 23032 13820 23044
rect 12926 23004 13820 23032
rect 11701 22995 11759 23001
rect 13814 22992 13820 23004
rect 13872 22992 13878 23044
rect 14369 23035 14427 23041
rect 14369 23001 14381 23035
rect 14415 23001 14427 23035
rect 14369 22995 14427 23001
rect 12618 22964 12624 22976
rect 11072 22936 12624 22964
rect 12618 22924 12624 22936
rect 12676 22924 12682 22976
rect 13170 22924 13176 22976
rect 13228 22924 13234 22976
rect 14384 22964 14412 22995
rect 15286 22992 15292 23044
rect 15344 23032 15350 23044
rect 17405 23035 17463 23041
rect 17405 23032 17417 23035
rect 15344 23004 17417 23032
rect 15344 22992 15350 23004
rect 17405 23001 17417 23004
rect 17451 23032 17463 23035
rect 17494 23032 17500 23044
rect 17451 23004 17500 23032
rect 17451 23001 17463 23004
rect 17405 22995 17463 23001
rect 17494 22992 17500 23004
rect 17552 22992 17558 23044
rect 18800 23004 20300 23032
rect 18800 22964 18828 23004
rect 14384 22936 18828 22964
rect 20272 22964 20300 23004
rect 20346 22992 20352 23044
rect 20404 22992 20410 23044
rect 21652 22964 21680 23140
rect 22557 23137 22569 23171
rect 22603 23168 22615 23171
rect 23768 23168 23796 23196
rect 22603 23140 23796 23168
rect 22603 23137 22615 23140
rect 22557 23131 22615 23137
rect 25130 23128 25136 23180
rect 25188 23128 25194 23180
rect 25682 23128 25688 23180
rect 25740 23168 25746 23180
rect 25866 23168 25872 23180
rect 25740 23140 25872 23168
rect 25740 23128 25746 23140
rect 25866 23128 25872 23140
rect 25924 23168 25930 23180
rect 26206 23168 26234 23208
rect 26988 23208 27476 23236
rect 26329 23171 26387 23177
rect 26329 23168 26341 23171
rect 25924 23140 26096 23168
rect 26206 23140 26341 23168
rect 25924 23128 25930 23140
rect 22278 23060 22284 23112
rect 22336 23060 22342 23112
rect 23842 23060 23848 23112
rect 23900 23100 23906 23112
rect 25958 23100 25964 23112
rect 23900 23072 25964 23100
rect 23900 23060 23906 23072
rect 25958 23060 25964 23072
rect 26016 23060 26022 23112
rect 26068 23100 26096 23140
rect 26329 23137 26341 23140
rect 26375 23137 26387 23171
rect 26329 23131 26387 23137
rect 26145 23103 26203 23109
rect 26145 23100 26157 23103
rect 26068 23072 26157 23100
rect 26145 23069 26157 23072
rect 26191 23069 26203 23103
rect 26145 23063 26203 23069
rect 24486 23032 24492 23044
rect 23782 23004 24492 23032
rect 24486 22992 24492 23004
rect 24544 22992 24550 23044
rect 25041 23035 25099 23041
rect 25041 23001 25053 23035
rect 25087 23032 25099 23035
rect 26988 23032 27016 23208
rect 27062 23128 27068 23180
rect 27120 23168 27126 23180
rect 27341 23171 27399 23177
rect 27341 23168 27353 23171
rect 27120 23140 27353 23168
rect 27120 23128 27126 23140
rect 27341 23137 27353 23140
rect 27387 23137 27399 23171
rect 27448 23168 27476 23208
rect 29086 23196 29092 23248
rect 29144 23196 29150 23248
rect 29178 23196 29184 23248
rect 29236 23236 29242 23248
rect 29840 23236 29868 23276
rect 30006 23264 30012 23276
rect 30064 23304 30070 23316
rect 30064 23276 31248 23304
rect 30064 23264 30070 23276
rect 29236 23208 29868 23236
rect 29236 23196 29242 23208
rect 31110 23196 31116 23248
rect 31168 23196 31174 23248
rect 31220 23236 31248 23276
rect 32122 23264 32128 23316
rect 32180 23264 32186 23316
rect 40034 23236 40040 23248
rect 31220 23208 40040 23236
rect 28258 23168 28264 23180
rect 27448 23140 28264 23168
rect 27341 23131 27399 23137
rect 28258 23128 28264 23140
rect 28316 23128 28322 23180
rect 28350 23128 28356 23180
rect 28408 23168 28414 23180
rect 29733 23171 29791 23177
rect 29733 23168 29745 23171
rect 28408 23140 29745 23168
rect 28408 23128 28414 23140
rect 29733 23137 29745 23140
rect 29779 23168 29791 23171
rect 31128 23168 31156 23196
rect 29779 23140 31156 23168
rect 29779 23137 29791 23140
rect 29733 23131 29791 23137
rect 28994 23100 29000 23112
rect 28750 23072 29000 23100
rect 28994 23060 29000 23072
rect 29052 23100 29058 23112
rect 29178 23100 29184 23112
rect 29052 23072 29184 23100
rect 29052 23060 29058 23072
rect 29178 23060 29184 23072
rect 29236 23060 29242 23112
rect 31220 23100 31248 23208
rect 40034 23196 40040 23208
rect 40092 23196 40098 23248
rect 33413 23103 33471 23109
rect 33413 23100 33425 23103
rect 31142 23072 31248 23100
rect 31312 23072 33425 23100
rect 25087 23004 27016 23032
rect 27617 23035 27675 23041
rect 25087 23001 25099 23004
rect 25041 22995 25099 23001
rect 27617 23001 27629 23035
rect 27663 23032 27675 23035
rect 27663 23004 28028 23032
rect 27663 23001 27675 23004
rect 27617 22995 27675 23001
rect 20272 22936 21680 22964
rect 21818 22924 21824 22976
rect 21876 22924 21882 22976
rect 23382 22924 23388 22976
rect 23440 22964 23446 22976
rect 24029 22967 24087 22973
rect 24029 22964 24041 22967
rect 23440 22936 24041 22964
rect 23440 22924 23446 22936
rect 24029 22933 24041 22936
rect 24075 22933 24087 22967
rect 24029 22927 24087 22933
rect 24578 22924 24584 22976
rect 24636 22924 24642 22976
rect 24946 22924 24952 22976
rect 25004 22924 25010 22976
rect 25774 22924 25780 22976
rect 25832 22924 25838 22976
rect 26237 22967 26295 22973
rect 26237 22933 26249 22967
rect 26283 22964 26295 22967
rect 27706 22964 27712 22976
rect 26283 22936 27712 22964
rect 26283 22933 26295 22936
rect 26237 22927 26295 22933
rect 27706 22924 27712 22936
rect 27764 22924 27770 22976
rect 28000 22964 28028 23004
rect 29086 22992 29092 23044
rect 29144 23032 29150 23044
rect 30009 23035 30067 23041
rect 30009 23032 30021 23035
rect 29144 23004 30021 23032
rect 29144 22992 29150 23004
rect 30009 23001 30021 23004
rect 30055 23001 30067 23035
rect 30009 22995 30067 23001
rect 28626 22964 28632 22976
rect 28000 22936 28632 22964
rect 28626 22924 28632 22936
rect 28684 22924 28690 22976
rect 29546 22924 29552 22976
rect 29604 22964 29610 22976
rect 31312 22964 31340 23072
rect 33413 23069 33425 23072
rect 33459 23069 33471 23103
rect 33413 23063 33471 23069
rect 48590 23060 48596 23112
rect 48648 23060 48654 23112
rect 49050 23060 49056 23112
rect 49108 23060 49114 23112
rect 32674 22992 32680 23044
rect 32732 22992 32738 23044
rect 34146 22992 34152 23044
rect 34204 22992 34210 23044
rect 45526 23004 49280 23032
rect 29604 22936 31340 22964
rect 29604 22924 29610 22936
rect 31478 22924 31484 22976
rect 31536 22924 31542 22976
rect 32766 22924 32772 22976
rect 32824 22924 32830 22976
rect 33502 22924 33508 22976
rect 33560 22924 33566 22976
rect 34238 22924 34244 22976
rect 34296 22924 34302 22976
rect 42794 22924 42800 22976
rect 42852 22964 42858 22976
rect 45526 22964 45554 23004
rect 42852 22936 45554 22964
rect 42852 22924 42858 22936
rect 48406 22924 48412 22976
rect 48464 22924 48470 22976
rect 49252 22973 49280 23004
rect 49237 22967 49295 22973
rect 49237 22933 49249 22967
rect 49283 22933 49295 22967
rect 49237 22927 49295 22933
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 14458 22760 14464 22772
rect 2746 22732 14464 22760
rect 1762 22652 1768 22704
rect 1820 22692 1826 22704
rect 2746 22692 2774 22732
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 19702 22760 19708 22772
rect 16868 22732 19708 22760
rect 1820 22664 2774 22692
rect 3789 22695 3847 22701
rect 1820 22652 1826 22664
rect 3789 22661 3801 22695
rect 3835 22692 3847 22695
rect 3835 22664 6868 22692
rect 3835 22661 3847 22664
rect 3789 22655 3847 22661
rect 1670 22584 1676 22636
rect 1728 22584 1734 22636
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22593 4767 22627
rect 6840 22624 6868 22664
rect 6914 22652 6920 22704
rect 6972 22692 6978 22704
rect 7101 22695 7159 22701
rect 7101 22692 7113 22695
rect 6972 22664 7113 22692
rect 6972 22652 6978 22664
rect 7101 22661 7113 22664
rect 7147 22692 7159 22695
rect 7929 22695 7987 22701
rect 7929 22692 7941 22695
rect 7147 22664 7941 22692
rect 7147 22661 7159 22664
rect 7101 22655 7159 22661
rect 7929 22661 7941 22664
rect 7975 22661 7987 22695
rect 7929 22655 7987 22661
rect 10686 22652 10692 22704
rect 10744 22652 10750 22704
rect 11882 22652 11888 22704
rect 11940 22692 11946 22704
rect 12618 22692 12624 22704
rect 11940 22664 12624 22692
rect 11940 22652 11946 22664
rect 12618 22652 12624 22664
rect 12676 22652 12682 22704
rect 16114 22652 16120 22704
rect 16172 22652 16178 22704
rect 7006 22624 7012 22636
rect 6840 22596 7012 22624
rect 4709 22587 4767 22593
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 2866 22556 2872 22568
rect 2823 22528 2872 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 3694 22516 3700 22568
rect 3752 22556 3758 22568
rect 3881 22559 3939 22565
rect 3881 22556 3893 22559
rect 3752 22528 3893 22556
rect 3752 22516 3758 22528
rect 3881 22525 3893 22528
rect 3927 22525 3939 22559
rect 3881 22519 3939 22525
rect 4065 22559 4123 22565
rect 4065 22525 4077 22559
rect 4111 22556 4123 22559
rect 4246 22556 4252 22568
rect 4111 22528 4252 22556
rect 4111 22525 4123 22528
rect 4065 22519 4123 22525
rect 4246 22516 4252 22528
rect 4304 22516 4310 22568
rect 3510 22448 3516 22500
rect 3568 22488 3574 22500
rect 4724 22488 4752 22587
rect 7006 22584 7012 22596
rect 7064 22584 7070 22636
rect 7193 22627 7251 22633
rect 7193 22593 7205 22627
rect 7239 22624 7251 22627
rect 7834 22624 7840 22636
rect 7239 22596 7840 22624
rect 7239 22593 7251 22596
rect 7193 22587 7251 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 8113 22627 8171 22633
rect 8113 22593 8125 22627
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 7374 22516 7380 22568
rect 7432 22516 7438 22568
rect 3568 22460 4752 22488
rect 3568 22448 3574 22460
rect 5350 22448 5356 22500
rect 5408 22488 5414 22500
rect 8128 22488 8156 22587
rect 9950 22584 9956 22636
rect 10008 22584 10014 22636
rect 11793 22627 11851 22633
rect 11793 22593 11805 22627
rect 11839 22624 11851 22627
rect 11974 22624 11980 22636
rect 11839 22596 11980 22624
rect 11839 22593 11851 22596
rect 11793 22587 11851 22593
rect 11974 22584 11980 22596
rect 12032 22584 12038 22636
rect 13814 22584 13820 22636
rect 13872 22584 13878 22636
rect 15105 22627 15163 22633
rect 15105 22593 15117 22627
rect 15151 22624 15163 22627
rect 16574 22624 16580 22636
rect 15151 22596 16580 22624
rect 15151 22593 15163 22596
rect 15105 22587 15163 22593
rect 16574 22584 16580 22596
rect 16632 22584 16638 22636
rect 16868 22633 16896 22732
rect 19702 22720 19708 22732
rect 19760 22720 19766 22772
rect 20346 22720 20352 22772
rect 20404 22760 20410 22772
rect 21453 22763 21511 22769
rect 21453 22760 21465 22763
rect 20404 22732 21465 22760
rect 20404 22720 20410 22732
rect 21453 22729 21465 22732
rect 21499 22760 21511 22763
rect 25130 22760 25136 22772
rect 21499 22732 25136 22760
rect 21499 22729 21511 22732
rect 21453 22723 21511 22729
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 25777 22763 25835 22769
rect 25777 22729 25789 22763
rect 25823 22760 25835 22763
rect 26142 22760 26148 22772
rect 25823 22732 26148 22760
rect 25823 22729 25835 22732
rect 25777 22723 25835 22729
rect 26142 22720 26148 22732
rect 26200 22720 26206 22772
rect 27614 22720 27620 22772
rect 27672 22720 27678 22772
rect 31478 22760 31484 22772
rect 28644 22732 31484 22760
rect 18506 22692 18512 22704
rect 18354 22664 18512 22692
rect 18506 22652 18512 22664
rect 18564 22652 18570 22704
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 19150 22584 19156 22636
rect 19208 22624 19214 22636
rect 19720 22633 19748 22720
rect 19981 22695 20039 22701
rect 19981 22661 19993 22695
rect 20027 22692 20039 22695
rect 20070 22692 20076 22704
rect 20027 22664 20076 22692
rect 20027 22661 20039 22664
rect 19981 22655 20039 22661
rect 20070 22652 20076 22664
rect 20128 22652 20134 22704
rect 23658 22692 23664 22704
rect 22664 22664 23664 22692
rect 19245 22627 19303 22633
rect 19245 22624 19257 22627
rect 19208 22596 19257 22624
rect 19208 22584 19214 22596
rect 19245 22593 19257 22596
rect 19291 22593 19303 22627
rect 19245 22587 19303 22593
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22593 19763 22627
rect 21450 22624 21456 22636
rect 21114 22596 21456 22624
rect 19705 22587 19763 22593
rect 21450 22584 21456 22596
rect 21508 22584 21514 22636
rect 22664 22633 22692 22664
rect 23658 22652 23664 22664
rect 23716 22652 23722 22704
rect 24670 22652 24676 22704
rect 24728 22692 24734 22704
rect 24728 22664 26004 22692
rect 24728 22652 24734 22664
rect 22649 22627 22707 22633
rect 22649 22593 22661 22627
rect 22695 22593 22707 22627
rect 22649 22587 22707 22593
rect 24486 22584 24492 22636
rect 24544 22624 24550 22636
rect 25222 22624 25228 22636
rect 24544 22596 25228 22624
rect 24544 22584 24550 22596
rect 25222 22584 25228 22596
rect 25280 22584 25286 22636
rect 25498 22584 25504 22636
rect 25556 22624 25562 22636
rect 25685 22627 25743 22633
rect 25685 22624 25697 22627
rect 25556 22596 25697 22624
rect 25556 22584 25562 22596
rect 25685 22593 25697 22596
rect 25731 22593 25743 22627
rect 25685 22587 25743 22593
rect 8662 22516 8668 22568
rect 8720 22516 8726 22568
rect 12434 22516 12440 22568
rect 12492 22516 12498 22568
rect 13832 22556 13860 22584
rect 17129 22559 17187 22565
rect 12544 22528 14320 22556
rect 5408 22460 8156 22488
rect 5408 22448 5414 22460
rect 10502 22448 10508 22500
rect 10560 22488 10566 22500
rect 10778 22488 10784 22500
rect 10560 22460 10784 22488
rect 10560 22448 10566 22460
rect 10778 22448 10784 22460
rect 10836 22488 10842 22500
rect 12544 22488 12572 22528
rect 10836 22460 12572 22488
rect 10836 22448 10842 22460
rect 3418 22380 3424 22432
rect 3476 22380 3482 22432
rect 3602 22380 3608 22432
rect 3660 22420 3666 22432
rect 4522 22420 4528 22432
rect 3660 22392 4528 22420
rect 3660 22380 3666 22392
rect 4522 22380 4528 22392
rect 4580 22380 4586 22432
rect 6638 22380 6644 22432
rect 6696 22420 6702 22432
rect 6733 22423 6791 22429
rect 6733 22420 6745 22423
rect 6696 22392 6745 22420
rect 6696 22380 6702 22392
rect 6733 22389 6745 22392
rect 6779 22389 6791 22423
rect 6733 22383 6791 22389
rect 6822 22380 6828 22432
rect 6880 22420 6886 22432
rect 11885 22423 11943 22429
rect 11885 22420 11897 22423
rect 6880 22392 11897 22420
rect 6880 22380 6886 22392
rect 11885 22389 11897 22392
rect 11931 22389 11943 22423
rect 11885 22383 11943 22389
rect 12250 22380 12256 22432
rect 12308 22420 12314 22432
rect 12694 22423 12752 22429
rect 12694 22420 12706 22423
rect 12308 22392 12706 22420
rect 12308 22380 12314 22392
rect 12694 22389 12706 22392
rect 12740 22420 12752 22423
rect 13170 22420 13176 22432
rect 12740 22392 13176 22420
rect 12740 22389 12752 22392
rect 12694 22383 12752 22389
rect 13170 22380 13176 22392
rect 13228 22380 13234 22432
rect 13446 22380 13452 22432
rect 13504 22420 13510 22432
rect 14185 22423 14243 22429
rect 14185 22420 14197 22423
rect 13504 22392 14197 22420
rect 13504 22380 13510 22392
rect 14185 22389 14197 22392
rect 14231 22389 14243 22423
rect 14292 22420 14320 22528
rect 17129 22525 17141 22559
rect 17175 22556 17187 22559
rect 17218 22556 17224 22568
rect 17175 22528 17224 22556
rect 17175 22525 17187 22528
rect 17129 22519 17187 22525
rect 17218 22516 17224 22528
rect 17276 22516 17282 22568
rect 18598 22516 18604 22568
rect 18656 22516 18662 22568
rect 22278 22516 22284 22568
rect 22336 22556 22342 22568
rect 23109 22559 23167 22565
rect 23109 22556 23121 22559
rect 22336 22528 23121 22556
rect 22336 22516 22342 22528
rect 23109 22525 23121 22528
rect 23155 22525 23167 22559
rect 23109 22519 23167 22525
rect 18506 22420 18512 22432
rect 14292 22392 18512 22420
rect 14185 22383 14243 22389
rect 18506 22380 18512 22392
rect 18564 22380 18570 22432
rect 19058 22380 19064 22432
rect 19116 22380 19122 22432
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 21818 22420 21824 22432
rect 19392 22392 21824 22420
rect 19392 22380 19398 22392
rect 21818 22380 21824 22392
rect 21876 22380 21882 22432
rect 23124 22420 23152 22519
rect 23382 22516 23388 22568
rect 23440 22516 23446 22568
rect 23474 22516 23480 22568
rect 23532 22556 23538 22568
rect 24578 22556 24584 22568
rect 23532 22528 24584 22556
rect 23532 22516 23538 22528
rect 24578 22516 24584 22528
rect 24636 22516 24642 22568
rect 25869 22559 25927 22565
rect 25869 22556 25881 22559
rect 24872 22528 25881 22556
rect 23382 22420 23388 22432
rect 23124 22392 23388 22420
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 23934 22380 23940 22432
rect 23992 22420 23998 22432
rect 24872 22429 24900 22528
rect 25869 22525 25881 22528
rect 25915 22525 25927 22559
rect 25869 22519 25927 22525
rect 25976 22488 26004 22664
rect 27430 22652 27436 22704
rect 27488 22692 27494 22704
rect 28644 22701 28672 22732
rect 31478 22720 31484 22732
rect 31536 22720 31542 22772
rect 32490 22720 32496 22772
rect 32548 22720 32554 22772
rect 28629 22695 28687 22701
rect 27488 22664 27752 22692
rect 27488 22652 27494 22664
rect 27338 22624 27344 22636
rect 26068 22596 27344 22624
rect 26068 22568 26096 22596
rect 27338 22584 27344 22596
rect 27396 22624 27402 22636
rect 27525 22627 27583 22633
rect 27525 22624 27537 22627
rect 27396 22596 27537 22624
rect 27396 22584 27402 22596
rect 27525 22593 27537 22596
rect 27571 22593 27583 22627
rect 27525 22587 27583 22593
rect 26050 22516 26056 22568
rect 26108 22516 26114 22568
rect 26142 22516 26148 22568
rect 26200 22556 26206 22568
rect 27724 22565 27752 22664
rect 28629 22661 28641 22695
rect 28675 22661 28687 22695
rect 30006 22692 30012 22704
rect 29854 22664 30012 22692
rect 28629 22655 28687 22661
rect 30006 22652 30012 22664
rect 30064 22652 30070 22704
rect 31018 22652 31024 22704
rect 31076 22652 31082 22704
rect 31110 22652 31116 22704
rect 31168 22692 31174 22704
rect 40034 22692 40040 22704
rect 31168 22664 35894 22692
rect 39422 22664 40040 22692
rect 31168 22652 31174 22664
rect 28350 22584 28356 22636
rect 28408 22584 28414 22636
rect 30926 22584 30932 22636
rect 30984 22584 30990 22636
rect 32398 22584 32404 22636
rect 32456 22584 32462 22636
rect 33137 22627 33195 22633
rect 33137 22593 33149 22627
rect 33183 22624 33195 22627
rect 33318 22624 33324 22636
rect 33183 22596 33324 22624
rect 33183 22593 33195 22596
rect 33137 22587 33195 22593
rect 33318 22584 33324 22596
rect 33376 22584 33382 22636
rect 33502 22584 33508 22636
rect 33560 22624 33566 22636
rect 34241 22627 34299 22633
rect 34241 22624 34253 22627
rect 33560 22596 34253 22624
rect 33560 22584 33566 22596
rect 34241 22593 34253 22596
rect 34287 22593 34299 22627
rect 35866 22624 35894 22664
rect 40034 22652 40040 22664
rect 40092 22652 40098 22704
rect 37921 22627 37979 22633
rect 37921 22624 37933 22627
rect 35866 22596 37933 22624
rect 34241 22587 34299 22593
rect 37921 22593 37933 22596
rect 37967 22593 37979 22627
rect 37921 22587 37979 22593
rect 27709 22559 27767 22565
rect 26200 22528 27568 22556
rect 26200 22516 26206 22528
rect 27157 22491 27215 22497
rect 27157 22488 27169 22491
rect 25976 22460 27169 22488
rect 27157 22457 27169 22460
rect 27203 22457 27215 22491
rect 27540 22488 27568 22528
rect 27709 22525 27721 22559
rect 27755 22525 27767 22559
rect 27709 22519 27767 22525
rect 28718 22516 28724 22568
rect 28776 22556 28782 22568
rect 31113 22559 31171 22565
rect 31113 22556 31125 22559
rect 28776 22528 31125 22556
rect 28776 22516 28782 22528
rect 31113 22525 31125 22528
rect 31159 22525 31171 22559
rect 31113 22519 31171 22525
rect 38197 22559 38255 22565
rect 38197 22525 38209 22559
rect 38243 22556 38255 22559
rect 48406 22556 48412 22568
rect 38243 22528 48412 22556
rect 38243 22525 38255 22528
rect 38197 22519 38255 22525
rect 48406 22516 48412 22528
rect 48464 22516 48470 22568
rect 27798 22488 27804 22500
rect 27540 22460 27804 22488
rect 27157 22451 27215 22457
rect 27798 22448 27804 22460
rect 27856 22448 27862 22500
rect 29914 22448 29920 22500
rect 29972 22488 29978 22500
rect 29972 22460 30236 22488
rect 29972 22448 29978 22460
rect 24857 22423 24915 22429
rect 24857 22420 24869 22423
rect 23992 22392 24869 22420
rect 23992 22380 23998 22392
rect 24857 22389 24869 22392
rect 24903 22389 24915 22423
rect 24857 22383 24915 22389
rect 25314 22380 25320 22432
rect 25372 22380 25378 22432
rect 25406 22380 25412 22432
rect 25464 22420 25470 22432
rect 26602 22420 26608 22432
rect 25464 22392 26608 22420
rect 25464 22380 25470 22392
rect 26602 22380 26608 22392
rect 26660 22380 26666 22432
rect 28994 22380 29000 22432
rect 29052 22420 29058 22432
rect 30101 22423 30159 22429
rect 30101 22420 30113 22423
rect 29052 22392 30113 22420
rect 29052 22380 29058 22392
rect 30101 22389 30113 22392
rect 30147 22389 30159 22423
rect 30208 22420 30236 22460
rect 30374 22448 30380 22500
rect 30432 22488 30438 22500
rect 30561 22491 30619 22497
rect 30561 22488 30573 22491
rect 30432 22460 30573 22488
rect 30432 22448 30438 22460
rect 30561 22457 30573 22460
rect 30607 22457 30619 22491
rect 30561 22451 30619 22457
rect 31662 22448 31668 22500
rect 31720 22488 31726 22500
rect 33965 22491 34023 22497
rect 33965 22488 33977 22491
rect 31720 22460 33977 22488
rect 31720 22448 31726 22460
rect 33965 22457 33977 22460
rect 34011 22488 34023 22491
rect 34701 22491 34759 22497
rect 34701 22488 34713 22491
rect 34011 22460 34713 22488
rect 34011 22457 34023 22460
rect 33965 22451 34023 22457
rect 34701 22457 34713 22460
rect 34747 22457 34759 22491
rect 34701 22451 34759 22457
rect 31570 22420 31576 22432
rect 30208 22392 31576 22420
rect 30101 22383 30159 22389
rect 31570 22380 31576 22392
rect 31628 22380 31634 22432
rect 33226 22380 33232 22432
rect 33284 22380 33290 22432
rect 34330 22380 34336 22432
rect 34388 22380 34394 22432
rect 39666 22380 39672 22432
rect 39724 22380 39730 22432
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 3602 22176 3608 22228
rect 3660 22216 3666 22228
rect 3786 22216 3792 22228
rect 3660 22188 3792 22216
rect 3660 22176 3666 22188
rect 3786 22176 3792 22188
rect 3844 22176 3850 22228
rect 6546 22176 6552 22228
rect 6604 22216 6610 22228
rect 6822 22216 6828 22228
rect 6604 22188 6828 22216
rect 6604 22176 6610 22188
rect 6822 22176 6828 22188
rect 6880 22176 6886 22228
rect 7006 22176 7012 22228
rect 7064 22216 7070 22228
rect 10318 22216 10324 22228
rect 7064 22188 10324 22216
rect 7064 22176 7070 22188
rect 10318 22176 10324 22188
rect 10376 22176 10382 22228
rect 14458 22176 14464 22228
rect 14516 22176 14522 22228
rect 19518 22216 19524 22228
rect 16546 22188 19524 22216
rect 6730 22108 6736 22160
rect 6788 22148 6794 22160
rect 10962 22148 10968 22160
rect 6788 22120 6914 22148
rect 6788 22108 6794 22120
rect 1302 22040 1308 22092
rect 1360 22080 1366 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1360 22052 2053 22080
rect 1360 22040 1366 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 4430 22040 4436 22092
rect 4488 22040 4494 22092
rect 6886 22080 6914 22120
rect 9968 22120 10968 22148
rect 9968 22089 9996 22120
rect 10962 22108 10968 22120
rect 11020 22108 11026 22160
rect 15102 22108 15108 22160
rect 15160 22148 15166 22160
rect 15160 22120 15700 22148
rect 15160 22108 15166 22120
rect 7285 22083 7343 22089
rect 7285 22080 7297 22083
rect 6886 22052 7297 22080
rect 7285 22049 7297 22052
rect 7331 22049 7343 22083
rect 7285 22043 7343 22049
rect 9953 22083 10011 22089
rect 9953 22049 9965 22083
rect 9999 22080 10011 22083
rect 9999 22052 10033 22080
rect 9999 22049 10011 22052
rect 9953 22043 10011 22049
rect 10594 22040 10600 22092
rect 10652 22040 10658 22092
rect 13354 22040 13360 22092
rect 13412 22040 13418 22092
rect 15672 22089 15700 22120
rect 15657 22083 15715 22089
rect 15657 22049 15669 22083
rect 15703 22049 15715 22083
rect 15657 22043 15715 22049
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 22012 1823 22015
rect 1811 21984 2268 22012
rect 1811 21981 1823 21984
rect 1765 21975 1823 21981
rect 2240 21876 2268 21984
rect 2314 21972 2320 22024
rect 2372 22012 2378 22024
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 2372 21984 3985 22012
rect 2372 21972 2378 21984
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 7006 21972 7012 22024
rect 7064 21972 7070 22024
rect 9677 22015 9735 22021
rect 9677 21981 9689 22015
rect 9723 22012 9735 22015
rect 10612 22012 10640 22040
rect 9723 21984 10640 22012
rect 10873 22015 10931 22021
rect 9723 21981 9735 21984
rect 9677 21975 9735 21981
rect 10873 21981 10885 22015
rect 10919 22012 10931 22015
rect 11146 22012 11152 22024
rect 10919 21984 11152 22012
rect 10919 21981 10931 21984
rect 10873 21975 10931 21981
rect 11146 21972 11152 21984
rect 11204 21972 11210 22024
rect 11238 21972 11244 22024
rect 11296 22012 11302 22024
rect 11609 22015 11667 22021
rect 11609 22012 11621 22015
rect 11296 21984 11621 22012
rect 11296 21972 11302 21984
rect 11609 21981 11621 21984
rect 11655 21981 11667 22015
rect 11609 21975 11667 21981
rect 12526 21972 12532 22024
rect 12584 21972 12590 22024
rect 15381 22015 15439 22021
rect 15381 21981 15393 22015
rect 15427 22012 15439 22015
rect 16546 22012 16574 22188
rect 19518 22176 19524 22188
rect 19576 22176 19582 22228
rect 19978 22176 19984 22228
rect 20036 22216 20042 22228
rect 32766 22216 32772 22228
rect 20036 22188 32772 22216
rect 20036 22176 20042 22188
rect 32766 22176 32772 22188
rect 32824 22176 32830 22228
rect 18874 22108 18880 22160
rect 18932 22148 18938 22160
rect 19334 22148 19340 22160
rect 18932 22120 19340 22148
rect 18932 22108 18938 22120
rect 19334 22108 19340 22120
rect 19392 22108 19398 22160
rect 22830 22108 22836 22160
rect 22888 22108 22894 22160
rect 25406 22148 25412 22160
rect 23952 22120 25412 22148
rect 17126 22040 17132 22092
rect 17184 22080 17190 22092
rect 18690 22080 18696 22092
rect 17184 22052 18696 22080
rect 17184 22040 17190 22052
rect 18690 22040 18696 22052
rect 18748 22040 18754 22092
rect 20162 22080 20168 22092
rect 18984 22052 20168 22080
rect 15427 21984 16574 22012
rect 15427 21981 15439 21984
rect 15381 21975 15439 21981
rect 18506 21972 18512 22024
rect 18564 22012 18570 22024
rect 18984 22012 19012 22052
rect 20162 22040 20168 22052
rect 20220 22040 20226 22092
rect 20254 22040 20260 22092
rect 20312 22080 20318 22092
rect 23952 22089 23980 22120
rect 25406 22108 25412 22120
rect 25464 22108 25470 22160
rect 27062 22108 27068 22160
rect 27120 22148 27126 22160
rect 28169 22151 28227 22157
rect 28169 22148 28181 22151
rect 27120 22120 28181 22148
rect 27120 22108 27126 22120
rect 28169 22117 28181 22120
rect 28215 22117 28227 22151
rect 31478 22148 31484 22160
rect 28169 22111 28227 22117
rect 30760 22120 31484 22148
rect 20809 22083 20867 22089
rect 20809 22080 20821 22083
rect 20312 22052 20821 22080
rect 20312 22040 20318 22052
rect 20809 22049 20821 22052
rect 20855 22049 20867 22083
rect 20809 22043 20867 22049
rect 23937 22083 23995 22089
rect 23937 22049 23949 22083
rect 23983 22080 23995 22083
rect 23983 22052 24017 22080
rect 23983 22049 23995 22052
rect 23937 22043 23995 22049
rect 25130 22040 25136 22092
rect 25188 22040 25194 22092
rect 27246 22040 27252 22092
rect 27304 22040 27310 22092
rect 27430 22040 27436 22092
rect 27488 22080 27494 22092
rect 27525 22083 27583 22089
rect 27525 22080 27537 22083
rect 27488 22052 27537 22080
rect 27488 22040 27494 22052
rect 27525 22049 27537 22052
rect 27571 22049 27583 22083
rect 29178 22080 29184 22092
rect 27525 22043 27583 22049
rect 27632 22052 29184 22080
rect 18564 21984 19012 22012
rect 18564 21972 18570 21984
rect 19058 21972 19064 22024
rect 19116 22012 19122 22024
rect 19288 22012 19294 22024
rect 19116 21984 19294 22012
rect 19116 21972 19122 21984
rect 19288 21972 19294 21984
rect 19346 21972 19352 22024
rect 19610 21972 19616 22024
rect 19668 22012 19674 22024
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 19668 22008 19748 22012
rect 19904 22008 20361 22012
rect 19668 21984 20361 22008
rect 19668 21972 19674 21984
rect 19720 21980 19932 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 23382 21972 23388 22024
rect 23440 22012 23446 22024
rect 24854 22012 24860 22024
rect 23440 21984 24860 22012
rect 23440 21972 23446 21984
rect 24854 21972 24860 21984
rect 24912 22012 24918 22024
rect 25774 22012 25780 22024
rect 24912 21984 25780 22012
rect 24912 21972 24918 21984
rect 25774 21972 25780 21984
rect 25832 21972 25838 22024
rect 27264 22012 27292 22040
rect 27632 22012 27660 22052
rect 29178 22040 29184 22052
rect 29236 22080 29242 22092
rect 29638 22080 29644 22092
rect 29236 22052 29644 22080
rect 29236 22040 29242 22052
rect 29638 22040 29644 22052
rect 29696 22040 29702 22092
rect 30760 22089 30788 22120
rect 31478 22108 31484 22120
rect 31536 22108 31542 22160
rect 31570 22108 31576 22160
rect 31628 22148 31634 22160
rect 39666 22148 39672 22160
rect 31628 22120 39672 22148
rect 31628 22108 31634 22120
rect 39666 22108 39672 22120
rect 39724 22108 39730 22160
rect 30745 22083 30803 22089
rect 30745 22049 30757 22083
rect 30791 22080 30803 22083
rect 34514 22080 34520 22092
rect 30791 22052 30825 22080
rect 32508 22052 34520 22080
rect 30791 22049 30803 22052
rect 30745 22043 30803 22049
rect 27264 21984 27660 22012
rect 27798 21972 27804 22024
rect 27856 22012 27862 22024
rect 28813 22015 28871 22021
rect 28813 22012 28825 22015
rect 27856 21984 28825 22012
rect 27856 21972 27862 21984
rect 28813 21981 28825 21984
rect 28859 21981 28871 22015
rect 28813 21975 28871 21981
rect 30561 22015 30619 22021
rect 30561 21981 30573 22015
rect 30607 22012 30619 22015
rect 32508 22012 32536 22052
rect 34514 22040 34520 22052
rect 34572 22040 34578 22092
rect 30607 21984 32536 22012
rect 30607 21981 30619 21984
rect 30561 21975 30619 21981
rect 32582 21972 32588 22024
rect 32640 21972 32646 22024
rect 32858 21972 32864 22024
rect 32916 21972 32922 22024
rect 49050 21972 49056 22024
rect 49108 21972 49114 22024
rect 6181 21947 6239 21953
rect 6181 21913 6193 21947
rect 6227 21944 6239 21947
rect 6454 21944 6460 21956
rect 6227 21916 6460 21944
rect 6227 21913 6239 21916
rect 6181 21907 6239 21913
rect 6454 21904 6460 21916
rect 6512 21904 6518 21956
rect 9769 21947 9827 21953
rect 9769 21913 9781 21947
rect 9815 21944 9827 21947
rect 11882 21944 11888 21956
rect 9815 21916 11888 21944
rect 9815 21913 9827 21916
rect 9769 21907 9827 21913
rect 11882 21904 11888 21916
rect 11940 21904 11946 21956
rect 14366 21904 14372 21956
rect 14424 21904 14430 21956
rect 16666 21904 16672 21956
rect 16724 21944 16730 21956
rect 17405 21947 17463 21953
rect 17405 21944 17417 21947
rect 16724 21916 17417 21944
rect 16724 21904 16730 21916
rect 17405 21913 17417 21916
rect 17451 21944 17463 21947
rect 17494 21944 17500 21956
rect 17451 21916 17500 21944
rect 17451 21913 17463 21916
rect 17405 21907 17463 21913
rect 17494 21904 17500 21916
rect 17552 21904 17558 21956
rect 18782 21904 18788 21956
rect 18840 21944 18846 21956
rect 19485 21947 19543 21953
rect 19485 21944 19497 21947
rect 18840 21916 19497 21944
rect 18840 21904 18846 21916
rect 19485 21913 19497 21916
rect 19531 21913 19543 21947
rect 19485 21907 19543 21913
rect 20530 21904 20536 21956
rect 20588 21944 20594 21956
rect 23474 21944 23480 21956
rect 20588 21916 23480 21944
rect 20588 21904 20594 21916
rect 23474 21904 23480 21916
rect 23532 21904 23538 21956
rect 23658 21904 23664 21956
rect 23716 21904 23722 21956
rect 23753 21947 23811 21953
rect 23753 21913 23765 21947
rect 23799 21944 23811 21947
rect 24670 21944 24676 21956
rect 23799 21916 24676 21944
rect 23799 21913 23811 21916
rect 23753 21907 23811 21913
rect 24670 21904 24676 21916
rect 24728 21904 24734 21956
rect 24949 21947 25007 21953
rect 24949 21913 24961 21947
rect 24995 21944 25007 21947
rect 25682 21944 25688 21956
rect 24995 21916 25688 21944
rect 24995 21913 25007 21916
rect 24949 21907 25007 21913
rect 25682 21904 25688 21916
rect 25740 21904 25746 21956
rect 25958 21904 25964 21956
rect 26016 21944 26022 21956
rect 26053 21947 26111 21953
rect 26053 21944 26065 21947
rect 26016 21916 26065 21944
rect 26016 21904 26022 21916
rect 26053 21913 26065 21916
rect 26099 21913 26111 21947
rect 26053 21907 26111 21913
rect 26786 21904 26792 21956
rect 26844 21904 26850 21956
rect 27448 21916 28672 21944
rect 5994 21876 6000 21888
rect 2240 21848 6000 21876
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 6270 21836 6276 21888
rect 6328 21836 6334 21888
rect 8938 21836 8944 21888
rect 8996 21876 9002 21888
rect 9309 21879 9367 21885
rect 9309 21876 9321 21879
rect 8996 21848 9321 21876
rect 8996 21836 9002 21848
rect 9309 21845 9321 21848
rect 9355 21845 9367 21879
rect 9309 21839 9367 21845
rect 9398 21836 9404 21888
rect 9456 21876 9462 21888
rect 14918 21876 14924 21888
rect 9456 21848 14924 21876
rect 9456 21836 9462 21848
rect 14918 21836 14924 21848
rect 14976 21836 14982 21888
rect 15010 21836 15016 21888
rect 15068 21836 15074 21888
rect 17218 21836 17224 21888
rect 17276 21876 17282 21888
rect 18877 21879 18935 21885
rect 18877 21876 18889 21879
rect 17276 21848 18889 21876
rect 17276 21836 17282 21848
rect 18877 21845 18889 21848
rect 18923 21845 18935 21879
rect 18877 21839 18935 21845
rect 18966 21836 18972 21888
rect 19024 21876 19030 21888
rect 19334 21876 19340 21888
rect 19024 21848 19340 21876
rect 19024 21836 19030 21848
rect 19334 21836 19340 21848
rect 19392 21836 19398 21888
rect 19613 21879 19671 21885
rect 19613 21845 19625 21879
rect 19659 21876 19671 21879
rect 20070 21876 20076 21888
rect 19659 21848 20076 21876
rect 19659 21845 19671 21848
rect 19613 21839 19671 21845
rect 20070 21836 20076 21848
rect 20128 21836 20134 21888
rect 23290 21836 23296 21888
rect 23348 21836 23354 21888
rect 23566 21836 23572 21888
rect 23624 21876 23630 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 23624 21848 24593 21876
rect 23624 21836 23630 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 25041 21879 25099 21885
rect 25041 21845 25053 21879
rect 25087 21876 25099 21879
rect 27448 21876 27476 21916
rect 28644 21885 28672 21916
rect 29178 21904 29184 21956
rect 29236 21944 29242 21956
rect 31389 21947 31447 21953
rect 31389 21944 31401 21947
rect 29236 21916 31401 21944
rect 29236 21904 29242 21916
rect 31389 21913 31401 21916
rect 31435 21913 31447 21947
rect 31389 21907 31447 21913
rect 25087 21848 27476 21876
rect 28629 21879 28687 21885
rect 25087 21845 25099 21848
rect 25041 21839 25099 21845
rect 28629 21845 28641 21879
rect 28675 21845 28687 21879
rect 28629 21839 28687 21845
rect 28994 21836 29000 21888
rect 29052 21876 29058 21888
rect 30101 21879 30159 21885
rect 30101 21876 30113 21879
rect 29052 21848 30113 21876
rect 29052 21836 29058 21848
rect 30101 21845 30113 21848
rect 30147 21845 30159 21879
rect 30101 21839 30159 21845
rect 30469 21879 30527 21885
rect 30469 21845 30481 21879
rect 30515 21876 30527 21879
rect 31294 21876 31300 21888
rect 30515 21848 31300 21876
rect 30515 21845 30527 21848
rect 30469 21839 30527 21845
rect 31294 21836 31300 21848
rect 31352 21836 31358 21888
rect 31478 21836 31484 21888
rect 31536 21836 31542 21888
rect 49234 21836 49240 21888
rect 49292 21836 49298 21888
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 1762 21632 1768 21684
rect 1820 21672 1826 21684
rect 6270 21672 6276 21684
rect 1820 21644 6276 21672
rect 1820 21632 1826 21644
rect 6270 21632 6276 21644
rect 6328 21632 6334 21684
rect 6380 21644 9720 21672
rect 2130 21564 2136 21616
rect 2188 21604 2194 21616
rect 5721 21607 5779 21613
rect 5721 21604 5733 21607
rect 2188 21576 5733 21604
rect 2188 21564 2194 21576
rect 5721 21573 5733 21576
rect 5767 21573 5779 21607
rect 5721 21567 5779 21573
rect 6086 21564 6092 21616
rect 6144 21604 6150 21616
rect 6380 21604 6408 21644
rect 6144 21576 6408 21604
rect 6144 21564 6150 21576
rect 6730 21564 6736 21616
rect 6788 21604 6794 21616
rect 7374 21604 7380 21616
rect 6788 21576 7380 21604
rect 6788 21564 6794 21576
rect 7374 21564 7380 21576
rect 7432 21564 7438 21616
rect 9582 21604 9588 21616
rect 8602 21576 9588 21604
rect 9582 21564 9588 21576
rect 9640 21564 9646 21616
rect 9692 21604 9720 21644
rect 11882 21632 11888 21684
rect 11940 21632 11946 21684
rect 12345 21675 12403 21681
rect 12345 21641 12357 21675
rect 12391 21672 12403 21675
rect 12802 21672 12808 21684
rect 12391 21644 12808 21672
rect 12391 21641 12403 21644
rect 12345 21635 12403 21641
rect 12802 21632 12808 21644
rect 12860 21632 12866 21684
rect 18782 21672 18788 21684
rect 13464 21644 18788 21672
rect 12253 21607 12311 21613
rect 12253 21604 12265 21607
rect 9692 21576 12265 21604
rect 12253 21573 12265 21576
rect 12299 21573 12311 21607
rect 13464 21604 13492 21644
rect 18782 21632 18788 21644
rect 18840 21632 18846 21684
rect 19702 21672 19708 21684
rect 18892 21644 19708 21672
rect 12253 21567 12311 21573
rect 12360 21576 13492 21604
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21536 1823 21539
rect 2314 21536 2320 21548
rect 1811 21508 2320 21536
rect 1811 21505 1823 21508
rect 1765 21499 1823 21505
rect 2314 21496 2320 21508
rect 2372 21496 2378 21548
rect 3602 21496 3608 21548
rect 3660 21496 3666 21548
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21536 5687 21539
rect 5675 21508 6776 21536
rect 5675 21505 5687 21508
rect 5629 21499 5687 21505
rect 2038 21428 2044 21480
rect 2096 21428 2102 21480
rect 4154 21428 4160 21480
rect 4212 21428 4218 21480
rect 5534 21428 5540 21480
rect 5592 21468 5598 21480
rect 5813 21471 5871 21477
rect 5813 21468 5825 21471
rect 5592 21440 5825 21468
rect 5592 21428 5598 21440
rect 5813 21437 5825 21440
rect 5859 21437 5871 21471
rect 6748 21468 6776 21508
rect 6822 21496 6828 21548
rect 6880 21496 6886 21548
rect 9306 21496 9312 21548
rect 9364 21536 9370 21548
rect 10229 21539 10287 21545
rect 10229 21536 10241 21539
rect 9364 21508 10241 21536
rect 9364 21496 9370 21508
rect 10229 21505 10241 21508
rect 10275 21505 10287 21539
rect 10229 21499 10287 21505
rect 10321 21539 10379 21545
rect 10321 21505 10333 21539
rect 10367 21536 10379 21539
rect 12066 21536 12072 21548
rect 10367 21508 12072 21536
rect 10367 21505 10379 21508
rect 10321 21499 10379 21505
rect 12066 21496 12072 21508
rect 12124 21496 12130 21548
rect 6748 21440 6960 21468
rect 5813 21431 5871 21437
rect 1946 21360 1952 21412
rect 2004 21400 2010 21412
rect 6932 21400 6960 21440
rect 7098 21428 7104 21480
rect 7156 21428 7162 21480
rect 9950 21468 9956 21480
rect 7208 21440 9956 21468
rect 7208 21400 7236 21440
rect 9950 21428 9956 21440
rect 10008 21428 10014 21480
rect 10042 21428 10048 21480
rect 10100 21468 10106 21480
rect 10413 21471 10471 21477
rect 10413 21468 10425 21471
rect 10100 21440 10425 21468
rect 10100 21428 10106 21440
rect 10413 21437 10425 21440
rect 10459 21437 10471 21471
rect 10413 21431 10471 21437
rect 10778 21428 10784 21480
rect 10836 21468 10842 21480
rect 12360 21468 12388 21576
rect 14918 21564 14924 21616
rect 14976 21604 14982 21616
rect 18892 21604 18920 21644
rect 19702 21632 19708 21644
rect 19760 21632 19766 21684
rect 20530 21632 20536 21684
rect 20588 21672 20594 21684
rect 25130 21672 25136 21684
rect 20588 21644 25136 21672
rect 20588 21632 20594 21644
rect 25130 21632 25136 21644
rect 25188 21632 25194 21684
rect 25961 21675 26019 21681
rect 25961 21641 25973 21675
rect 26007 21672 26019 21675
rect 26694 21672 26700 21684
rect 26007 21644 26700 21672
rect 26007 21641 26019 21644
rect 25961 21635 26019 21641
rect 26694 21632 26700 21644
rect 26752 21632 26758 21684
rect 26786 21632 26792 21684
rect 26844 21672 26850 21684
rect 27246 21672 27252 21684
rect 26844 21644 27252 21672
rect 26844 21632 26850 21644
rect 27246 21632 27252 21644
rect 27304 21632 27310 21684
rect 27709 21675 27767 21681
rect 27709 21641 27721 21675
rect 27755 21672 27767 21675
rect 27755 21644 30972 21672
rect 27755 21641 27767 21644
rect 27709 21635 27767 21641
rect 20254 21604 20260 21616
rect 14976 21576 18920 21604
rect 20194 21576 20260 21604
rect 14976 21564 14982 21576
rect 20254 21564 20260 21576
rect 20312 21604 20318 21616
rect 21082 21604 21088 21616
rect 20312 21576 21088 21604
rect 20312 21564 20318 21576
rect 21082 21564 21088 21576
rect 21140 21564 21146 21616
rect 23661 21607 23719 21613
rect 23661 21573 23673 21607
rect 23707 21604 23719 21607
rect 23934 21604 23940 21616
rect 23707 21576 23940 21604
rect 23707 21573 23719 21576
rect 23661 21567 23719 21573
rect 23934 21564 23940 21576
rect 23992 21564 23998 21616
rect 25222 21604 25228 21616
rect 24886 21576 25228 21604
rect 25222 21564 25228 21576
rect 25280 21564 25286 21616
rect 28994 21604 29000 21616
rect 26068 21576 29000 21604
rect 12526 21496 12532 21548
rect 12584 21536 12590 21548
rect 12805 21539 12863 21545
rect 12805 21536 12817 21539
rect 12584 21508 12817 21536
rect 12584 21496 12590 21508
rect 12805 21505 12817 21508
rect 12851 21505 12863 21539
rect 14214 21508 14320 21536
rect 12805 21499 12863 21505
rect 14292 21480 14320 21508
rect 15010 21496 15016 21548
rect 15068 21536 15074 21548
rect 15933 21539 15991 21545
rect 15933 21536 15945 21539
rect 15068 21508 15945 21536
rect 15068 21496 15074 21508
rect 15933 21505 15945 21508
rect 15979 21536 15991 21539
rect 15979 21508 16160 21536
rect 15979 21505 15991 21508
rect 15933 21499 15991 21505
rect 10836 21440 12388 21468
rect 12437 21471 12495 21477
rect 10836 21428 10842 21440
rect 12437 21437 12449 21471
rect 12483 21437 12495 21471
rect 12437 21431 12495 21437
rect 13081 21471 13139 21477
rect 13081 21437 13093 21471
rect 13127 21468 13139 21471
rect 13446 21468 13452 21480
rect 13127 21440 13452 21468
rect 13127 21437 13139 21440
rect 13081 21431 13139 21437
rect 2004 21372 5396 21400
rect 6932 21372 7236 21400
rect 8849 21403 8907 21409
rect 2004 21360 2010 21372
rect 1486 21292 1492 21344
rect 1544 21332 1550 21344
rect 3326 21332 3332 21344
rect 1544 21304 3332 21332
rect 1544 21292 1550 21304
rect 3326 21292 3332 21304
rect 3384 21292 3390 21344
rect 4430 21292 4436 21344
rect 4488 21332 4494 21344
rect 5261 21335 5319 21341
rect 5261 21332 5273 21335
rect 4488 21304 5273 21332
rect 4488 21292 4494 21304
rect 5261 21301 5273 21304
rect 5307 21301 5319 21335
rect 5368 21332 5396 21372
rect 8849 21369 8861 21403
rect 8895 21400 8907 21403
rect 9490 21400 9496 21412
rect 8895 21372 9496 21400
rect 8895 21369 8907 21372
rect 8849 21363 8907 21369
rect 9490 21360 9496 21372
rect 9548 21400 9554 21412
rect 12452 21400 12480 21431
rect 13446 21428 13452 21440
rect 13504 21428 13510 21480
rect 13814 21428 13820 21480
rect 13872 21468 13878 21480
rect 14274 21468 14280 21480
rect 13872 21440 14280 21468
rect 13872 21428 13878 21440
rect 14274 21428 14280 21440
rect 14332 21428 14338 21480
rect 15194 21428 15200 21480
rect 15252 21468 15258 21480
rect 16025 21471 16083 21477
rect 16025 21468 16037 21471
rect 15252 21440 16037 21468
rect 15252 21428 15258 21440
rect 16025 21437 16037 21440
rect 16071 21437 16083 21471
rect 16025 21431 16083 21437
rect 9548 21372 12480 21400
rect 9548 21360 9554 21372
rect 6917 21335 6975 21341
rect 6917 21332 6929 21335
rect 5368 21304 6929 21332
rect 5261 21295 5319 21301
rect 6917 21301 6929 21304
rect 6963 21301 6975 21335
rect 6917 21295 6975 21301
rect 7098 21292 7104 21344
rect 7156 21332 7162 21344
rect 8478 21332 8484 21344
rect 7156 21304 8484 21332
rect 7156 21292 7162 21304
rect 8478 21292 8484 21304
rect 8536 21292 8542 21344
rect 9306 21292 9312 21344
rect 9364 21292 9370 21344
rect 9858 21292 9864 21344
rect 9916 21292 9922 21344
rect 9950 21292 9956 21344
rect 10008 21332 10014 21344
rect 10778 21332 10784 21344
rect 10008 21304 10784 21332
rect 10008 21292 10014 21304
rect 10778 21292 10784 21304
rect 10836 21292 10842 21344
rect 12802 21292 12808 21344
rect 12860 21332 12866 21344
rect 13814 21332 13820 21344
rect 12860 21304 13820 21332
rect 12860 21292 12866 21304
rect 13814 21292 13820 21304
rect 13872 21292 13878 21344
rect 14090 21292 14096 21344
rect 14148 21332 14154 21344
rect 14553 21335 14611 21341
rect 14553 21332 14565 21335
rect 14148 21304 14565 21332
rect 14148 21292 14154 21304
rect 14553 21301 14565 21304
rect 14599 21301 14611 21335
rect 14553 21295 14611 21301
rect 14734 21292 14740 21344
rect 14792 21332 14798 21344
rect 15381 21335 15439 21341
rect 15381 21332 15393 21335
rect 14792 21304 15393 21332
rect 14792 21292 14798 21304
rect 15381 21301 15393 21304
rect 15427 21301 15439 21335
rect 15381 21295 15439 21301
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 15565 21335 15623 21341
rect 15565 21332 15577 21335
rect 15528 21304 15577 21332
rect 15528 21292 15534 21304
rect 15565 21301 15577 21304
rect 15611 21301 15623 21335
rect 16132 21332 16160 21508
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 17221 21539 17279 21545
rect 17221 21536 17233 21539
rect 16632 21508 17233 21536
rect 16632 21496 16638 21508
rect 17221 21505 17233 21508
rect 17267 21505 17279 21539
rect 17221 21499 17279 21505
rect 21453 21539 21511 21545
rect 21453 21505 21465 21539
rect 21499 21536 21511 21539
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 21499 21508 22385 21536
rect 21499 21505 21511 21508
rect 21453 21499 21511 21505
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 22462 21496 22468 21548
rect 22520 21496 22526 21548
rect 23198 21536 23204 21548
rect 22572 21508 23204 21536
rect 16209 21471 16267 21477
rect 16209 21437 16221 21471
rect 16255 21437 16267 21471
rect 16209 21431 16267 21437
rect 16224 21400 16252 21431
rect 17034 21428 17040 21480
rect 17092 21468 17098 21480
rect 17681 21471 17739 21477
rect 17681 21468 17693 21471
rect 17092 21440 17693 21468
rect 17092 21428 17098 21440
rect 17681 21437 17693 21440
rect 17727 21437 17739 21471
rect 17681 21431 17739 21437
rect 18690 21428 18696 21480
rect 18748 21428 18754 21480
rect 18969 21471 19027 21477
rect 18969 21468 18981 21471
rect 18800 21440 18981 21468
rect 17218 21400 17224 21412
rect 16224 21372 17224 21400
rect 17218 21360 17224 21372
rect 17276 21360 17282 21412
rect 18322 21360 18328 21412
rect 18380 21400 18386 21412
rect 18800 21400 18828 21440
rect 18969 21437 18981 21440
rect 19015 21437 19027 21471
rect 18969 21431 19027 21437
rect 19058 21428 19064 21480
rect 19116 21468 19122 21480
rect 22572 21468 22600 21508
rect 23198 21496 23204 21508
rect 23256 21496 23262 21548
rect 23382 21496 23388 21548
rect 23440 21496 23446 21548
rect 26068 21545 26096 21576
rect 28994 21564 29000 21576
rect 29052 21564 29058 21616
rect 29730 21564 29736 21616
rect 29788 21564 29794 21616
rect 26053 21539 26111 21545
rect 26053 21505 26065 21539
rect 26099 21505 26111 21539
rect 27617 21539 27675 21545
rect 26053 21499 26111 21505
rect 26160 21508 27568 21536
rect 19116 21440 22600 21468
rect 22649 21471 22707 21477
rect 19116 21428 19122 21440
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 24670 21468 24676 21480
rect 22695 21440 24676 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 24670 21428 24676 21440
rect 24728 21468 24734 21480
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24728 21440 25145 21468
rect 24728 21428 24734 21440
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 25958 21428 25964 21480
rect 26016 21468 26022 21480
rect 26160 21468 26188 21508
rect 26016 21440 26188 21468
rect 26237 21471 26295 21477
rect 26016 21428 26022 21440
rect 26237 21437 26249 21471
rect 26283 21437 26295 21471
rect 27540 21468 27568 21508
rect 27617 21505 27629 21539
rect 27663 21536 27675 21539
rect 27890 21536 27896 21548
rect 27663 21508 27896 21536
rect 27663 21505 27675 21508
rect 27617 21499 27675 21505
rect 27890 21496 27896 21508
rect 27948 21496 27954 21548
rect 27706 21468 27712 21480
rect 27540 21440 27712 21468
rect 26237 21431 26295 21437
rect 18380 21372 18828 21400
rect 20441 21403 20499 21409
rect 18380 21360 18386 21372
rect 20441 21369 20453 21403
rect 20487 21400 20499 21403
rect 20530 21400 20536 21412
rect 20487 21372 20536 21400
rect 20487 21369 20499 21372
rect 20441 21363 20499 21369
rect 20530 21360 20536 21372
rect 20588 21360 20594 21412
rect 20898 21360 20904 21412
rect 20956 21400 20962 21412
rect 22005 21403 22063 21409
rect 22005 21400 22017 21403
rect 20956 21372 22017 21400
rect 20956 21360 20962 21372
rect 22005 21369 22017 21372
rect 22051 21369 22063 21403
rect 22005 21363 22063 21369
rect 25590 21360 25596 21412
rect 25648 21360 25654 21412
rect 26252 21400 26280 21431
rect 27706 21428 27712 21440
rect 27764 21428 27770 21480
rect 27798 21428 27804 21480
rect 27856 21428 27862 21480
rect 28350 21428 28356 21480
rect 28408 21468 28414 21480
rect 28445 21471 28503 21477
rect 28445 21468 28457 21471
rect 28408 21440 28457 21468
rect 28408 21428 28414 21440
rect 28445 21437 28457 21440
rect 28491 21437 28503 21471
rect 28721 21471 28779 21477
rect 28721 21468 28733 21471
rect 28445 21431 28503 21437
rect 28552 21440 28733 21468
rect 28552 21400 28580 21440
rect 28721 21437 28733 21440
rect 28767 21468 28779 21471
rect 29086 21468 29092 21480
rect 28767 21440 29092 21468
rect 28767 21437 28779 21440
rect 28721 21431 28779 21437
rect 29086 21428 29092 21440
rect 29144 21428 29150 21480
rect 30944 21468 30972 21644
rect 32030 21632 32036 21684
rect 32088 21672 32094 21684
rect 32493 21675 32551 21681
rect 32493 21672 32505 21675
rect 32088 21644 32505 21672
rect 32088 21632 32094 21644
rect 32493 21641 32505 21644
rect 32539 21641 32551 21675
rect 32493 21635 32551 21641
rect 33045 21675 33103 21681
rect 33045 21641 33057 21675
rect 33091 21672 33103 21675
rect 34146 21672 34152 21684
rect 33091 21644 34152 21672
rect 33091 21641 33103 21644
rect 33045 21635 33103 21641
rect 34146 21632 34152 21644
rect 34204 21632 34210 21684
rect 31113 21607 31171 21613
rect 31113 21573 31125 21607
rect 31159 21604 31171 21607
rect 35250 21604 35256 21616
rect 31159 21576 35256 21604
rect 31159 21573 31171 21576
rect 31113 21567 31171 21573
rect 35250 21564 35256 21576
rect 35308 21564 35314 21616
rect 31018 21496 31024 21548
rect 31076 21496 31082 21548
rect 31754 21536 31760 21548
rect 31128 21508 31760 21536
rect 31128 21468 31156 21508
rect 31754 21496 31760 21508
rect 31812 21496 31818 21548
rect 32214 21496 32220 21548
rect 32272 21536 32278 21548
rect 32401 21539 32459 21545
rect 32401 21536 32413 21539
rect 32272 21508 32413 21536
rect 32272 21496 32278 21508
rect 32401 21505 32413 21508
rect 32447 21505 32459 21539
rect 32401 21499 32459 21505
rect 33229 21539 33287 21545
rect 33229 21505 33241 21539
rect 33275 21536 33287 21539
rect 33410 21536 33416 21548
rect 33275 21508 33416 21536
rect 33275 21505 33287 21508
rect 33229 21499 33287 21505
rect 33410 21496 33416 21508
rect 33468 21496 33474 21548
rect 47854 21496 47860 21548
rect 47912 21536 47918 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 47912 21508 47961 21536
rect 47912 21496 47918 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 30944 21440 31156 21468
rect 31205 21471 31263 21477
rect 31205 21437 31217 21471
rect 31251 21437 31263 21471
rect 31205 21431 31263 21437
rect 31220 21400 31248 21431
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 26252 21372 28580 21400
rect 30208 21372 31248 21400
rect 30208 21344 30236 21372
rect 17037 21335 17095 21341
rect 17037 21332 17049 21335
rect 16132 21304 17049 21332
rect 15565 21295 15623 21301
rect 17037 21301 17049 21304
rect 17083 21301 17095 21335
rect 17037 21295 17095 21301
rect 17494 21292 17500 21344
rect 17552 21332 17558 21344
rect 21450 21332 21456 21344
rect 17552 21304 21456 21332
rect 17552 21292 17558 21304
rect 21450 21292 21456 21304
rect 21508 21292 21514 21344
rect 22462 21292 22468 21344
rect 22520 21332 22526 21344
rect 25314 21332 25320 21344
rect 22520 21304 25320 21332
rect 22520 21292 22526 21304
rect 25314 21292 25320 21304
rect 25372 21292 25378 21344
rect 27246 21292 27252 21344
rect 27304 21292 27310 21344
rect 30190 21292 30196 21344
rect 30248 21292 30254 21344
rect 30650 21292 30656 21344
rect 30708 21292 30714 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 5994 21088 6000 21140
rect 6052 21128 6058 21140
rect 11425 21131 11483 21137
rect 11425 21128 11437 21131
rect 6052 21100 11437 21128
rect 6052 21088 6058 21100
rect 11425 21097 11437 21100
rect 11471 21097 11483 21131
rect 11425 21091 11483 21097
rect 12250 21088 12256 21140
rect 12308 21128 12314 21140
rect 12802 21128 12808 21140
rect 12308 21100 12808 21128
rect 12308 21088 12314 21100
rect 12802 21088 12808 21100
rect 12860 21088 12866 21140
rect 14369 21131 14427 21137
rect 14369 21097 14381 21131
rect 14415 21128 14427 21131
rect 17862 21128 17868 21140
rect 14415 21100 17868 21128
rect 14415 21097 14427 21100
rect 14369 21091 14427 21097
rect 17862 21088 17868 21100
rect 17920 21088 17926 21140
rect 19518 21088 19524 21140
rect 19576 21088 19582 21140
rect 19692 21131 19750 21137
rect 19692 21097 19704 21131
rect 19738 21128 19750 21131
rect 20438 21128 20444 21140
rect 19738 21100 20444 21128
rect 19738 21097 19750 21100
rect 19692 21091 19750 21097
rect 20438 21088 20444 21100
rect 20496 21088 20502 21140
rect 20714 21088 20720 21140
rect 20772 21128 20778 21140
rect 21177 21131 21235 21137
rect 21177 21128 21189 21131
rect 20772 21100 21189 21128
rect 20772 21088 20778 21100
rect 21177 21097 21189 21100
rect 21223 21097 21235 21131
rect 21177 21091 21235 21097
rect 21910 21088 21916 21140
rect 21968 21128 21974 21140
rect 24673 21131 24731 21137
rect 24673 21128 24685 21131
rect 21968 21100 24685 21128
rect 21968 21088 21974 21100
rect 24673 21097 24685 21100
rect 24719 21097 24731 21131
rect 30650 21128 30656 21140
rect 24673 21091 24731 21097
rect 25240 21100 30656 21128
rect 4982 21020 4988 21072
rect 5040 21060 5046 21072
rect 5353 21063 5411 21069
rect 5353 21060 5365 21063
rect 5040 21032 5365 21060
rect 5040 21020 5046 21032
rect 5353 21029 5365 21032
rect 5399 21029 5411 21063
rect 5353 21023 5411 21029
rect 6822 21020 6828 21072
rect 6880 21060 6886 21072
rect 7653 21063 7711 21069
rect 7653 21060 7665 21063
rect 6880 21032 7665 21060
rect 6880 21020 6886 21032
rect 7653 21029 7665 21032
rect 7699 21029 7711 21063
rect 7653 21023 7711 21029
rect 12342 21020 12348 21072
rect 12400 21060 12406 21072
rect 19536 21060 19564 21088
rect 12400 21032 15700 21060
rect 12400 21020 12406 21032
rect 4709 20995 4767 21001
rect 4709 20961 4721 20995
rect 4755 20992 4767 20995
rect 5166 20992 5172 21004
rect 4755 20964 5172 20992
rect 4755 20961 4767 20964
rect 4709 20955 4767 20961
rect 5166 20952 5172 20964
rect 5224 20952 5230 21004
rect 5813 20995 5871 21001
rect 5813 20961 5825 20995
rect 5859 20992 5871 20995
rect 8205 20995 8263 21001
rect 8205 20992 8217 20995
rect 5859 20964 8217 20992
rect 5859 20961 5871 20964
rect 5813 20955 5871 20961
rect 8205 20961 8217 20964
rect 8251 20961 8263 20995
rect 8205 20955 8263 20961
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 4338 20924 4344 20936
rect 1811 20896 4344 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 4338 20884 4344 20896
rect 4396 20884 4402 20936
rect 4798 20884 4804 20936
rect 4856 20924 4862 20936
rect 5537 20927 5595 20933
rect 5537 20924 5549 20927
rect 4856 20896 5549 20924
rect 4856 20884 4862 20896
rect 5537 20893 5549 20896
rect 5583 20893 5595 20927
rect 7558 20924 7564 20936
rect 5537 20887 5595 20893
rect 7116 20896 7564 20924
rect 2777 20859 2835 20865
rect 2777 20825 2789 20859
rect 2823 20856 2835 20859
rect 2866 20856 2872 20868
rect 2823 20828 2872 20856
rect 2823 20825 2835 20828
rect 2777 20819 2835 20825
rect 2866 20816 2872 20828
rect 2924 20816 2930 20868
rect 4525 20859 4583 20865
rect 4525 20825 4537 20859
rect 4571 20856 4583 20859
rect 4982 20856 4988 20868
rect 4571 20828 4988 20856
rect 4571 20825 4583 20828
rect 4525 20819 4583 20825
rect 4982 20816 4988 20828
rect 5040 20816 5046 20868
rect 5092 20828 6224 20856
rect 4154 20748 4160 20800
rect 4212 20748 4218 20800
rect 4617 20791 4675 20797
rect 4617 20757 4629 20791
rect 4663 20788 4675 20791
rect 5092 20788 5120 20828
rect 4663 20760 5120 20788
rect 6196 20788 6224 20828
rect 6270 20816 6276 20868
rect 6328 20816 6334 20868
rect 7116 20788 7144 20896
rect 7558 20884 7564 20896
rect 7616 20884 7622 20936
rect 8220 20924 8248 20955
rect 8386 20952 8392 21004
rect 8444 20992 8450 21004
rect 9585 20995 9643 21001
rect 9585 20992 9597 20995
rect 8444 20964 9597 20992
rect 8444 20952 8450 20964
rect 9585 20961 9597 20964
rect 9631 20961 9643 20995
rect 9585 20955 9643 20961
rect 12618 20952 12624 21004
rect 12676 20952 12682 21004
rect 14826 20952 14832 21004
rect 14884 20952 14890 21004
rect 15672 21001 15700 21032
rect 17604 21032 19564 21060
rect 15013 20995 15071 21001
rect 15013 20961 15025 20995
rect 15059 20961 15071 20995
rect 15013 20955 15071 20961
rect 15657 20995 15715 21001
rect 15657 20961 15669 20995
rect 15703 20961 15715 20995
rect 15657 20955 15715 20961
rect 15841 20995 15899 21001
rect 15841 20961 15853 20995
rect 15887 20992 15899 20995
rect 16666 20992 16672 21004
rect 15887 20964 16672 20992
rect 15887 20961 15899 20964
rect 15841 20955 15899 20961
rect 8754 20924 8760 20936
rect 8220 20896 8760 20924
rect 8754 20884 8760 20896
rect 8812 20884 8818 20936
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20924 9367 20927
rect 9398 20924 9404 20936
rect 9355 20896 9404 20924
rect 9355 20893 9367 20896
rect 9309 20887 9367 20893
rect 9398 20884 9404 20896
rect 9456 20884 9462 20936
rect 12161 20927 12219 20933
rect 12161 20893 12173 20927
rect 12207 20924 12219 20927
rect 12710 20924 12716 20936
rect 12207 20896 12716 20924
rect 12207 20893 12219 20896
rect 12161 20887 12219 20893
rect 12710 20884 12716 20896
rect 12768 20884 12774 20936
rect 15028 20924 15056 20955
rect 16666 20952 16672 20964
rect 16724 20952 16730 21004
rect 17604 21001 17632 21032
rect 20806 21020 20812 21072
rect 20864 21060 20870 21072
rect 23293 21063 23351 21069
rect 23293 21060 23305 21063
rect 20864 21032 23305 21060
rect 20864 21020 20870 21032
rect 23293 21029 23305 21032
rect 23339 21029 23351 21063
rect 25240 21060 25268 21100
rect 30650 21088 30656 21100
rect 30708 21088 30714 21140
rect 31846 21088 31852 21140
rect 31904 21128 31910 21140
rect 32493 21131 32551 21137
rect 32493 21128 32505 21131
rect 31904 21100 32505 21128
rect 31904 21088 31910 21100
rect 32493 21097 32505 21100
rect 32539 21097 32551 21131
rect 32493 21091 32551 21097
rect 25958 21060 25964 21072
rect 23293 21023 23351 21029
rect 25148 21032 25268 21060
rect 25332 21032 25964 21060
rect 17589 20995 17647 21001
rect 16776 20964 17540 20992
rect 16776 20924 16804 20964
rect 15028 20896 16804 20924
rect 17034 20884 17040 20936
rect 17092 20924 17098 20936
rect 17313 20927 17371 20933
rect 17313 20924 17325 20927
rect 17092 20896 17325 20924
rect 17092 20884 17098 20896
rect 17313 20893 17325 20896
rect 17359 20924 17371 20927
rect 17402 20924 17408 20936
rect 17359 20896 17408 20924
rect 17359 20893 17371 20896
rect 17313 20887 17371 20893
rect 17402 20884 17408 20896
rect 17460 20884 17466 20936
rect 7466 20816 7472 20868
rect 7524 20856 7530 20868
rect 8113 20859 8171 20865
rect 8113 20856 8125 20859
rect 7524 20828 8125 20856
rect 7524 20816 7530 20828
rect 8113 20825 8125 20828
rect 8159 20825 8171 20859
rect 8113 20819 8171 20825
rect 11330 20816 11336 20868
rect 11388 20816 11394 20868
rect 15470 20856 15476 20868
rect 12406 20828 15476 20856
rect 6196 20760 7144 20788
rect 4663 20757 4675 20760
rect 4617 20751 4675 20757
rect 7190 20748 7196 20800
rect 7248 20788 7254 20800
rect 7285 20791 7343 20797
rect 7285 20788 7297 20791
rect 7248 20760 7297 20788
rect 7248 20748 7254 20760
rect 7285 20757 7297 20760
rect 7331 20757 7343 20791
rect 7285 20751 7343 20757
rect 7374 20748 7380 20800
rect 7432 20788 7438 20800
rect 8021 20791 8079 20797
rect 8021 20788 8033 20791
rect 7432 20760 8033 20788
rect 7432 20748 7438 20760
rect 8021 20757 8033 20760
rect 8067 20757 8079 20791
rect 8021 20751 8079 20757
rect 11146 20748 11152 20800
rect 11204 20788 11210 20800
rect 12406 20788 12434 20828
rect 15470 20816 15476 20828
rect 15528 20816 15534 20868
rect 16850 20856 16856 20868
rect 15580 20828 16856 20856
rect 11204 20760 12434 20788
rect 11204 20748 11210 20760
rect 13998 20748 14004 20800
rect 14056 20788 14062 20800
rect 14734 20788 14740 20800
rect 14056 20760 14740 20788
rect 14056 20748 14062 20760
rect 14734 20748 14740 20760
rect 14792 20748 14798 20800
rect 15194 20748 15200 20800
rect 15252 20748 15258 20800
rect 15580 20797 15608 20828
rect 16850 20816 16856 20828
rect 16908 20816 16914 20868
rect 17126 20856 17132 20868
rect 16960 20828 17132 20856
rect 15565 20791 15623 20797
rect 15565 20757 15577 20791
rect 15611 20757 15623 20791
rect 15565 20751 15623 20757
rect 16390 20748 16396 20800
rect 16448 20748 16454 20800
rect 16960 20797 16988 20828
rect 17126 20816 17132 20828
rect 17184 20816 17190 20868
rect 17512 20856 17540 20964
rect 17589 20961 17601 20995
rect 17635 20961 17647 20995
rect 17589 20955 17647 20961
rect 18598 20952 18604 21004
rect 18656 20952 18662 21004
rect 18785 20995 18843 21001
rect 18785 20961 18797 20995
rect 18831 20992 18843 20995
rect 19058 20992 19064 21004
rect 18831 20964 19064 20992
rect 18831 20961 18843 20964
rect 18785 20955 18843 20961
rect 19058 20952 19064 20964
rect 19116 20952 19122 21004
rect 19429 20995 19487 21001
rect 19429 20961 19441 20995
rect 19475 20992 19487 20995
rect 19702 20992 19708 21004
rect 19475 20964 19708 20992
rect 19475 20961 19487 20964
rect 19429 20955 19487 20961
rect 19702 20952 19708 20964
rect 19760 20992 19766 21004
rect 20346 20992 20352 21004
rect 19760 20964 20352 20992
rect 19760 20952 19766 20964
rect 20346 20952 20352 20964
rect 20404 20992 20410 21004
rect 21174 20992 21180 21004
rect 20404 20964 21180 20992
rect 20404 20952 20410 20964
rect 21174 20952 21180 20964
rect 21232 20992 21238 21004
rect 22097 20995 22155 21001
rect 22097 20992 22109 20995
rect 21232 20964 22109 20992
rect 21232 20952 21238 20964
rect 22097 20961 22109 20964
rect 22143 20961 22155 20995
rect 22097 20955 22155 20961
rect 23198 20952 23204 21004
rect 23256 20992 23262 21004
rect 23658 20992 23664 21004
rect 23256 20964 23664 20992
rect 23256 20952 23262 20964
rect 23658 20952 23664 20964
rect 23716 20952 23722 21004
rect 23842 20952 23848 21004
rect 23900 20952 23906 21004
rect 25148 21001 25176 21032
rect 25332 21001 25360 21032
rect 25958 21020 25964 21032
rect 26016 21020 26022 21072
rect 27522 21020 27528 21072
rect 27580 21060 27586 21072
rect 27580 21032 30052 21060
rect 27580 21020 27586 21032
rect 25133 20995 25191 21001
rect 25133 20961 25145 20995
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 25317 20995 25375 21001
rect 25317 20961 25329 20995
rect 25363 20961 25375 20995
rect 25317 20955 25375 20961
rect 25774 20952 25780 21004
rect 25832 20992 25838 21004
rect 26050 20992 26056 21004
rect 25832 20964 26056 20992
rect 25832 20952 25838 20964
rect 26050 20952 26056 20964
rect 26108 20992 26114 21004
rect 28350 20992 28356 21004
rect 26108 20964 28356 20992
rect 26108 20952 26114 20964
rect 28350 20952 28356 20964
rect 28408 20952 28414 21004
rect 30024 21001 30052 21032
rect 30009 20995 30067 21001
rect 30009 20961 30021 20995
rect 30055 20961 30067 20995
rect 30009 20955 30067 20961
rect 21082 20924 21088 20936
rect 20838 20896 21088 20924
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 21542 20884 21548 20936
rect 21600 20924 21606 20936
rect 22741 20927 22799 20933
rect 22741 20924 22753 20927
rect 21600 20896 22753 20924
rect 21600 20884 21606 20896
rect 22741 20893 22753 20896
rect 22787 20893 22799 20927
rect 22741 20887 22799 20893
rect 19978 20856 19984 20868
rect 17512 20828 19984 20856
rect 19978 20816 19984 20828
rect 20036 20816 20042 20868
rect 21361 20859 21419 20865
rect 21361 20856 21373 20859
rect 21008 20828 21373 20856
rect 16945 20791 17003 20797
rect 16945 20757 16957 20791
rect 16991 20757 17003 20791
rect 16945 20751 17003 20757
rect 17402 20748 17408 20800
rect 17460 20748 17466 20800
rect 18141 20791 18199 20797
rect 18141 20757 18153 20791
rect 18187 20788 18199 20791
rect 18414 20788 18420 20800
rect 18187 20760 18420 20788
rect 18187 20757 18199 20760
rect 18141 20751 18199 20757
rect 18414 20748 18420 20760
rect 18472 20748 18478 20800
rect 18509 20791 18567 20797
rect 18509 20757 18521 20791
rect 18555 20788 18567 20791
rect 19242 20788 19248 20800
rect 18555 20760 19248 20788
rect 18555 20757 18567 20760
rect 18509 20751 18567 20757
rect 19242 20748 19248 20760
rect 19300 20748 19306 20800
rect 19334 20748 19340 20800
rect 19392 20788 19398 20800
rect 20622 20788 20628 20800
rect 19392 20760 20628 20788
rect 19392 20748 19398 20760
rect 20622 20748 20628 20760
rect 20680 20748 20686 20800
rect 20714 20748 20720 20800
rect 20772 20788 20778 20800
rect 21008 20788 21036 20828
rect 21361 20825 21373 20828
rect 21407 20825 21419 20859
rect 22756 20856 22784 20887
rect 23474 20884 23480 20936
rect 23532 20924 23538 20936
rect 24946 20924 24952 20936
rect 23532 20896 24952 20924
rect 23532 20884 23538 20896
rect 24946 20884 24952 20896
rect 25004 20884 25010 20936
rect 27706 20884 27712 20936
rect 27764 20884 27770 20936
rect 28261 20927 28319 20933
rect 28261 20893 28273 20927
rect 28307 20924 28319 20927
rect 28442 20924 28448 20936
rect 28307 20896 28448 20924
rect 28307 20893 28319 20896
rect 28261 20887 28319 20893
rect 28442 20884 28448 20896
rect 28500 20884 28506 20936
rect 28534 20884 28540 20936
rect 28592 20884 28598 20936
rect 29362 20884 29368 20936
rect 29420 20924 29426 20936
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 29420 20896 29745 20924
rect 29420 20884 29426 20896
rect 29733 20893 29745 20896
rect 29779 20893 29791 20927
rect 29733 20887 29791 20893
rect 29822 20884 29828 20936
rect 29880 20924 29886 20936
rect 31021 20927 31079 20933
rect 31021 20924 31033 20927
rect 29880 20896 31033 20924
rect 29880 20884 29886 20896
rect 31021 20893 31033 20896
rect 31067 20893 31079 20927
rect 31021 20887 31079 20893
rect 31294 20884 31300 20936
rect 31352 20884 31358 20936
rect 23753 20859 23811 20865
rect 23753 20856 23765 20859
rect 22756 20828 23765 20856
rect 21361 20819 21419 20825
rect 23753 20825 23765 20828
rect 23799 20825 23811 20859
rect 23753 20819 23811 20825
rect 25041 20859 25099 20865
rect 25041 20825 25053 20859
rect 25087 20856 25099 20859
rect 26234 20856 26240 20868
rect 25087 20828 26240 20856
rect 25087 20825 25099 20828
rect 25041 20819 25099 20825
rect 26234 20816 26240 20828
rect 26292 20816 26298 20868
rect 26329 20859 26387 20865
rect 26329 20825 26341 20859
rect 26375 20825 26387 20859
rect 26329 20819 26387 20825
rect 20772 20760 21036 20788
rect 20772 20748 20778 20760
rect 23658 20748 23664 20800
rect 23716 20748 23722 20800
rect 26344 20788 26372 20819
rect 27062 20816 27068 20868
rect 27120 20816 27126 20868
rect 27724 20856 27752 20884
rect 27724 20828 27844 20856
rect 27706 20788 27712 20800
rect 26344 20760 27712 20788
rect 27706 20748 27712 20760
rect 27764 20748 27770 20800
rect 27816 20797 27844 20828
rect 32306 20816 32312 20868
rect 32364 20856 32370 20868
rect 32401 20859 32459 20865
rect 32401 20856 32413 20859
rect 32364 20828 32413 20856
rect 32364 20816 32370 20828
rect 32401 20825 32413 20828
rect 32447 20825 32459 20859
rect 32401 20819 32459 20825
rect 27801 20791 27859 20797
rect 27801 20757 27813 20791
rect 27847 20757 27859 20791
rect 27801 20751 27859 20757
rect 27890 20748 27896 20800
rect 27948 20788 27954 20800
rect 28534 20788 28540 20800
rect 27948 20760 28540 20788
rect 27948 20748 27954 20760
rect 28534 20748 28540 20760
rect 28592 20788 28598 20800
rect 31018 20788 31024 20800
rect 28592 20760 31024 20788
rect 28592 20748 28598 20760
rect 31018 20748 31024 20760
rect 31076 20748 31082 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 5629 20587 5687 20593
rect 5629 20553 5641 20587
rect 5675 20584 5687 20587
rect 6086 20584 6092 20596
rect 5675 20556 6092 20584
rect 5675 20553 5687 20556
rect 5629 20547 5687 20553
rect 6086 20544 6092 20556
rect 6144 20584 6150 20596
rect 10410 20584 10416 20596
rect 6144 20556 10416 20584
rect 6144 20544 6150 20556
rect 10410 20544 10416 20556
rect 10468 20544 10474 20596
rect 11882 20544 11888 20596
rect 11940 20544 11946 20596
rect 12989 20587 13047 20593
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 17218 20584 17224 20596
rect 13035 20556 17224 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 17310 20544 17316 20596
rect 17368 20544 17374 20596
rect 17405 20587 17463 20593
rect 17405 20553 17417 20587
rect 17451 20584 17463 20587
rect 17451 20556 21312 20584
rect 17451 20553 17463 20556
rect 17405 20547 17463 20553
rect 6914 20516 6920 20528
rect 3620 20488 6920 20516
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20448 1823 20451
rect 1854 20448 1860 20460
rect 1811 20420 1860 20448
rect 1811 20417 1823 20420
rect 1765 20411 1823 20417
rect 1854 20408 1860 20420
rect 1912 20408 1918 20460
rect 3620 20457 3648 20488
rect 6914 20476 6920 20488
rect 6972 20476 6978 20528
rect 10226 20476 10232 20528
rect 10284 20516 10290 20528
rect 12897 20519 12955 20525
rect 12897 20516 12909 20519
rect 10284 20488 12909 20516
rect 10284 20476 10290 20488
rect 12897 20485 12909 20488
rect 12943 20485 12955 20519
rect 12897 20479 12955 20485
rect 13354 20476 13360 20528
rect 13412 20516 13418 20528
rect 14274 20516 14280 20528
rect 13412 20488 14280 20516
rect 13412 20476 13418 20488
rect 14274 20476 14280 20488
rect 14332 20516 14338 20528
rect 18601 20519 18659 20525
rect 14332 20488 14490 20516
rect 14332 20476 14338 20488
rect 18601 20485 18613 20519
rect 18647 20516 18659 20519
rect 18966 20516 18972 20528
rect 18647 20488 18972 20516
rect 18647 20485 18659 20488
rect 18601 20479 18659 20485
rect 18966 20476 18972 20488
rect 19024 20476 19030 20528
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20417 3663 20451
rect 3605 20411 3663 20417
rect 6546 20408 6552 20460
rect 6604 20408 6610 20460
rect 8386 20408 8392 20460
rect 8444 20408 8450 20460
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 10502 20448 10508 20460
rect 9732 20420 10508 20448
rect 9732 20408 9738 20420
rect 10502 20408 10508 20420
rect 10560 20408 10566 20460
rect 10689 20451 10747 20457
rect 10689 20417 10701 20451
rect 10735 20448 10747 20451
rect 11054 20448 11060 20460
rect 10735 20420 11060 20448
rect 10735 20417 10747 20420
rect 10689 20411 10747 20417
rect 11054 20408 11060 20420
rect 11112 20408 11118 20460
rect 11606 20408 11612 20460
rect 11664 20448 11670 20460
rect 11793 20451 11851 20457
rect 11793 20448 11805 20451
rect 11664 20420 11805 20448
rect 11664 20408 11670 20420
rect 11793 20417 11805 20420
rect 11839 20448 11851 20451
rect 12250 20448 12256 20460
rect 11839 20420 12256 20448
rect 11839 20417 11851 20420
rect 11793 20411 11851 20417
rect 12250 20408 12256 20420
rect 12308 20408 12314 20460
rect 15286 20408 15292 20460
rect 15344 20448 15350 20460
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15344 20420 16037 20448
rect 15344 20408 15350 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 16390 20408 16396 20460
rect 16448 20448 16454 20460
rect 17402 20448 17408 20460
rect 16448 20420 17408 20448
rect 16448 20408 16454 20420
rect 17402 20408 17408 20420
rect 17460 20408 17466 20460
rect 18414 20448 18420 20460
rect 17512 20420 18420 20448
rect 2774 20340 2780 20392
rect 2832 20340 2838 20392
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 5718 20340 5724 20392
rect 5776 20340 5782 20392
rect 5810 20340 5816 20392
rect 5868 20340 5874 20392
rect 5902 20340 5908 20392
rect 5960 20380 5966 20392
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 5960 20352 7021 20380
rect 5960 20340 5966 20352
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 7009 20343 7067 20349
rect 7098 20340 7104 20392
rect 7156 20380 7162 20392
rect 7466 20380 7472 20392
rect 7156 20352 7472 20380
rect 7156 20340 7162 20352
rect 7466 20340 7472 20352
rect 7524 20340 7530 20392
rect 8665 20383 8723 20389
rect 8665 20349 8677 20383
rect 8711 20380 8723 20383
rect 11698 20380 11704 20392
rect 8711 20352 11704 20380
rect 8711 20349 8723 20352
rect 8665 20343 8723 20349
rect 11698 20340 11704 20352
rect 11756 20340 11762 20392
rect 13173 20383 13231 20389
rect 13173 20349 13185 20383
rect 13219 20380 13231 20383
rect 13446 20380 13452 20392
rect 13219 20352 13452 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 13446 20340 13452 20352
rect 13504 20340 13510 20392
rect 13722 20340 13728 20392
rect 13780 20340 13786 20392
rect 14001 20383 14059 20389
rect 14001 20349 14013 20383
rect 14047 20380 14059 20383
rect 14090 20380 14096 20392
rect 14047 20352 14096 20380
rect 14047 20349 14059 20352
rect 14001 20343 14059 20349
rect 14090 20340 14096 20352
rect 14148 20380 14154 20392
rect 17512 20380 17540 20420
rect 18414 20408 18420 20420
rect 18472 20408 18478 20460
rect 18506 20408 18512 20460
rect 18564 20408 18570 20460
rect 19702 20408 19708 20460
rect 19760 20408 19766 20460
rect 21082 20408 21088 20460
rect 21140 20408 21146 20460
rect 14148 20352 17540 20380
rect 17589 20383 17647 20389
rect 14148 20340 14154 20352
rect 17589 20349 17601 20383
rect 17635 20349 17647 20383
rect 17589 20343 17647 20349
rect 18785 20383 18843 20389
rect 18785 20349 18797 20383
rect 18831 20380 18843 20383
rect 18874 20380 18880 20392
rect 18831 20352 18880 20380
rect 18831 20349 18843 20352
rect 18785 20343 18843 20349
rect 5261 20315 5319 20321
rect 5261 20281 5273 20315
rect 5307 20312 5319 20315
rect 7190 20312 7196 20324
rect 5307 20284 7196 20312
rect 5307 20281 5319 20284
rect 5261 20275 5319 20281
rect 7190 20272 7196 20284
rect 7248 20272 7254 20324
rect 10873 20315 10931 20321
rect 10873 20312 10885 20315
rect 9692 20284 10885 20312
rect 5626 20204 5632 20256
rect 5684 20244 5690 20256
rect 9692 20244 9720 20284
rect 10873 20281 10885 20284
rect 10919 20281 10931 20315
rect 10873 20275 10931 20281
rect 12526 20272 12532 20324
rect 12584 20272 12590 20324
rect 15286 20272 15292 20324
rect 15344 20312 15350 20324
rect 15930 20312 15936 20324
rect 15344 20284 15936 20312
rect 15344 20272 15350 20284
rect 15930 20272 15936 20284
rect 15988 20272 15994 20324
rect 17604 20312 17632 20343
rect 18874 20340 18880 20352
rect 18932 20340 18938 20392
rect 19978 20340 19984 20392
rect 20036 20340 20042 20392
rect 21100 20312 21128 20408
rect 21284 20380 21312 20556
rect 21450 20544 21456 20596
rect 21508 20544 21514 20596
rect 22830 20544 22836 20596
rect 22888 20584 22894 20596
rect 23477 20587 23535 20593
rect 23477 20584 23489 20587
rect 22888 20556 23489 20584
rect 22888 20544 22894 20556
rect 23477 20553 23489 20556
rect 23523 20553 23535 20587
rect 23477 20547 23535 20553
rect 23569 20587 23627 20593
rect 23569 20553 23581 20587
rect 23615 20584 23627 20587
rect 27246 20584 27252 20596
rect 23615 20556 27252 20584
rect 23615 20553 23627 20556
rect 23569 20547 23627 20553
rect 27246 20544 27252 20556
rect 27304 20544 27310 20596
rect 27617 20587 27675 20593
rect 27617 20553 27629 20587
rect 27663 20584 27675 20587
rect 28902 20584 28908 20596
rect 27663 20556 28908 20584
rect 27663 20553 27675 20556
rect 27617 20547 27675 20553
rect 28902 20544 28908 20556
rect 28960 20544 28966 20596
rect 30101 20587 30159 20593
rect 30101 20584 30113 20587
rect 29012 20556 30113 20584
rect 22097 20519 22155 20525
rect 22097 20485 22109 20519
rect 22143 20516 22155 20519
rect 23382 20516 23388 20528
rect 22143 20488 23388 20516
rect 22143 20485 22155 20488
rect 22097 20479 22155 20485
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 24854 20516 24860 20528
rect 24320 20488 24860 20516
rect 24320 20457 24348 20488
rect 24854 20476 24860 20488
rect 24912 20476 24918 20528
rect 26418 20476 26424 20528
rect 26476 20516 26482 20528
rect 29012 20516 29040 20556
rect 30101 20553 30113 20556
rect 30147 20553 30159 20587
rect 30101 20547 30159 20553
rect 31021 20587 31079 20593
rect 31021 20553 31033 20587
rect 31067 20584 31079 20587
rect 34698 20584 34704 20596
rect 31067 20556 34704 20584
rect 31067 20553 31079 20556
rect 31021 20547 31079 20553
rect 34698 20544 34704 20556
rect 34756 20544 34762 20596
rect 26476 20488 29040 20516
rect 26476 20476 26482 20488
rect 29638 20476 29644 20528
rect 29696 20476 29702 20528
rect 30116 20488 31156 20516
rect 30116 20460 30144 20488
rect 24305 20451 24363 20457
rect 24305 20417 24317 20451
rect 24351 20417 24363 20451
rect 27062 20448 27068 20460
rect 25714 20434 27068 20448
rect 24305 20411 24363 20417
rect 25700 20420 27068 20434
rect 23566 20380 23572 20392
rect 21284 20352 23572 20380
rect 23566 20340 23572 20352
rect 23624 20340 23630 20392
rect 23753 20383 23811 20389
rect 23753 20349 23765 20383
rect 23799 20349 23811 20383
rect 23753 20343 23811 20349
rect 24581 20383 24639 20389
rect 24581 20349 24593 20383
rect 24627 20380 24639 20383
rect 24670 20380 24676 20392
rect 24627 20352 24676 20380
rect 24627 20349 24639 20352
rect 24581 20343 24639 20349
rect 21634 20312 21640 20324
rect 17604 20284 19748 20312
rect 21100 20284 21640 20312
rect 5684 20216 9720 20244
rect 5684 20204 5690 20216
rect 10042 20204 10048 20256
rect 10100 20244 10106 20256
rect 10137 20247 10195 20253
rect 10137 20244 10149 20247
rect 10100 20216 10149 20244
rect 10100 20204 10106 20216
rect 10137 20213 10149 20216
rect 10183 20213 10195 20247
rect 10137 20207 10195 20213
rect 10410 20204 10416 20256
rect 10468 20244 10474 20256
rect 14642 20244 14648 20256
rect 10468 20216 14648 20244
rect 10468 20204 10474 20216
rect 14642 20204 14648 20216
rect 14700 20244 14706 20256
rect 15102 20244 15108 20256
rect 14700 20216 15108 20244
rect 14700 20204 14706 20216
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 15470 20204 15476 20256
rect 15528 20204 15534 20256
rect 15562 20204 15568 20256
rect 15620 20244 15626 20256
rect 16117 20247 16175 20253
rect 16117 20244 16129 20247
rect 15620 20216 16129 20244
rect 15620 20204 15626 20216
rect 16117 20213 16129 20216
rect 16163 20213 16175 20247
rect 16117 20207 16175 20213
rect 16945 20247 17003 20253
rect 16945 20213 16957 20247
rect 16991 20244 17003 20247
rect 17310 20244 17316 20256
rect 16991 20216 17316 20244
rect 16991 20213 17003 20216
rect 16945 20207 17003 20213
rect 17310 20204 17316 20216
rect 17368 20204 17374 20256
rect 18141 20247 18199 20253
rect 18141 20213 18153 20247
rect 18187 20244 18199 20247
rect 19058 20244 19064 20256
rect 18187 20216 19064 20244
rect 18187 20213 18199 20216
rect 18141 20207 18199 20213
rect 19058 20204 19064 20216
rect 19116 20204 19122 20256
rect 19720 20244 19748 20284
rect 21634 20272 21640 20284
rect 21692 20272 21698 20324
rect 23109 20315 23167 20321
rect 23109 20312 23121 20315
rect 22066 20284 23121 20312
rect 20530 20244 20536 20256
rect 19720 20216 20536 20244
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 20714 20204 20720 20256
rect 20772 20244 20778 20256
rect 22066 20244 22094 20284
rect 23109 20281 23121 20284
rect 23155 20281 23167 20315
rect 23109 20275 23167 20281
rect 20772 20216 22094 20244
rect 20772 20204 20778 20216
rect 22186 20204 22192 20256
rect 22244 20204 22250 20256
rect 23768 20244 23796 20343
rect 24670 20340 24676 20352
rect 24728 20340 24734 20392
rect 25222 20340 25228 20392
rect 25280 20380 25286 20392
rect 25700 20380 25728 20420
rect 27062 20408 27068 20420
rect 27120 20408 27126 20460
rect 27154 20408 27160 20460
rect 27212 20448 27218 20460
rect 27522 20448 27528 20460
rect 27212 20420 27528 20448
rect 27212 20408 27218 20420
rect 27522 20408 27528 20420
rect 27580 20408 27586 20460
rect 28350 20408 28356 20460
rect 28408 20408 28414 20460
rect 30098 20408 30104 20460
rect 30156 20408 30162 20460
rect 30929 20451 30987 20457
rect 30929 20417 30941 20451
rect 30975 20417 30987 20451
rect 30929 20411 30987 20417
rect 25280 20352 25728 20380
rect 27709 20383 27767 20389
rect 25280 20340 25286 20352
rect 27709 20349 27721 20383
rect 27755 20349 27767 20383
rect 27709 20343 27767 20349
rect 28629 20383 28687 20389
rect 28629 20349 28641 20383
rect 28675 20380 28687 20383
rect 30190 20380 30196 20392
rect 28675 20352 30196 20380
rect 28675 20349 28687 20352
rect 28629 20343 28687 20349
rect 25682 20272 25688 20324
rect 25740 20312 25746 20324
rect 26053 20315 26111 20321
rect 26053 20312 26065 20315
rect 25740 20284 26065 20312
rect 25740 20272 25746 20284
rect 26053 20281 26065 20284
rect 26099 20312 26111 20315
rect 27724 20312 27752 20343
rect 30190 20340 30196 20352
rect 30248 20340 30254 20392
rect 30944 20312 30972 20411
rect 31128 20389 31156 20488
rect 31113 20383 31171 20389
rect 31113 20349 31125 20383
rect 31159 20349 31171 20383
rect 31113 20343 31171 20349
rect 26099 20284 27752 20312
rect 30208 20284 30972 20312
rect 26099 20281 26111 20284
rect 26053 20275 26111 20281
rect 25866 20244 25872 20256
rect 23768 20216 25872 20244
rect 25866 20204 25872 20216
rect 25924 20204 25930 20256
rect 27154 20204 27160 20256
rect 27212 20204 27218 20256
rect 27338 20204 27344 20256
rect 27396 20244 27402 20256
rect 30208 20244 30236 20284
rect 27396 20216 30236 20244
rect 27396 20204 27402 20216
rect 30282 20204 30288 20256
rect 30340 20244 30346 20256
rect 30561 20247 30619 20253
rect 30561 20244 30573 20247
rect 30340 20216 30573 20244
rect 30340 20204 30346 20216
rect 30561 20213 30573 20216
rect 30607 20213 30619 20247
rect 30561 20207 30619 20213
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 2498 20000 2504 20052
rect 2556 20040 2562 20052
rect 5902 20040 5908 20052
rect 2556 20012 5908 20040
rect 2556 20000 2562 20012
rect 5902 20000 5908 20012
rect 5960 20000 5966 20052
rect 6273 20043 6331 20049
rect 6273 20009 6285 20043
rect 6319 20040 6331 20043
rect 6730 20040 6736 20052
rect 6319 20012 6736 20040
rect 6319 20009 6331 20012
rect 6273 20003 6331 20009
rect 6730 20000 6736 20012
rect 6788 20000 6794 20052
rect 6996 20043 7054 20049
rect 6996 20009 7008 20043
rect 7042 20040 7054 20043
rect 10042 20040 10048 20052
rect 7042 20012 10048 20040
rect 7042 20009 7054 20012
rect 6996 20003 7054 20009
rect 10042 20000 10048 20012
rect 10100 20000 10106 20052
rect 11698 20000 11704 20052
rect 11756 20040 11762 20052
rect 12526 20040 12532 20052
rect 11756 20012 12532 20040
rect 11756 20000 11762 20012
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 16301 20043 16359 20049
rect 16301 20040 16313 20043
rect 15436 20012 16313 20040
rect 15436 20000 15442 20012
rect 16301 20009 16313 20012
rect 16347 20009 16359 20043
rect 16301 20003 16359 20009
rect 16945 20043 17003 20049
rect 16945 20009 16957 20043
rect 16991 20009 17003 20043
rect 16945 20003 17003 20009
rect 8386 19932 8392 19984
rect 8444 19972 8450 19984
rect 9214 19972 9220 19984
rect 8444 19944 9220 19972
rect 8444 19932 8450 19944
rect 9214 19932 9220 19944
rect 9272 19932 9278 19984
rect 12434 19972 12440 19984
rect 12406 19932 12440 19972
rect 12492 19972 12498 19984
rect 13722 19972 13728 19984
rect 12492 19944 13728 19972
rect 12492 19932 12498 19944
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 16960 19972 16988 20003
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 23293 20043 23351 20049
rect 23293 20040 23305 20043
rect 18932 20012 23305 20040
rect 18932 20000 18938 20012
rect 23293 20009 23305 20012
rect 23339 20009 23351 20043
rect 23293 20003 23351 20009
rect 23566 20000 23572 20052
rect 23624 20040 23630 20052
rect 27154 20040 27160 20052
rect 23624 20012 27160 20040
rect 23624 20000 23630 20012
rect 27154 20000 27160 20012
rect 27212 20000 27218 20052
rect 27617 20043 27675 20049
rect 27617 20009 27629 20043
rect 27663 20040 27675 20043
rect 27798 20040 27804 20052
rect 27663 20012 27804 20040
rect 27663 20009 27675 20012
rect 27617 20003 27675 20009
rect 27798 20000 27804 20012
rect 27856 20000 27862 20052
rect 19518 19972 19524 19984
rect 16960 19944 19524 19972
rect 19518 19932 19524 19944
rect 19576 19932 19582 19984
rect 21542 19932 21548 19984
rect 21600 19972 21606 19984
rect 22005 19975 22063 19981
rect 22005 19972 22017 19975
rect 21600 19944 22017 19972
rect 21600 19932 21606 19944
rect 22005 19941 22017 19944
rect 22051 19941 22063 19975
rect 22005 19935 22063 19941
rect 1394 19864 1400 19916
rect 1452 19904 1458 19916
rect 2041 19907 2099 19913
rect 2041 19904 2053 19907
rect 1452 19876 2053 19904
rect 1452 19864 1458 19876
rect 2041 19873 2053 19876
rect 2087 19873 2099 19907
rect 2041 19867 2099 19873
rect 4525 19907 4583 19913
rect 4525 19873 4537 19907
rect 4571 19904 4583 19907
rect 6733 19907 6791 19913
rect 6733 19904 6745 19907
rect 4571 19876 6745 19904
rect 4571 19873 4583 19876
rect 4525 19867 4583 19873
rect 6733 19873 6745 19876
rect 6779 19904 6791 19907
rect 7006 19904 7012 19916
rect 6779 19876 7012 19904
rect 6779 19873 6791 19876
rect 6733 19867 6791 19873
rect 7006 19864 7012 19876
rect 7064 19864 7070 19916
rect 7466 19864 7472 19916
rect 7524 19904 7530 19916
rect 8478 19904 8484 19916
rect 7524 19876 8484 19904
rect 7524 19864 7530 19876
rect 1762 19796 1768 19848
rect 1820 19796 1826 19848
rect 8128 19822 8156 19876
rect 8478 19864 8484 19876
rect 8536 19904 8542 19916
rect 9674 19904 9680 19916
rect 8536 19876 9680 19904
rect 8536 19864 8542 19876
rect 9674 19864 9680 19876
rect 9732 19864 9738 19916
rect 9953 19907 10011 19913
rect 9953 19873 9965 19907
rect 9999 19904 10011 19907
rect 12406 19904 12434 19932
rect 9999 19876 12434 19904
rect 13633 19907 13691 19913
rect 9999 19873 10011 19876
rect 9953 19867 10011 19873
rect 13633 19873 13645 19907
rect 13679 19904 13691 19907
rect 14829 19907 14887 19913
rect 14829 19904 14841 19907
rect 13679 19876 14841 19904
rect 13679 19873 13691 19876
rect 13633 19867 13691 19873
rect 14829 19873 14841 19876
rect 14875 19904 14887 19907
rect 15470 19904 15476 19916
rect 14875 19876 15476 19904
rect 14875 19873 14887 19876
rect 14829 19867 14887 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 17126 19864 17132 19916
rect 17184 19904 17190 19916
rect 17405 19907 17463 19913
rect 17405 19904 17417 19907
rect 17184 19876 17417 19904
rect 17184 19864 17190 19876
rect 17405 19873 17417 19876
rect 17451 19873 17463 19907
rect 17405 19867 17463 19873
rect 17589 19907 17647 19913
rect 17589 19873 17601 19907
rect 17635 19904 17647 19907
rect 18230 19904 18236 19916
rect 17635 19876 18236 19904
rect 17635 19873 17647 19876
rect 17589 19867 17647 19873
rect 18230 19864 18236 19876
rect 18288 19864 18294 19916
rect 18414 19864 18420 19916
rect 18472 19904 18478 19916
rect 18693 19907 18751 19913
rect 18693 19904 18705 19907
rect 18472 19876 18705 19904
rect 18472 19864 18478 19876
rect 18693 19873 18705 19876
rect 18739 19873 18751 19907
rect 18693 19867 18751 19873
rect 19702 19864 19708 19916
rect 19760 19904 19766 19916
rect 20257 19907 20315 19913
rect 20257 19904 20269 19907
rect 19760 19876 20269 19904
rect 19760 19864 19766 19876
rect 20257 19873 20269 19876
rect 20303 19873 20315 19907
rect 20257 19867 20315 19873
rect 20530 19864 20536 19916
rect 20588 19864 20594 19916
rect 22020 19904 22048 19935
rect 22554 19932 22560 19984
rect 22612 19972 22618 19984
rect 22833 19975 22891 19981
rect 22833 19972 22845 19975
rect 22612 19944 22845 19972
rect 22612 19932 22618 19944
rect 22833 19941 22845 19944
rect 22879 19941 22891 19975
rect 22833 19935 22891 19941
rect 22922 19932 22928 19984
rect 22980 19972 22986 19984
rect 24673 19975 24731 19981
rect 24673 19972 24685 19975
rect 22980 19944 24685 19972
rect 22980 19932 22986 19944
rect 24673 19941 24685 19944
rect 24719 19941 24731 19975
rect 24673 19935 24731 19941
rect 27522 19932 27528 19984
rect 27580 19972 27586 19984
rect 31386 19972 31392 19984
rect 27580 19944 31392 19972
rect 27580 19932 27586 19944
rect 31386 19932 31392 19944
rect 31444 19932 31450 19984
rect 23842 19904 23848 19916
rect 22020 19876 23848 19904
rect 23842 19864 23848 19876
rect 23900 19864 23906 19916
rect 25314 19864 25320 19916
rect 25372 19864 25378 19916
rect 26234 19864 26240 19916
rect 26292 19904 26298 19916
rect 28353 19907 28411 19913
rect 28353 19904 28365 19907
rect 26292 19876 28365 19904
rect 26292 19864 26298 19876
rect 28353 19873 28365 19876
rect 28399 19873 28411 19907
rect 29733 19907 29791 19913
rect 29733 19904 29745 19907
rect 28353 19867 28411 19873
rect 28460 19876 29745 19904
rect 9766 19836 9772 19848
rect 8404 19808 9772 19836
rect 4801 19771 4859 19777
rect 4801 19737 4813 19771
rect 4847 19737 4859 19771
rect 6270 19768 6276 19780
rect 6026 19740 6276 19768
rect 4801 19731 4859 19737
rect 4816 19700 4844 19731
rect 6270 19728 6276 19740
rect 6328 19768 6334 19780
rect 7466 19768 7472 19780
rect 6328 19740 7472 19768
rect 6328 19728 6334 19740
rect 7466 19728 7472 19740
rect 7524 19728 7530 19780
rect 6546 19700 6552 19712
rect 4816 19672 6552 19700
rect 6546 19660 6552 19672
rect 6604 19660 6610 19712
rect 6730 19660 6736 19712
rect 6788 19700 6794 19712
rect 8404 19700 8432 19808
rect 9766 19796 9772 19808
rect 9824 19796 9830 19848
rect 13262 19836 13268 19848
rect 11362 19808 13268 19836
rect 13262 19796 13268 19808
rect 13320 19836 13326 19848
rect 13320 19808 14320 19836
rect 13320 19796 13326 19808
rect 9306 19728 9312 19780
rect 9364 19728 9370 19780
rect 10229 19771 10287 19777
rect 10229 19737 10241 19771
rect 10275 19737 10287 19771
rect 10229 19731 10287 19737
rect 6788 19672 8432 19700
rect 8481 19703 8539 19709
rect 6788 19660 6794 19672
rect 8481 19669 8493 19703
rect 8527 19700 8539 19703
rect 8846 19700 8852 19712
rect 8527 19672 8852 19700
rect 8527 19669 8539 19672
rect 8481 19663 8539 19669
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 9398 19660 9404 19712
rect 9456 19660 9462 19712
rect 10244 19700 10272 19731
rect 11790 19728 11796 19780
rect 11848 19768 11854 19780
rect 12158 19768 12164 19780
rect 11848 19740 12164 19768
rect 11848 19728 11854 19740
rect 12158 19728 12164 19740
rect 12216 19768 12222 19780
rect 12253 19771 12311 19777
rect 12253 19768 12265 19771
rect 12216 19740 12265 19768
rect 12216 19728 12222 19740
rect 12253 19737 12265 19740
rect 12299 19737 12311 19771
rect 12253 19731 12311 19737
rect 13357 19771 13415 19777
rect 13357 19737 13369 19771
rect 13403 19768 13415 19771
rect 13538 19768 13544 19780
rect 13403 19740 13544 19768
rect 13403 19737 13415 19740
rect 13357 19731 13415 19737
rect 13538 19728 13544 19740
rect 13596 19728 13602 19780
rect 14292 19768 14320 19808
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 17313 19839 17371 19845
rect 17313 19805 17325 19839
rect 17359 19836 17371 19839
rect 18782 19836 18788 19848
rect 17359 19808 18788 19836
rect 17359 19805 17371 19808
rect 17313 19799 17371 19805
rect 18782 19796 18788 19808
rect 18840 19796 18846 19848
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19836 19671 19839
rect 19886 19836 19892 19848
rect 19659 19808 19892 19836
rect 19659 19805 19671 19808
rect 19613 19799 19671 19805
rect 19886 19796 19892 19808
rect 19944 19796 19950 19848
rect 21634 19796 21640 19848
rect 21692 19836 21698 19848
rect 23382 19836 23388 19848
rect 21692 19808 23388 19836
rect 21692 19796 21698 19808
rect 23382 19796 23388 19808
rect 23440 19796 23446 19848
rect 23753 19839 23811 19845
rect 23753 19805 23765 19839
rect 23799 19836 23811 19839
rect 25774 19836 25780 19848
rect 23799 19808 25780 19836
rect 23799 19805 23811 19808
rect 23753 19799 23811 19805
rect 25774 19796 25780 19808
rect 25832 19796 25838 19848
rect 25866 19796 25872 19848
rect 25924 19796 25930 19848
rect 27246 19796 27252 19848
rect 27304 19796 27310 19848
rect 27430 19796 27436 19848
rect 27488 19836 27494 19848
rect 28460 19836 28488 19876
rect 29733 19873 29745 19876
rect 29779 19873 29791 19907
rect 29733 19867 29791 19873
rect 31570 19864 31576 19916
rect 31628 19864 31634 19916
rect 27488 19808 28488 19836
rect 27488 19796 27494 19808
rect 29914 19796 29920 19848
rect 29972 19836 29978 19848
rect 30009 19839 30067 19845
rect 30009 19836 30021 19839
rect 29972 19808 30021 19836
rect 29972 19796 29978 19808
rect 30009 19805 30021 19808
rect 30055 19805 30067 19839
rect 30009 19799 30067 19805
rect 15286 19768 15292 19780
rect 14292 19740 15292 19768
rect 15286 19728 15292 19740
rect 15344 19728 15350 19780
rect 16132 19740 18184 19768
rect 11238 19700 11244 19712
rect 10244 19672 11244 19700
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 11514 19660 11520 19712
rect 11572 19700 11578 19712
rect 12345 19703 12403 19709
rect 12345 19700 12357 19703
rect 11572 19672 12357 19700
rect 11572 19660 11578 19672
rect 12345 19669 12357 19672
rect 12391 19669 12403 19703
rect 12345 19663 12403 19669
rect 12986 19660 12992 19712
rect 13044 19660 13050 19712
rect 13449 19703 13507 19709
rect 13449 19669 13461 19703
rect 13495 19700 13507 19703
rect 16132 19700 16160 19740
rect 18156 19709 18184 19740
rect 18230 19728 18236 19780
rect 18288 19768 18294 19780
rect 20806 19768 20812 19780
rect 18288 19740 20812 19768
rect 18288 19728 18294 19740
rect 20806 19728 20812 19740
rect 20864 19728 20870 19780
rect 24026 19768 24032 19780
rect 21836 19740 24032 19768
rect 13495 19672 16160 19700
rect 18141 19703 18199 19709
rect 13495 19669 13507 19672
rect 13449 19663 13507 19669
rect 18141 19669 18153 19703
rect 18187 19669 18199 19703
rect 18141 19663 18199 19669
rect 18414 19660 18420 19712
rect 18472 19700 18478 19712
rect 18509 19703 18567 19709
rect 18509 19700 18521 19703
rect 18472 19672 18521 19700
rect 18472 19660 18478 19672
rect 18509 19669 18521 19672
rect 18555 19669 18567 19703
rect 18509 19663 18567 19669
rect 18601 19703 18659 19709
rect 18601 19669 18613 19703
rect 18647 19700 18659 19703
rect 19518 19700 19524 19712
rect 18647 19672 19524 19700
rect 18647 19669 18659 19672
rect 18601 19663 18659 19669
rect 19518 19660 19524 19672
rect 19576 19660 19582 19712
rect 19705 19703 19763 19709
rect 19705 19669 19717 19703
rect 19751 19700 19763 19703
rect 19886 19700 19892 19712
rect 19751 19672 19892 19700
rect 19751 19669 19763 19672
rect 19705 19663 19763 19669
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 21358 19660 21364 19712
rect 21416 19700 21422 19712
rect 21836 19700 21864 19740
rect 24026 19728 24032 19740
rect 24084 19728 24090 19780
rect 25041 19771 25099 19777
rect 25041 19737 25053 19771
rect 25087 19768 25099 19771
rect 25498 19768 25504 19780
rect 25087 19740 25504 19768
rect 25087 19737 25099 19740
rect 25041 19731 25099 19737
rect 25498 19728 25504 19740
rect 25556 19728 25562 19780
rect 26142 19728 26148 19780
rect 26200 19728 26206 19780
rect 31481 19771 31539 19777
rect 27540 19740 31064 19768
rect 21416 19672 21864 19700
rect 21416 19660 21422 19672
rect 23658 19660 23664 19712
rect 23716 19660 23722 19712
rect 25133 19703 25191 19709
rect 25133 19669 25145 19703
rect 25179 19700 25191 19703
rect 27540 19700 27568 19740
rect 25179 19672 27568 19700
rect 25179 19669 25191 19672
rect 25133 19663 25191 19669
rect 27614 19660 27620 19712
rect 27672 19700 27678 19712
rect 31036 19709 31064 19740
rect 31481 19737 31493 19771
rect 31527 19768 31539 19771
rect 41322 19768 41328 19780
rect 31527 19740 41328 19768
rect 31527 19737 31539 19740
rect 31481 19731 31539 19737
rect 41322 19728 41328 19740
rect 41380 19728 41386 19780
rect 28583 19703 28641 19709
rect 28583 19700 28595 19703
rect 27672 19672 28595 19700
rect 27672 19660 27678 19672
rect 28583 19669 28595 19672
rect 28629 19669 28641 19703
rect 28583 19663 28641 19669
rect 31021 19703 31079 19709
rect 31021 19669 31033 19703
rect 31067 19669 31079 19703
rect 31021 19663 31079 19669
rect 31386 19660 31392 19712
rect 31444 19660 31450 19712
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 5626 19496 5632 19508
rect 2746 19468 5632 19496
rect 2746 19428 2774 19468
rect 5626 19456 5632 19468
rect 5684 19456 5690 19508
rect 5721 19499 5779 19505
rect 5721 19465 5733 19499
rect 5767 19496 5779 19499
rect 6822 19496 6828 19508
rect 5767 19468 6828 19496
rect 5767 19465 5779 19468
rect 5721 19459 5779 19465
rect 6822 19456 6828 19468
rect 6880 19456 6886 19508
rect 8754 19456 8760 19508
rect 8812 19496 8818 19508
rect 9950 19496 9956 19508
rect 8812 19468 9956 19496
rect 8812 19456 8818 19468
rect 9950 19456 9956 19468
rect 10008 19456 10014 19508
rect 14550 19496 14556 19508
rect 11992 19468 14556 19496
rect 11992 19440 12020 19468
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 20622 19496 20628 19508
rect 14752 19468 20628 19496
rect 1780 19400 2774 19428
rect 1780 19369 1808 19400
rect 4522 19388 4528 19440
rect 4580 19388 4586 19440
rect 6914 19428 6920 19440
rect 5368 19400 6920 19428
rect 1765 19363 1823 19369
rect 1765 19329 1777 19363
rect 1811 19329 1823 19363
rect 1765 19323 1823 19329
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19360 3663 19363
rect 5368 19360 5396 19400
rect 6914 19388 6920 19400
rect 6972 19388 6978 19440
rect 8570 19388 8576 19440
rect 8628 19428 8634 19440
rect 10137 19431 10195 19437
rect 10137 19428 10149 19431
rect 8628 19400 10149 19428
rect 8628 19388 8634 19400
rect 10137 19397 10149 19400
rect 10183 19397 10195 19431
rect 11974 19428 11980 19440
rect 10137 19391 10195 19397
rect 11716 19400 11980 19428
rect 3651 19332 5396 19360
rect 5629 19363 5687 19369
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 5629 19329 5641 19363
rect 5675 19360 5687 19363
rect 6730 19360 6736 19372
rect 5675 19332 6736 19360
rect 5675 19329 5687 19332
rect 5629 19323 5687 19329
rect 6730 19320 6736 19332
rect 6788 19320 6794 19372
rect 7006 19360 7012 19372
rect 7064 19369 7070 19372
rect 6974 19332 7012 19360
rect 7006 19320 7012 19332
rect 7064 19323 7074 19369
rect 7064 19320 7070 19323
rect 8386 19320 8392 19372
rect 8444 19320 8450 19372
rect 8662 19320 8668 19372
rect 8720 19360 8726 19372
rect 11716 19369 11744 19400
rect 11974 19388 11980 19400
rect 12032 19388 12038 19440
rect 13354 19428 13360 19440
rect 13202 19400 13360 19428
rect 13354 19388 13360 19400
rect 13412 19388 13418 19440
rect 13722 19388 13728 19440
rect 13780 19428 13786 19440
rect 14645 19431 14703 19437
rect 14645 19428 14657 19431
rect 13780 19400 14657 19428
rect 13780 19388 13786 19400
rect 14645 19397 14657 19400
rect 14691 19397 14703 19431
rect 14645 19391 14703 19397
rect 9217 19363 9275 19369
rect 9217 19360 9229 19363
rect 8720 19332 9229 19360
rect 8720 19320 8726 19332
rect 9217 19329 9229 19332
rect 9263 19329 9275 19363
rect 9217 19323 9275 19329
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19329 11759 19363
rect 13909 19363 13967 19369
rect 13909 19360 13921 19363
rect 11701 19323 11759 19329
rect 13740 19332 13921 19360
rect 13740 19304 13768 19332
rect 13909 19329 13921 19332
rect 13955 19360 13967 19363
rect 14752 19360 14780 19468
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 21453 19499 21511 19505
rect 21453 19496 21465 19499
rect 20864 19468 21465 19496
rect 20864 19456 20870 19468
rect 21453 19465 21465 19468
rect 21499 19465 21511 19499
rect 21453 19459 21511 19465
rect 22370 19456 22376 19508
rect 22428 19496 22434 19508
rect 22465 19499 22523 19505
rect 22465 19496 22477 19499
rect 22428 19468 22477 19496
rect 22428 19456 22434 19468
rect 22465 19465 22477 19468
rect 22511 19465 22523 19499
rect 22465 19459 22523 19465
rect 22554 19456 22560 19508
rect 22612 19496 22618 19508
rect 22833 19499 22891 19505
rect 22833 19496 22845 19499
rect 22612 19468 22845 19496
rect 22612 19456 22618 19468
rect 22833 19465 22845 19468
rect 22879 19465 22891 19499
rect 22833 19459 22891 19465
rect 22925 19499 22983 19505
rect 22925 19465 22937 19499
rect 22971 19496 22983 19499
rect 23566 19496 23572 19508
rect 22971 19468 23572 19496
rect 22971 19465 22983 19468
rect 22925 19459 22983 19465
rect 23566 19456 23572 19468
rect 23624 19456 23630 19508
rect 23661 19499 23719 19505
rect 23661 19465 23673 19499
rect 23707 19465 23719 19499
rect 23661 19459 23719 19465
rect 15378 19388 15384 19440
rect 15436 19428 15442 19440
rect 15749 19431 15807 19437
rect 15749 19428 15761 19431
rect 15436 19400 15761 19428
rect 15436 19388 15442 19400
rect 15749 19397 15761 19400
rect 15795 19428 15807 19431
rect 15838 19428 15844 19440
rect 15795 19400 15844 19428
rect 15795 19397 15807 19400
rect 15749 19391 15807 19397
rect 15838 19388 15844 19400
rect 15896 19388 15902 19440
rect 17126 19388 17132 19440
rect 17184 19428 17190 19440
rect 18690 19428 18696 19440
rect 17184 19400 17356 19428
rect 17184 19388 17190 19400
rect 13955 19332 14780 19360
rect 13955 19329 13967 19332
rect 13909 19323 13967 19329
rect 15654 19320 15660 19372
rect 15712 19320 15718 19372
rect 16758 19320 16764 19372
rect 16816 19360 16822 19372
rect 17328 19369 17356 19400
rect 17420 19400 18696 19428
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 16816 19332 17233 19360
rect 16816 19320 16822 19332
rect 17221 19329 17233 19332
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19329 17371 19363
rect 17313 19323 17371 19329
rect 2038 19252 2044 19304
rect 2096 19252 2102 19304
rect 3418 19252 3424 19304
rect 3476 19292 3482 19304
rect 5813 19295 5871 19301
rect 5813 19292 5825 19295
rect 3476 19264 5825 19292
rect 3476 19252 3482 19264
rect 5813 19261 5825 19264
rect 5859 19261 5871 19295
rect 5813 19255 5871 19261
rect 7285 19295 7343 19301
rect 7285 19261 7297 19295
rect 7331 19292 7343 19295
rect 7650 19292 7656 19304
rect 7331 19264 7656 19292
rect 7331 19261 7343 19264
rect 7285 19255 7343 19261
rect 4246 19116 4252 19168
rect 4304 19156 4310 19168
rect 5261 19159 5319 19165
rect 5261 19156 5273 19159
rect 4304 19128 5273 19156
rect 4304 19116 4310 19128
rect 5261 19125 5273 19128
rect 5307 19125 5319 19159
rect 5828 19156 5856 19255
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 11977 19295 12035 19301
rect 11977 19261 11989 19295
rect 12023 19292 12035 19295
rect 13630 19292 13636 19304
rect 12023 19264 13636 19292
rect 12023 19261 12035 19264
rect 11977 19255 12035 19261
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 13722 19252 13728 19304
rect 13780 19252 13786 19304
rect 15838 19252 15844 19304
rect 15896 19252 15902 19304
rect 16298 19252 16304 19304
rect 16356 19292 16362 19304
rect 17420 19292 17448 19400
rect 18690 19388 18696 19400
rect 18748 19428 18754 19440
rect 21634 19428 21640 19440
rect 18748 19400 19748 19428
rect 21206 19400 21640 19428
rect 18748 19388 18754 19400
rect 18509 19363 18567 19369
rect 18509 19329 18521 19363
rect 18555 19360 18567 19363
rect 18874 19360 18880 19372
rect 18555 19332 18880 19360
rect 18555 19329 18567 19332
rect 18509 19323 18567 19329
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 19334 19360 19340 19372
rect 18984 19332 19340 19360
rect 18984 19304 19012 19332
rect 19334 19320 19340 19332
rect 19392 19320 19398 19372
rect 19720 19304 19748 19400
rect 21634 19388 21640 19400
rect 21692 19388 21698 19440
rect 21726 19388 21732 19440
rect 21784 19428 21790 19440
rect 22646 19428 22652 19440
rect 21784 19400 22652 19428
rect 21784 19388 21790 19400
rect 22646 19388 22652 19400
rect 22704 19388 22710 19440
rect 23676 19428 23704 19459
rect 24026 19456 24032 19508
rect 24084 19456 24090 19508
rect 27617 19499 27675 19505
rect 27617 19465 27629 19499
rect 27663 19496 27675 19499
rect 35066 19496 35072 19508
rect 27663 19468 35072 19496
rect 27663 19465 27675 19468
rect 27617 19459 27675 19465
rect 35066 19456 35072 19468
rect 35124 19456 35130 19508
rect 23584 19400 23704 19428
rect 23584 19360 23612 19400
rect 29638 19388 29644 19440
rect 29696 19388 29702 19440
rect 23584 19332 23704 19360
rect 16356 19264 17448 19292
rect 17497 19295 17555 19301
rect 16356 19252 16362 19264
rect 17497 19261 17509 19295
rect 17543 19292 17555 19295
rect 18046 19292 18052 19304
rect 17543 19264 18052 19292
rect 17543 19261 17555 19264
rect 17497 19255 17555 19261
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 18598 19252 18604 19304
rect 18656 19252 18662 19304
rect 18785 19295 18843 19301
rect 18785 19261 18797 19295
rect 18831 19261 18843 19295
rect 18785 19255 18843 19261
rect 8478 19184 8484 19236
rect 8536 19224 8542 19236
rect 11422 19224 11428 19236
rect 8536 19196 11428 19224
rect 8536 19184 8542 19196
rect 11422 19184 11428 19196
rect 11480 19184 11486 19236
rect 12986 19184 12992 19236
rect 13044 19224 13050 19236
rect 18322 19224 18328 19236
rect 13044 19196 16988 19224
rect 13044 19184 13050 19196
rect 7282 19156 7288 19168
rect 5828 19128 7288 19156
rect 5261 19119 5319 19125
rect 7282 19116 7288 19128
rect 7340 19116 7346 19168
rect 11238 19116 11244 19168
rect 11296 19156 11302 19168
rect 13449 19159 13507 19165
rect 13449 19156 13461 19159
rect 11296 19128 13461 19156
rect 11296 19116 11302 19128
rect 13449 19125 13461 19128
rect 13495 19125 13507 19159
rect 13449 19119 13507 19125
rect 15286 19116 15292 19168
rect 15344 19116 15350 19168
rect 15930 19116 15936 19168
rect 15988 19156 15994 19168
rect 16666 19156 16672 19168
rect 15988 19128 16672 19156
rect 15988 19116 15994 19128
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 16850 19116 16856 19168
rect 16908 19116 16914 19168
rect 16960 19156 16988 19196
rect 18064 19196 18328 19224
rect 18064 19156 18092 19196
rect 18322 19184 18328 19196
rect 18380 19184 18386 19236
rect 18800 19224 18828 19255
rect 18966 19252 18972 19304
rect 19024 19252 19030 19304
rect 19702 19252 19708 19304
rect 19760 19252 19766 19304
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 19812 19264 19993 19292
rect 18800 19196 19334 19224
rect 16960 19128 18092 19156
rect 18138 19116 18144 19168
rect 18196 19116 18202 19168
rect 19306 19156 19334 19196
rect 19610 19184 19616 19236
rect 19668 19224 19674 19236
rect 19812 19224 19840 19264
rect 19981 19261 19993 19264
rect 20027 19292 20039 19295
rect 20346 19292 20352 19304
rect 20027 19264 20352 19292
rect 20027 19261 20039 19264
rect 19981 19255 20039 19261
rect 20346 19252 20352 19264
rect 20404 19252 20410 19304
rect 23109 19295 23167 19301
rect 23109 19261 23121 19295
rect 23155 19261 23167 19295
rect 23109 19255 23167 19261
rect 19668 19196 19840 19224
rect 23124 19224 23152 19255
rect 23566 19252 23572 19304
rect 23624 19292 23630 19304
rect 23676 19292 23704 19332
rect 24118 19320 24124 19372
rect 24176 19320 24182 19372
rect 25038 19320 25044 19372
rect 25096 19320 25102 19372
rect 27614 19320 27620 19372
rect 27672 19360 27678 19372
rect 27801 19363 27859 19369
rect 27801 19360 27813 19363
rect 27672 19332 27813 19360
rect 27672 19320 27678 19332
rect 27801 19329 27813 19332
rect 27847 19329 27859 19363
rect 27801 19323 27859 19329
rect 23624 19264 23704 19292
rect 24305 19295 24363 19301
rect 23624 19252 23630 19264
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 24946 19292 24952 19304
rect 24351 19264 24952 19292
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 24946 19252 24952 19264
rect 25004 19252 25010 19304
rect 25866 19252 25872 19304
rect 25924 19252 25930 19304
rect 26326 19252 26332 19304
rect 26384 19292 26390 19304
rect 26605 19295 26663 19301
rect 26605 19292 26617 19295
rect 26384 19264 26617 19292
rect 26384 19252 26390 19264
rect 26605 19261 26617 19264
rect 26651 19261 26663 19295
rect 26605 19255 26663 19261
rect 28350 19252 28356 19304
rect 28408 19252 28414 19304
rect 28629 19295 28687 19301
rect 28629 19292 28641 19295
rect 28460 19264 28641 19292
rect 26142 19224 26148 19236
rect 23124 19196 26148 19224
rect 19668 19184 19674 19196
rect 26142 19184 26148 19196
rect 26200 19184 26206 19236
rect 26418 19184 26424 19236
rect 26476 19224 26482 19236
rect 28460 19224 28488 19264
rect 28629 19261 28641 19264
rect 28675 19261 28687 19295
rect 28629 19255 28687 19261
rect 30926 19224 30932 19236
rect 26476 19196 28488 19224
rect 29656 19196 30932 19224
rect 26476 19184 26482 19196
rect 19978 19156 19984 19168
rect 19306 19128 19984 19156
rect 19978 19116 19984 19128
rect 20036 19116 20042 19168
rect 20162 19116 20168 19168
rect 20220 19156 20226 19168
rect 25406 19156 25412 19168
rect 20220 19128 25412 19156
rect 20220 19116 20226 19128
rect 25406 19116 25412 19128
rect 25464 19116 25470 19168
rect 25774 19116 25780 19168
rect 25832 19156 25838 19168
rect 28442 19156 28448 19168
rect 25832 19128 28448 19156
rect 25832 19116 25838 19128
rect 28442 19116 28448 19128
rect 28500 19156 28506 19168
rect 29656 19156 29684 19196
rect 30926 19184 30932 19196
rect 30984 19184 30990 19236
rect 28500 19128 29684 19156
rect 28500 19116 28506 19128
rect 30098 19116 30104 19168
rect 30156 19116 30162 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 11514 18952 11520 18964
rect 2746 18924 11520 18952
rect 2746 18816 2774 18924
rect 11514 18912 11520 18924
rect 11572 18912 11578 18964
rect 12066 18912 12072 18964
rect 12124 18912 12130 18964
rect 18138 18952 18144 18964
rect 12406 18924 14320 18952
rect 12406 18884 12434 18924
rect 6104 18856 7512 18884
rect 1780 18788 2774 18816
rect 1780 18757 1808 18788
rect 3326 18776 3332 18828
rect 3384 18816 3390 18828
rect 6104 18816 6132 18856
rect 6270 18816 6276 18828
rect 3384 18788 6132 18816
rect 6196 18788 6276 18816
rect 3384 18776 3390 18788
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18717 1823 18751
rect 1765 18711 1823 18717
rect 4341 18751 4399 18757
rect 4341 18717 4353 18751
rect 4387 18748 4399 18751
rect 4706 18748 4712 18760
rect 4387 18720 4712 18748
rect 4387 18717 4399 18720
rect 4341 18711 4399 18717
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 4798 18708 4804 18760
rect 4856 18708 4862 18760
rect 6196 18734 6224 18788
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 6546 18776 6552 18828
rect 6604 18816 6610 18828
rect 7484 18825 7512 18856
rect 8220 18856 12434 18884
rect 7469 18819 7527 18825
rect 6604 18788 7144 18816
rect 6604 18776 6610 18788
rect 2498 18640 2504 18692
rect 2556 18640 2562 18692
rect 5077 18683 5135 18689
rect 5077 18649 5089 18683
rect 5123 18680 5135 18683
rect 5166 18680 5172 18692
rect 5123 18652 5172 18680
rect 5123 18649 5135 18652
rect 5077 18643 5135 18649
rect 5166 18640 5172 18652
rect 5224 18640 5230 18692
rect 7116 18680 7144 18788
rect 7469 18785 7481 18819
rect 7515 18785 7527 18819
rect 7469 18779 7527 18785
rect 7193 18751 7251 18757
rect 7193 18717 7205 18751
rect 7239 18748 7251 18751
rect 8220 18748 8248 18856
rect 12526 18844 12532 18896
rect 12584 18884 12590 18896
rect 14090 18884 14096 18896
rect 12584 18856 14096 18884
rect 12584 18844 12590 18856
rect 14090 18844 14096 18856
rect 14148 18844 14154 18896
rect 8294 18776 8300 18828
rect 8352 18816 8358 18828
rect 8754 18816 8760 18828
rect 8352 18788 8760 18816
rect 8352 18776 8358 18788
rect 8754 18776 8760 18788
rect 8812 18816 8818 18828
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 8812 18788 9689 18816
rect 8812 18776 8818 18788
rect 9677 18785 9689 18788
rect 9723 18785 9735 18819
rect 9677 18779 9735 18785
rect 11238 18776 11244 18828
rect 11296 18816 11302 18828
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 11296 18788 11437 18816
rect 11296 18776 11302 18788
rect 11425 18785 11437 18788
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11882 18816 11888 18828
rect 11572 18788 11888 18816
rect 11572 18776 11578 18788
rect 11882 18776 11888 18788
rect 11940 18816 11946 18828
rect 12250 18816 12256 18828
rect 11940 18788 12256 18816
rect 11940 18776 11946 18788
rect 12250 18776 12256 18788
rect 12308 18776 12314 18828
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 12621 18819 12679 18825
rect 12621 18816 12633 18819
rect 12492 18788 12633 18816
rect 12492 18776 12498 18788
rect 12621 18785 12633 18788
rect 12667 18785 12679 18819
rect 12621 18779 12679 18785
rect 12894 18776 12900 18828
rect 12952 18816 12958 18828
rect 13538 18816 13544 18828
rect 12952 18788 13544 18816
rect 12952 18776 12958 18788
rect 13538 18776 13544 18788
rect 13596 18776 13602 18828
rect 7239 18720 8248 18748
rect 9493 18751 9551 18757
rect 7239 18717 7251 18720
rect 7193 18711 7251 18717
rect 9493 18717 9505 18751
rect 9539 18748 9551 18751
rect 10502 18748 10508 18760
rect 9539 18720 10508 18748
rect 9539 18717 9551 18720
rect 9493 18711 9551 18717
rect 10502 18708 10508 18720
rect 10560 18708 10566 18760
rect 13170 18748 13176 18760
rect 11256 18720 13176 18748
rect 8570 18680 8576 18692
rect 7116 18652 8576 18680
rect 8570 18640 8576 18652
rect 8628 18640 8634 18692
rect 11256 18689 11284 18720
rect 13170 18708 13176 18720
rect 13228 18708 13234 18760
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18748 13415 18751
rect 13906 18748 13912 18760
rect 13403 18720 13912 18748
rect 13403 18717 13415 18720
rect 13357 18711 13415 18717
rect 13906 18708 13912 18720
rect 13964 18708 13970 18760
rect 10413 18683 10471 18689
rect 10413 18649 10425 18683
rect 10459 18680 10471 18683
rect 11241 18683 11299 18689
rect 11241 18680 11253 18683
rect 10459 18652 11253 18680
rect 10459 18649 10471 18652
rect 10413 18643 10471 18649
rect 11241 18649 11253 18652
rect 11287 18649 11299 18683
rect 11241 18643 11299 18649
rect 11422 18640 11428 18692
rect 11480 18680 11486 18692
rect 13541 18683 13599 18689
rect 13541 18680 13553 18683
rect 11480 18652 13553 18680
rect 11480 18640 11486 18652
rect 13541 18649 13553 18652
rect 13587 18649 13599 18683
rect 14292 18680 14320 18924
rect 14476 18924 18144 18952
rect 14476 18757 14504 18924
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 19978 18912 19984 18964
rect 20036 18952 20042 18964
rect 22925 18955 22983 18961
rect 22925 18952 22937 18955
rect 20036 18924 22937 18952
rect 20036 18912 20042 18924
rect 22925 18921 22937 18924
rect 22971 18921 22983 18955
rect 22925 18915 22983 18921
rect 23658 18912 23664 18964
rect 23716 18952 23722 18964
rect 24765 18955 24823 18961
rect 24765 18952 24777 18955
rect 23716 18924 24777 18952
rect 23716 18912 23722 18924
rect 24765 18921 24777 18924
rect 24811 18921 24823 18955
rect 24765 18915 24823 18921
rect 26142 18912 26148 18964
rect 26200 18952 26206 18964
rect 27157 18955 27215 18961
rect 27157 18952 27169 18955
rect 26200 18924 27169 18952
rect 26200 18912 26206 18924
rect 27157 18921 27169 18924
rect 27203 18921 27215 18955
rect 27157 18915 27215 18921
rect 28810 18912 28816 18964
rect 28868 18912 28874 18964
rect 29840 18924 35894 18952
rect 14642 18844 14648 18896
rect 14700 18844 14706 18896
rect 17218 18844 17224 18896
rect 17276 18884 17282 18896
rect 17865 18887 17923 18893
rect 17865 18884 17877 18887
rect 17276 18856 17877 18884
rect 17276 18844 17282 18856
rect 17865 18853 17877 18856
rect 17911 18853 17923 18887
rect 20806 18884 20812 18896
rect 17865 18847 17923 18853
rect 18156 18856 20812 18884
rect 15105 18819 15163 18825
rect 15105 18785 15117 18819
rect 15151 18816 15163 18819
rect 16114 18816 16120 18828
rect 15151 18788 16120 18816
rect 15151 18785 15163 18788
rect 15105 18779 15163 18785
rect 16114 18776 16120 18788
rect 16172 18776 16178 18828
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18717 14519 18751
rect 14461 18711 14519 18717
rect 16666 18708 16672 18760
rect 16724 18708 16730 18760
rect 17770 18708 17776 18760
rect 17828 18748 17834 18760
rect 18156 18748 18184 18856
rect 20806 18844 20812 18856
rect 20864 18844 20870 18896
rect 23385 18887 23443 18893
rect 23385 18853 23397 18887
rect 23431 18853 23443 18887
rect 23385 18847 23443 18853
rect 18322 18776 18328 18828
rect 18380 18816 18386 18828
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 18380 18788 18429 18816
rect 18380 18776 18386 18788
rect 18417 18785 18429 18788
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 20441 18819 20499 18825
rect 20441 18816 20453 18819
rect 19760 18788 20453 18816
rect 19760 18776 19766 18788
rect 20441 18785 20453 18788
rect 20487 18785 20499 18819
rect 20441 18779 20499 18785
rect 21174 18776 21180 18828
rect 21232 18776 21238 18828
rect 21450 18776 21456 18828
rect 21508 18776 21514 18828
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 23400 18816 23428 18847
rect 27062 18844 27068 18896
rect 27120 18884 27126 18896
rect 29733 18887 29791 18893
rect 29733 18884 29745 18887
rect 27120 18856 29745 18884
rect 27120 18844 27126 18856
rect 29733 18853 29745 18856
rect 29779 18853 29791 18887
rect 29733 18847 29791 18853
rect 22152 18788 23428 18816
rect 25409 18819 25467 18825
rect 22152 18776 22158 18788
rect 25409 18785 25421 18819
rect 25455 18816 25467 18819
rect 25774 18816 25780 18828
rect 25455 18788 25780 18816
rect 25455 18785 25467 18788
rect 25409 18779 25467 18785
rect 25774 18776 25780 18788
rect 25832 18776 25838 18828
rect 27522 18776 27528 18828
rect 27580 18816 27586 18828
rect 28169 18819 28227 18825
rect 28169 18816 28181 18819
rect 27580 18788 28181 18816
rect 27580 18776 27586 18788
rect 28169 18785 28181 18788
rect 28215 18785 28227 18819
rect 29840 18816 29868 18924
rect 31021 18887 31079 18893
rect 31021 18853 31033 18887
rect 31067 18884 31079 18887
rect 34422 18884 34428 18896
rect 31067 18856 34428 18884
rect 31067 18853 31079 18856
rect 31021 18847 31079 18853
rect 28169 18779 28227 18785
rect 28276 18788 29868 18816
rect 17828 18720 18184 18748
rect 18233 18751 18291 18757
rect 17828 18708 17834 18720
rect 18233 18717 18245 18751
rect 18279 18748 18291 18751
rect 18690 18748 18696 18760
rect 18279 18720 18696 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 23566 18708 23572 18760
rect 23624 18708 23630 18760
rect 27154 18708 27160 18760
rect 27212 18748 27218 18760
rect 28276 18748 28304 18788
rect 30006 18776 30012 18828
rect 30064 18816 30070 18828
rect 30285 18819 30343 18825
rect 30285 18816 30297 18819
rect 30064 18788 30297 18816
rect 30064 18776 30070 18788
rect 30285 18785 30297 18788
rect 30331 18785 30343 18819
rect 30285 18779 30343 18785
rect 27212 18720 28304 18748
rect 27212 18708 27218 18720
rect 28994 18708 29000 18760
rect 29052 18708 29058 18760
rect 29086 18708 29092 18760
rect 29144 18748 29150 18760
rect 30101 18751 30159 18757
rect 30101 18748 30113 18751
rect 29144 18720 30113 18748
rect 29144 18708 29150 18720
rect 30101 18717 30113 18720
rect 30147 18748 30159 18751
rect 31036 18748 31064 18847
rect 34422 18844 34428 18856
rect 34480 18844 34486 18896
rect 35866 18884 35894 18924
rect 45370 18884 45376 18896
rect 35866 18856 45376 18884
rect 45370 18844 45376 18856
rect 45428 18844 45434 18896
rect 30147 18720 31064 18748
rect 30147 18717 30159 18720
rect 30101 18711 30159 18717
rect 14292 18652 14688 18680
rect 13541 18643 13599 18649
rect 3326 18572 3332 18624
rect 3384 18612 3390 18624
rect 4157 18615 4215 18621
rect 4157 18612 4169 18615
rect 3384 18584 4169 18612
rect 3384 18572 3390 18584
rect 4157 18581 4169 18584
rect 4203 18581 4215 18615
rect 4157 18575 4215 18581
rect 7282 18572 7288 18624
rect 7340 18612 7346 18624
rect 9125 18615 9183 18621
rect 9125 18612 9137 18615
rect 7340 18584 9137 18612
rect 7340 18572 7346 18584
rect 9125 18581 9137 18584
rect 9171 18581 9183 18615
rect 9125 18575 9183 18581
rect 9585 18615 9643 18621
rect 9585 18581 9597 18615
rect 9631 18612 9643 18615
rect 9674 18612 9680 18624
rect 9631 18584 9680 18612
rect 9631 18581 9643 18584
rect 9585 18575 9643 18581
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 10870 18572 10876 18624
rect 10928 18572 10934 18624
rect 11333 18615 11391 18621
rect 11333 18581 11345 18615
rect 11379 18612 11391 18615
rect 11882 18612 11888 18624
rect 11379 18584 11888 18612
rect 11379 18581 11391 18584
rect 11333 18575 11391 18581
rect 11882 18572 11888 18584
rect 11940 18572 11946 18624
rect 12066 18572 12072 18624
rect 12124 18612 12130 18624
rect 12437 18615 12495 18621
rect 12437 18612 12449 18615
rect 12124 18584 12449 18612
rect 12124 18572 12130 18584
rect 12437 18581 12449 18584
rect 12483 18581 12495 18615
rect 12437 18575 12495 18581
rect 12529 18615 12587 18621
rect 12529 18581 12541 18615
rect 12575 18612 12587 18615
rect 14458 18612 14464 18624
rect 12575 18584 14464 18612
rect 12575 18581 12587 18584
rect 12529 18575 12587 18581
rect 14458 18572 14464 18584
rect 14516 18572 14522 18624
rect 14660 18612 14688 18652
rect 15010 18640 15016 18692
rect 15068 18680 15074 18692
rect 15381 18683 15439 18689
rect 15381 18680 15393 18683
rect 15068 18652 15393 18680
rect 15068 18640 15074 18652
rect 15381 18649 15393 18652
rect 15427 18680 15439 18683
rect 15470 18680 15476 18692
rect 15427 18652 15476 18680
rect 15427 18649 15439 18652
rect 15381 18643 15439 18649
rect 15470 18640 15476 18652
rect 15528 18640 15534 18692
rect 16684 18680 16712 18708
rect 17678 18680 17684 18692
rect 16606 18652 17684 18680
rect 17678 18640 17684 18652
rect 17736 18640 17742 18692
rect 18046 18640 18052 18692
rect 18104 18680 18110 18692
rect 18874 18680 18880 18692
rect 18104 18652 18880 18680
rect 18104 18640 18110 18652
rect 18874 18640 18880 18652
rect 18932 18640 18938 18692
rect 19702 18640 19708 18692
rect 19760 18680 19766 18692
rect 20622 18680 20628 18692
rect 19760 18652 20628 18680
rect 19760 18640 19766 18652
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 23842 18680 23848 18692
rect 22678 18652 23848 18680
rect 23842 18640 23848 18652
rect 23900 18680 23906 18692
rect 24486 18680 24492 18692
rect 23900 18652 24492 18680
rect 23900 18640 23906 18652
rect 24486 18640 24492 18652
rect 24544 18640 24550 18692
rect 25682 18640 25688 18692
rect 25740 18640 25746 18692
rect 27246 18680 27252 18692
rect 26910 18652 27252 18680
rect 27246 18640 27252 18652
rect 27304 18640 27310 18692
rect 28077 18683 28135 18689
rect 28077 18649 28089 18683
rect 28123 18680 28135 18683
rect 30282 18680 30288 18692
rect 28123 18652 30288 18680
rect 28123 18649 28135 18652
rect 28077 18643 28135 18649
rect 30282 18640 30288 18652
rect 30340 18640 30346 18692
rect 30374 18640 30380 18692
rect 30432 18680 30438 18692
rect 48498 18680 48504 18692
rect 30432 18652 48504 18680
rect 30432 18640 30438 18652
rect 48498 18640 48504 18652
rect 48556 18640 48562 18692
rect 15562 18612 15568 18624
rect 14660 18584 15568 18612
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 16666 18572 16672 18624
rect 16724 18612 16730 18624
rect 16853 18615 16911 18621
rect 16853 18612 16865 18615
rect 16724 18584 16865 18612
rect 16724 18572 16730 18584
rect 16853 18581 16865 18584
rect 16899 18581 16911 18615
rect 16853 18575 16911 18581
rect 18322 18572 18328 18624
rect 18380 18612 18386 18624
rect 21818 18612 21824 18624
rect 18380 18584 21824 18612
rect 18380 18572 18386 18584
rect 21818 18572 21824 18584
rect 21876 18572 21882 18624
rect 22922 18572 22928 18624
rect 22980 18612 22986 18624
rect 24854 18612 24860 18624
rect 22980 18584 24860 18612
rect 22980 18572 22986 18584
rect 24854 18572 24860 18584
rect 24912 18572 24918 18624
rect 25314 18572 25320 18624
rect 25372 18612 25378 18624
rect 26602 18612 26608 18624
rect 25372 18584 26608 18612
rect 25372 18572 25378 18584
rect 26602 18572 26608 18584
rect 26660 18572 26666 18624
rect 26694 18572 26700 18624
rect 26752 18612 26758 18624
rect 27617 18615 27675 18621
rect 27617 18612 27629 18615
rect 26752 18584 27629 18612
rect 26752 18572 26758 18584
rect 27617 18581 27629 18584
rect 27663 18581 27675 18615
rect 27617 18575 27675 18581
rect 27706 18572 27712 18624
rect 27764 18612 27770 18624
rect 27985 18615 28043 18621
rect 27985 18612 27997 18615
rect 27764 18584 27997 18612
rect 27764 18572 27770 18584
rect 27985 18581 27997 18584
rect 28031 18581 28043 18615
rect 27985 18575 28043 18581
rect 29454 18572 29460 18624
rect 29512 18612 29518 18624
rect 30193 18615 30251 18621
rect 30193 18612 30205 18615
rect 29512 18584 30205 18612
rect 29512 18572 29518 18584
rect 30193 18581 30205 18584
rect 30239 18581 30251 18615
rect 30193 18575 30251 18581
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 5074 18368 5080 18420
rect 5132 18408 5138 18420
rect 5721 18411 5779 18417
rect 5721 18408 5733 18411
rect 5132 18380 5733 18408
rect 5132 18368 5138 18380
rect 5721 18377 5733 18380
rect 5767 18408 5779 18411
rect 10873 18411 10931 18417
rect 10873 18408 10885 18411
rect 5767 18380 10885 18408
rect 5767 18377 5779 18380
rect 5721 18371 5779 18377
rect 10873 18377 10885 18380
rect 10919 18377 10931 18411
rect 10873 18371 10931 18377
rect 10962 18368 10968 18420
rect 11020 18408 11026 18420
rect 12066 18408 12072 18420
rect 11020 18380 12072 18408
rect 11020 18368 11026 18380
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 12492 18380 14688 18408
rect 12492 18368 12498 18380
rect 2222 18300 2228 18352
rect 2280 18340 2286 18352
rect 8573 18343 8631 18349
rect 2280 18312 3924 18340
rect 2280 18300 2286 18312
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 1946 18272 1952 18284
rect 1811 18244 1952 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 3418 18232 3424 18284
rect 3476 18232 3482 18284
rect 2774 18164 2780 18216
rect 2832 18164 2838 18216
rect 3896 18213 3924 18312
rect 8573 18309 8585 18343
rect 8619 18340 8631 18343
rect 9122 18340 9128 18352
rect 8619 18312 9128 18340
rect 8619 18309 8631 18312
rect 8573 18303 8631 18309
rect 9122 18300 9128 18312
rect 9180 18340 9186 18352
rect 13722 18340 13728 18352
rect 9180 18312 13728 18340
rect 9180 18300 9186 18312
rect 13722 18300 13728 18312
rect 13780 18300 13786 18352
rect 14550 18300 14556 18352
rect 14608 18300 14614 18352
rect 14660 18340 14688 18380
rect 15102 18368 15108 18420
rect 15160 18368 15166 18420
rect 15565 18411 15623 18417
rect 15565 18377 15577 18411
rect 15611 18408 15623 18411
rect 19705 18411 19763 18417
rect 19705 18408 19717 18411
rect 15611 18380 19717 18408
rect 15611 18377 15623 18380
rect 15565 18371 15623 18377
rect 19705 18377 19717 18380
rect 19751 18377 19763 18411
rect 19705 18371 19763 18377
rect 20073 18411 20131 18417
rect 20073 18377 20085 18411
rect 20119 18408 20131 18411
rect 20162 18408 20168 18420
rect 20119 18380 20168 18408
rect 20119 18377 20131 18380
rect 20073 18371 20131 18377
rect 20162 18368 20168 18380
rect 20220 18368 20226 18420
rect 20346 18368 20352 18420
rect 20404 18408 20410 18420
rect 24857 18411 24915 18417
rect 24857 18408 24869 18411
rect 20404 18380 24869 18408
rect 20404 18368 20410 18380
rect 24857 18377 24869 18380
rect 24903 18377 24915 18411
rect 24857 18371 24915 18377
rect 25130 18368 25136 18420
rect 25188 18408 25194 18420
rect 30285 18411 30343 18417
rect 30285 18408 30297 18411
rect 25188 18380 30297 18408
rect 25188 18368 25194 18380
rect 30285 18377 30297 18380
rect 30331 18377 30343 18411
rect 30285 18371 30343 18377
rect 30745 18411 30803 18417
rect 30745 18377 30757 18411
rect 30791 18408 30803 18411
rect 37734 18408 37740 18420
rect 30791 18380 37740 18408
rect 30791 18377 30803 18380
rect 30745 18371 30803 18377
rect 37734 18368 37740 18380
rect 37792 18368 37798 18420
rect 17405 18343 17463 18349
rect 17405 18340 17417 18343
rect 14660 18312 17417 18340
rect 17405 18309 17417 18312
rect 17451 18309 17463 18343
rect 17405 18303 17463 18309
rect 17494 18300 17500 18352
rect 17552 18340 17558 18352
rect 17552 18312 18368 18340
rect 17552 18300 17558 18312
rect 5626 18232 5632 18284
rect 5684 18232 5690 18284
rect 6362 18232 6368 18284
rect 6420 18272 6426 18284
rect 6549 18275 6607 18281
rect 6549 18272 6561 18275
rect 6420 18244 6561 18272
rect 6420 18232 6426 18244
rect 6549 18241 6561 18244
rect 6595 18241 6607 18275
rect 6549 18235 6607 18241
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8076 18244 9444 18272
rect 8076 18232 8082 18244
rect 3881 18207 3939 18213
rect 3881 18173 3893 18207
rect 3927 18173 3939 18207
rect 3881 18167 3939 18173
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 5905 18207 5963 18213
rect 5905 18204 5917 18207
rect 4212 18176 5917 18204
rect 4212 18164 4218 18176
rect 5905 18173 5917 18176
rect 5951 18173 5963 18207
rect 5905 18167 5963 18173
rect 5920 18136 5948 18167
rect 7006 18164 7012 18216
rect 7064 18164 7070 18216
rect 8386 18164 8392 18216
rect 8444 18204 8450 18216
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 8444 18176 9321 18204
rect 8444 18164 8450 18176
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9416 18204 9444 18244
rect 9490 18232 9496 18284
rect 9548 18272 9554 18284
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 9548 18244 10793 18272
rect 9548 18232 9554 18244
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 11422 18272 11428 18284
rect 10781 18235 10839 18241
rect 10888 18244 11428 18272
rect 10888 18204 10916 18244
rect 11422 18232 11428 18244
rect 11480 18232 11486 18284
rect 12437 18275 12495 18281
rect 12437 18241 12449 18275
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18272 12587 18275
rect 12802 18272 12808 18284
rect 12575 18244 12808 18272
rect 12575 18241 12587 18244
rect 12529 18235 12587 18241
rect 9416 18176 10916 18204
rect 10965 18207 11023 18213
rect 9309 18167 9367 18173
rect 10965 18173 10977 18207
rect 11011 18204 11023 18207
rect 12452 18204 12480 18235
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 13538 18232 13544 18284
rect 13596 18272 13602 18284
rect 15473 18275 15531 18281
rect 15473 18272 15485 18275
rect 13596 18244 15485 18272
rect 13596 18232 13602 18244
rect 15473 18241 15485 18244
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 17221 18275 17279 18281
rect 17221 18241 17233 18275
rect 17267 18241 17279 18275
rect 18340 18272 18368 18312
rect 18414 18300 18420 18352
rect 18472 18340 18478 18352
rect 18598 18340 18604 18352
rect 18472 18312 18604 18340
rect 18472 18300 18478 18312
rect 18598 18300 18604 18312
rect 18656 18300 18662 18352
rect 19242 18300 19248 18352
rect 19300 18340 19306 18352
rect 19300 18312 22048 18340
rect 19300 18300 19306 18312
rect 18693 18275 18751 18281
rect 18340 18244 18552 18272
rect 17221 18235 17279 18241
rect 12713 18207 12771 18213
rect 11011 18176 12296 18204
rect 12452 18176 12572 18204
rect 11011 18173 11023 18176
rect 10965 18167 11023 18173
rect 9582 18136 9588 18148
rect 5920 18108 9588 18136
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 10413 18139 10471 18145
rect 10413 18105 10425 18139
rect 10459 18136 10471 18139
rect 12268 18136 12296 18176
rect 12544 18148 12572 18176
rect 12713 18173 12725 18207
rect 12759 18204 12771 18207
rect 13354 18204 13360 18216
rect 12759 18176 13360 18204
rect 12759 18173 12771 18176
rect 12713 18167 12771 18173
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 15749 18207 15807 18213
rect 15749 18173 15761 18207
rect 15795 18204 15807 18207
rect 16666 18204 16672 18216
rect 15795 18176 16672 18204
rect 15795 18173 15807 18176
rect 15749 18167 15807 18173
rect 16666 18164 16672 18176
rect 16724 18164 16730 18216
rect 17236 18204 17264 18235
rect 17236 18176 18276 18204
rect 12434 18136 12440 18148
rect 10459 18108 12204 18136
rect 12268 18108 12440 18136
rect 10459 18105 10471 18108
rect 10413 18099 10471 18105
rect 1578 18028 1584 18080
rect 1636 18068 1642 18080
rect 5074 18068 5080 18080
rect 1636 18040 5080 18068
rect 1636 18028 1642 18040
rect 5074 18028 5080 18040
rect 5132 18028 5138 18080
rect 5261 18071 5319 18077
rect 5261 18037 5273 18071
rect 5307 18068 5319 18071
rect 6362 18068 6368 18080
rect 5307 18040 6368 18068
rect 5307 18037 5319 18040
rect 5261 18031 5319 18037
rect 6362 18028 6368 18040
rect 6420 18028 6426 18080
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 9490 18068 9496 18080
rect 7524 18040 9496 18068
rect 7524 18028 7530 18040
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 12066 18028 12072 18080
rect 12124 18028 12130 18080
rect 12176 18068 12204 18108
rect 12434 18096 12440 18108
rect 12492 18096 12498 18148
rect 12526 18096 12532 18148
rect 12584 18136 12590 18148
rect 13265 18139 13323 18145
rect 13265 18136 13277 18139
rect 12584 18108 13277 18136
rect 12584 18096 12590 18108
rect 13265 18105 13277 18108
rect 13311 18105 13323 18139
rect 13265 18099 13323 18105
rect 14458 18096 14464 18148
rect 14516 18136 14522 18148
rect 17770 18136 17776 18148
rect 14516 18108 17776 18136
rect 14516 18096 14522 18108
rect 17770 18096 17776 18108
rect 17828 18096 17834 18148
rect 18248 18136 18276 18176
rect 18414 18164 18420 18216
rect 18472 18164 18478 18216
rect 18524 18204 18552 18244
rect 18693 18241 18705 18275
rect 18739 18272 18751 18275
rect 19794 18272 19800 18284
rect 18739 18244 19800 18272
rect 18739 18241 18751 18244
rect 18693 18235 18751 18241
rect 19794 18232 19800 18244
rect 19852 18232 19858 18284
rect 22020 18281 22048 18312
rect 22462 18300 22468 18352
rect 22520 18340 22526 18352
rect 22830 18340 22836 18352
rect 22520 18312 22836 18340
rect 22520 18300 22526 18312
rect 22830 18300 22836 18312
rect 22888 18300 22894 18352
rect 23842 18300 23848 18352
rect 23900 18300 23906 18352
rect 25038 18300 25044 18352
rect 25096 18340 25102 18352
rect 25317 18343 25375 18349
rect 25317 18340 25329 18343
rect 25096 18312 25329 18340
rect 25096 18300 25102 18312
rect 25317 18309 25329 18312
rect 25363 18309 25375 18343
rect 25317 18303 25375 18309
rect 26050 18300 26056 18352
rect 26108 18300 26114 18352
rect 28350 18340 28356 18352
rect 28092 18312 28356 18340
rect 22005 18275 22063 18281
rect 20088 18244 20300 18272
rect 20088 18204 20116 18244
rect 18524 18176 20116 18204
rect 20162 18164 20168 18216
rect 20220 18164 20226 18216
rect 20272 18213 20300 18244
rect 22005 18241 22017 18275
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 22557 18275 22615 18281
rect 22557 18241 22569 18275
rect 22603 18272 22615 18275
rect 22922 18272 22928 18284
rect 22603 18244 22928 18272
rect 22603 18241 22615 18244
rect 22557 18235 22615 18241
rect 20257 18207 20315 18213
rect 20257 18173 20269 18207
rect 20303 18173 20315 18207
rect 20257 18167 20315 18173
rect 20806 18164 20812 18216
rect 20864 18204 20870 18216
rect 21634 18204 21640 18216
rect 20864 18176 21640 18204
rect 20864 18164 20870 18176
rect 21634 18164 21640 18176
rect 21692 18204 21698 18216
rect 22572 18204 22600 18235
rect 22922 18232 22928 18244
rect 22980 18232 22986 18284
rect 24670 18232 24676 18284
rect 24728 18272 24734 18284
rect 26694 18272 26700 18284
rect 24728 18244 26700 18272
rect 24728 18232 24734 18244
rect 26694 18232 26700 18244
rect 26752 18232 26758 18284
rect 27341 18275 27399 18281
rect 27341 18241 27353 18275
rect 27387 18272 27399 18275
rect 27706 18272 27712 18284
rect 27387 18244 27712 18272
rect 27387 18241 27399 18244
rect 27341 18235 27399 18241
rect 27706 18232 27712 18244
rect 27764 18232 27770 18284
rect 27798 18232 27804 18284
rect 27856 18272 27862 18284
rect 28092 18281 28120 18312
rect 28350 18300 28356 18312
rect 28408 18300 28414 18352
rect 30653 18343 30711 18349
rect 30653 18309 30665 18343
rect 30699 18340 30711 18343
rect 30926 18340 30932 18352
rect 30699 18312 30932 18340
rect 30699 18309 30711 18312
rect 30653 18303 30711 18309
rect 30926 18300 30932 18312
rect 30984 18300 30990 18352
rect 28077 18275 28135 18281
rect 28077 18272 28089 18275
rect 27856 18244 28089 18272
rect 27856 18232 27862 18244
rect 28077 18241 28089 18244
rect 28123 18241 28135 18275
rect 28077 18235 28135 18241
rect 29454 18232 29460 18284
rect 29512 18272 29518 18284
rect 29638 18272 29644 18284
rect 29512 18244 29644 18272
rect 29512 18232 29518 18244
rect 29638 18232 29644 18244
rect 29696 18232 29702 18284
rect 21692 18176 22600 18204
rect 21692 18164 21698 18176
rect 22646 18164 22652 18216
rect 22704 18164 22710 18216
rect 23109 18207 23167 18213
rect 23109 18173 23121 18207
rect 23155 18173 23167 18207
rect 23109 18167 23167 18173
rect 23385 18207 23443 18213
rect 23385 18173 23397 18207
rect 23431 18204 23443 18207
rect 25314 18204 25320 18216
rect 23431 18176 25320 18204
rect 23431 18173 23443 18176
rect 23385 18167 23443 18173
rect 22738 18136 22744 18148
rect 18248 18108 22744 18136
rect 22738 18096 22744 18108
rect 22796 18096 22802 18148
rect 12894 18068 12900 18080
rect 12176 18040 12900 18068
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 13170 18028 13176 18080
rect 13228 18068 13234 18080
rect 21266 18068 21272 18080
rect 13228 18040 21272 18068
rect 13228 18028 13234 18040
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 21450 18028 21456 18080
rect 21508 18028 21514 18080
rect 22094 18028 22100 18080
rect 22152 18028 22158 18080
rect 23124 18068 23152 18167
rect 25314 18164 25320 18176
rect 25372 18164 25378 18216
rect 28353 18207 28411 18213
rect 28353 18173 28365 18207
rect 28399 18204 28411 18207
rect 30098 18204 30104 18216
rect 28399 18176 30104 18204
rect 28399 18173 28411 18176
rect 28353 18167 28411 18173
rect 30098 18164 30104 18176
rect 30156 18164 30162 18216
rect 30834 18164 30840 18216
rect 30892 18164 30898 18216
rect 24762 18068 24768 18080
rect 23124 18040 24768 18068
rect 24762 18028 24768 18040
rect 24820 18028 24826 18080
rect 27522 18028 27528 18080
rect 27580 18068 27586 18080
rect 29825 18071 29883 18077
rect 29825 18068 29837 18071
rect 27580 18040 29837 18068
rect 27580 18028 27586 18040
rect 29825 18037 29837 18040
rect 29871 18037 29883 18071
rect 29825 18031 29883 18037
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 1946 17864 1952 17876
rect 1728 17836 1952 17864
rect 1728 17824 1734 17836
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 4338 17824 4344 17876
rect 4396 17824 4402 17876
rect 5166 17824 5172 17876
rect 5224 17864 5230 17876
rect 6641 17867 6699 17873
rect 6641 17864 6653 17867
rect 5224 17836 6653 17864
rect 5224 17824 5230 17836
rect 6641 17833 6653 17836
rect 6687 17833 6699 17867
rect 6641 17827 6699 17833
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7285 17867 7343 17873
rect 7285 17864 7297 17867
rect 6972 17836 7297 17864
rect 6972 17824 6978 17836
rect 7285 17833 7297 17836
rect 7331 17833 7343 17867
rect 12342 17864 12348 17876
rect 7285 17827 7343 17833
rect 9646 17836 12348 17864
rect 7837 17799 7895 17805
rect 7837 17765 7849 17799
rect 7883 17796 7895 17799
rect 9646 17796 9674 17836
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 13814 17824 13820 17876
rect 13872 17864 13878 17876
rect 14461 17867 14519 17873
rect 14461 17864 14473 17867
rect 13872 17836 14473 17864
rect 13872 17824 13878 17836
rect 14461 17833 14473 17836
rect 14507 17833 14519 17867
rect 14461 17827 14519 17833
rect 15013 17867 15071 17873
rect 15013 17833 15025 17867
rect 15059 17864 15071 17867
rect 18322 17864 18328 17876
rect 15059 17836 18328 17864
rect 15059 17833 15071 17836
rect 15013 17827 15071 17833
rect 18322 17824 18328 17836
rect 18380 17824 18386 17876
rect 18414 17824 18420 17876
rect 18472 17864 18478 17876
rect 19429 17867 19487 17873
rect 19429 17864 19441 17867
rect 18472 17836 19441 17864
rect 18472 17824 18478 17836
rect 19429 17833 19441 17836
rect 19475 17833 19487 17867
rect 19429 17827 19487 17833
rect 24486 17824 24492 17876
rect 24544 17864 24550 17876
rect 26418 17864 26424 17876
rect 24544 17836 26424 17864
rect 24544 17824 24550 17836
rect 26418 17824 26424 17836
rect 26476 17824 26482 17876
rect 26602 17824 26608 17876
rect 26660 17824 26666 17876
rect 26960 17867 27018 17873
rect 26960 17833 26972 17867
rect 27006 17864 27018 17867
rect 27522 17864 27528 17876
rect 27006 17836 27528 17864
rect 27006 17833 27018 17836
rect 26960 17827 27018 17833
rect 27522 17824 27528 17836
rect 27580 17824 27586 17876
rect 27614 17824 27620 17876
rect 27672 17864 27678 17876
rect 29733 17867 29791 17873
rect 29733 17864 29745 17867
rect 27672 17836 29745 17864
rect 27672 17824 27678 17836
rect 29733 17833 29745 17836
rect 29779 17833 29791 17867
rect 29733 17827 29791 17833
rect 7883 17768 8248 17796
rect 7883 17765 7895 17768
rect 7837 17759 7895 17765
rect 1210 17688 1216 17740
rect 1268 17728 1274 17740
rect 2041 17731 2099 17737
rect 2041 17728 2053 17731
rect 1268 17700 2053 17728
rect 1268 17688 1274 17700
rect 2041 17697 2053 17700
rect 2087 17697 2099 17731
rect 2041 17691 2099 17697
rect 5810 17688 5816 17740
rect 5868 17728 5874 17740
rect 7926 17728 7932 17740
rect 5868 17700 7932 17728
rect 5868 17688 5874 17700
rect 7926 17688 7932 17700
rect 7984 17688 7990 17740
rect 8220 17728 8248 17768
rect 9048 17768 9674 17796
rect 8481 17731 8539 17737
rect 8220 17700 8340 17728
rect 1762 17620 1768 17672
rect 1820 17620 1826 17672
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4798 17660 4804 17672
rect 4212 17632 4804 17660
rect 4212 17620 4218 17632
rect 4798 17620 4804 17632
rect 4856 17660 4862 17672
rect 4893 17663 4951 17669
rect 4893 17660 4905 17663
rect 4856 17632 4905 17660
rect 4856 17620 4862 17632
rect 4893 17629 4905 17632
rect 4939 17629 4951 17663
rect 4893 17623 4951 17629
rect 6270 17620 6276 17672
rect 6328 17620 6334 17672
rect 6914 17620 6920 17672
rect 6972 17660 6978 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 6972 17632 8217 17660
rect 6972 17620 6978 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8312 17660 8340 17700
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 9048 17728 9076 17768
rect 9766 17756 9772 17808
rect 9824 17796 9830 17808
rect 10597 17799 10655 17805
rect 10597 17796 10609 17799
rect 9824 17768 10609 17796
rect 9824 17756 9830 17768
rect 10597 17765 10609 17768
rect 10643 17765 10655 17799
rect 10597 17759 10655 17765
rect 13630 17756 13636 17808
rect 13688 17796 13694 17808
rect 13725 17799 13783 17805
rect 13725 17796 13737 17799
rect 13688 17768 13737 17796
rect 13688 17756 13694 17768
rect 13725 17765 13737 17768
rect 13771 17765 13783 17799
rect 20717 17799 20775 17805
rect 20717 17796 20729 17799
rect 13725 17759 13783 17765
rect 18340 17768 20729 17796
rect 8527 17700 9076 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 9306 17688 9312 17740
rect 9364 17728 9370 17740
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 9364 17700 9873 17728
rect 9364 17688 9370 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 9950 17688 9956 17740
rect 10008 17728 10014 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10008 17700 11161 17728
rect 10008 17688 10014 17700
rect 11149 17697 11161 17700
rect 11195 17697 11207 17731
rect 11149 17691 11207 17697
rect 12253 17731 12311 17737
rect 12253 17697 12265 17731
rect 12299 17728 12311 17731
rect 13262 17728 13268 17740
rect 12299 17700 13268 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 13262 17688 13268 17700
rect 13320 17688 13326 17740
rect 16298 17688 16304 17740
rect 16356 17688 16362 17740
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 16666 17728 16672 17740
rect 16623 17700 16672 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 16666 17688 16672 17700
rect 16724 17688 16730 17740
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 18340 17728 18368 17768
rect 20717 17765 20729 17768
rect 20763 17765 20775 17799
rect 20717 17759 20775 17765
rect 17184 17700 18368 17728
rect 17184 17688 17190 17700
rect 18414 17688 18420 17740
rect 18472 17728 18478 17740
rect 21269 17731 21327 17737
rect 21269 17728 21281 17731
rect 18472 17700 21281 17728
rect 18472 17688 18478 17700
rect 21269 17697 21281 17700
rect 21315 17697 21327 17731
rect 22557 17731 22615 17737
rect 22557 17728 22569 17731
rect 21269 17691 21327 17697
rect 21376 17700 22569 17728
rect 8312 17632 9076 17660
rect 8205 17623 8263 17629
rect 4249 17595 4307 17601
rect 4249 17561 4261 17595
rect 4295 17592 4307 17595
rect 5074 17592 5080 17604
rect 4295 17564 5080 17592
rect 4295 17561 4307 17564
rect 4249 17555 4307 17561
rect 5074 17552 5080 17564
rect 5132 17552 5138 17604
rect 5169 17595 5227 17601
rect 5169 17561 5181 17595
rect 5215 17561 5227 17595
rect 5169 17555 5227 17561
rect 5184 17524 5212 17555
rect 7006 17552 7012 17604
rect 7064 17592 7070 17604
rect 7193 17595 7251 17601
rect 7193 17592 7205 17595
rect 7064 17564 7205 17592
rect 7064 17552 7070 17564
rect 7193 17561 7205 17564
rect 7239 17561 7251 17595
rect 7193 17555 7251 17561
rect 7742 17552 7748 17604
rect 7800 17592 7806 17604
rect 8846 17592 8852 17604
rect 7800 17564 8852 17592
rect 7800 17552 7806 17564
rect 8846 17552 8852 17564
rect 8904 17552 8910 17604
rect 9048 17592 9076 17632
rect 9122 17620 9128 17672
rect 9180 17620 9186 17672
rect 11974 17620 11980 17672
rect 12032 17620 12038 17672
rect 15197 17663 15255 17669
rect 15197 17629 15209 17663
rect 15243 17660 15255 17663
rect 15562 17660 15568 17672
rect 15243 17632 15568 17660
rect 15243 17629 15255 17632
rect 15197 17623 15255 17629
rect 15562 17620 15568 17632
rect 15620 17620 15626 17672
rect 15746 17620 15752 17672
rect 15804 17660 15810 17672
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15804 17632 15853 17660
rect 15804 17620 15810 17632
rect 15841 17629 15853 17632
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 17678 17620 17684 17672
rect 17736 17620 17742 17672
rect 18877 17663 18935 17669
rect 18877 17629 18889 17663
rect 18923 17660 18935 17663
rect 19242 17660 19248 17672
rect 18923 17632 19248 17660
rect 18923 17629 18935 17632
rect 18877 17623 18935 17629
rect 19242 17620 19248 17632
rect 19300 17620 19306 17672
rect 19610 17620 19616 17672
rect 19668 17620 19674 17672
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17660 20591 17663
rect 21082 17660 21088 17672
rect 20579 17632 21088 17660
rect 20579 17629 20591 17632
rect 20533 17623 20591 17629
rect 21082 17620 21088 17632
rect 21140 17620 21146 17672
rect 10226 17592 10232 17604
rect 9048 17564 10232 17592
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 10965 17595 11023 17601
rect 10965 17561 10977 17595
rect 11011 17592 11023 17595
rect 11011 17564 11744 17592
rect 11011 17561 11023 17564
rect 10965 17555 11023 17561
rect 7760 17524 7788 17552
rect 5184 17496 7788 17524
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 8297 17527 8355 17533
rect 8297 17524 8309 17527
rect 7984 17496 8309 17524
rect 7984 17484 7990 17496
rect 8297 17493 8309 17496
rect 8343 17493 8355 17527
rect 8297 17487 8355 17493
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 9732 17496 11069 17524
rect 9732 17484 9738 17496
rect 11057 17493 11069 17496
rect 11103 17493 11115 17527
rect 11716 17524 11744 17564
rect 12710 17552 12716 17604
rect 12768 17552 12774 17604
rect 14369 17595 14427 17601
rect 14369 17561 14381 17595
rect 14415 17592 14427 17595
rect 15378 17592 15384 17604
rect 14415 17564 15384 17592
rect 14415 17561 14427 17564
rect 14369 17555 14427 17561
rect 15378 17552 15384 17564
rect 15436 17552 15442 17604
rect 15930 17552 15936 17604
rect 15988 17592 15994 17604
rect 21376 17592 21404 17700
rect 22557 17697 22569 17700
rect 22603 17697 22615 17731
rect 22557 17691 22615 17697
rect 24762 17688 24768 17740
rect 24820 17728 24826 17740
rect 24857 17731 24915 17737
rect 24857 17728 24869 17731
rect 24820 17700 24869 17728
rect 24820 17688 24826 17700
rect 24857 17697 24869 17700
rect 24903 17728 24915 17731
rect 25866 17728 25872 17740
rect 24903 17700 25872 17728
rect 24903 17697 24915 17700
rect 24857 17691 24915 17697
rect 25866 17688 25872 17700
rect 25924 17728 25930 17740
rect 26697 17731 26755 17737
rect 26697 17728 26709 17731
rect 25924 17700 26709 17728
rect 25924 17688 25930 17700
rect 26697 17697 26709 17700
rect 26743 17728 26755 17731
rect 27706 17728 27712 17740
rect 26743 17700 27712 17728
rect 26743 17697 26755 17700
rect 26697 17691 26755 17697
rect 27706 17688 27712 17700
rect 27764 17688 27770 17740
rect 29454 17728 29460 17740
rect 28092 17700 29460 17728
rect 21910 17620 21916 17672
rect 21968 17660 21974 17672
rect 22281 17663 22339 17669
rect 22281 17660 22293 17663
rect 21968 17632 22293 17660
rect 21968 17620 21974 17632
rect 22281 17629 22293 17632
rect 22327 17629 22339 17663
rect 24394 17660 24400 17672
rect 23690 17632 24400 17660
rect 22281 17623 22339 17629
rect 24394 17620 24400 17632
rect 24452 17620 24458 17672
rect 28092 17646 28120 17700
rect 29454 17688 29460 17700
rect 29512 17688 29518 17740
rect 30006 17688 30012 17740
rect 30064 17728 30070 17740
rect 30285 17731 30343 17737
rect 30285 17728 30297 17731
rect 30064 17700 30297 17728
rect 30064 17688 30070 17700
rect 30285 17697 30297 17700
rect 30331 17697 30343 17731
rect 30285 17691 30343 17697
rect 28810 17620 28816 17672
rect 28868 17660 28874 17672
rect 28997 17663 29055 17669
rect 28997 17660 29009 17663
rect 28868 17632 29009 17660
rect 28868 17620 28874 17632
rect 28997 17629 29009 17632
rect 29043 17660 29055 17663
rect 30101 17663 30159 17669
rect 30101 17660 30113 17663
rect 29043 17632 30113 17660
rect 29043 17629 29055 17632
rect 28997 17623 29055 17629
rect 30101 17629 30113 17632
rect 30147 17660 30159 17663
rect 30147 17632 31754 17660
rect 30147 17629 30159 17632
rect 30101 17623 30159 17629
rect 25133 17595 25191 17601
rect 25133 17592 25145 17595
rect 15988 17564 16988 17592
rect 15988 17552 15994 17564
rect 13722 17524 13728 17536
rect 11716 17496 13728 17524
rect 11057 17487 11115 17493
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 15657 17527 15715 17533
rect 15657 17493 15669 17527
rect 15703 17524 15715 17527
rect 16206 17524 16212 17536
rect 15703 17496 16212 17524
rect 15703 17493 15715 17496
rect 15657 17487 15715 17493
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 16960 17524 16988 17564
rect 17880 17564 18736 17592
rect 17880 17524 17908 17564
rect 16960 17496 17908 17524
rect 18049 17527 18107 17533
rect 18049 17493 18061 17527
rect 18095 17524 18107 17527
rect 18414 17524 18420 17536
rect 18095 17496 18420 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 18708 17533 18736 17564
rect 18892 17564 21404 17592
rect 24044 17564 25145 17592
rect 18892 17536 18920 17564
rect 18693 17527 18751 17533
rect 18693 17493 18705 17527
rect 18739 17493 18751 17527
rect 18693 17487 18751 17493
rect 18874 17484 18880 17536
rect 18932 17484 18938 17536
rect 20162 17484 20168 17536
rect 20220 17524 20226 17536
rect 20990 17524 20996 17536
rect 20220 17496 20996 17524
rect 20220 17484 20226 17496
rect 20990 17484 20996 17496
rect 21048 17524 21054 17536
rect 21085 17527 21143 17533
rect 21085 17524 21097 17527
rect 21048 17496 21097 17524
rect 21048 17484 21054 17496
rect 21085 17493 21097 17496
rect 21131 17493 21143 17527
rect 21085 17487 21143 17493
rect 21174 17484 21180 17536
rect 21232 17484 21238 17536
rect 22462 17484 22468 17536
rect 22520 17524 22526 17536
rect 23842 17524 23848 17536
rect 22520 17496 23848 17524
rect 22520 17484 22526 17496
rect 23842 17484 23848 17496
rect 23900 17484 23906 17536
rect 24044 17533 24072 17564
rect 25133 17561 25145 17564
rect 25179 17592 25191 17595
rect 25222 17592 25228 17604
rect 25179 17564 25228 17592
rect 25179 17561 25191 17564
rect 25133 17555 25191 17561
rect 25222 17552 25228 17564
rect 25280 17552 25286 17604
rect 26418 17592 26424 17604
rect 26358 17564 26424 17592
rect 26418 17552 26424 17564
rect 26476 17552 26482 17604
rect 26694 17552 26700 17604
rect 26752 17592 26758 17604
rect 30834 17592 30840 17604
rect 26752 17564 27384 17592
rect 26752 17552 26758 17564
rect 24029 17527 24087 17533
rect 24029 17493 24041 17527
rect 24075 17493 24087 17527
rect 24029 17487 24087 17493
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 27154 17524 27160 17536
rect 24268 17496 27160 17524
rect 24268 17484 24274 17496
rect 27154 17484 27160 17496
rect 27212 17484 27218 17536
rect 27356 17524 27384 17564
rect 28966 17564 30840 17592
rect 28445 17527 28503 17533
rect 28445 17524 28457 17527
rect 27356 17496 28457 17524
rect 28445 17493 28457 17496
rect 28491 17524 28503 17527
rect 28966 17524 28994 17564
rect 30834 17552 30840 17564
rect 30892 17552 30898 17604
rect 31726 17592 31754 17632
rect 42794 17592 42800 17604
rect 31726 17564 42800 17592
rect 42794 17552 42800 17564
rect 42852 17552 42858 17604
rect 28491 17496 28994 17524
rect 28491 17493 28503 17496
rect 28445 17487 28503 17493
rect 30190 17484 30196 17536
rect 30248 17524 30254 17536
rect 30929 17527 30987 17533
rect 30929 17524 30941 17527
rect 30248 17496 30941 17524
rect 30248 17484 30254 17496
rect 30929 17493 30941 17496
rect 30975 17524 30987 17527
rect 46382 17524 46388 17536
rect 30975 17496 46388 17524
rect 30975 17493 30987 17496
rect 30929 17487 30987 17493
rect 46382 17484 46388 17496
rect 46440 17484 46446 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 6825 17323 6883 17329
rect 6825 17289 6837 17323
rect 6871 17320 6883 17323
rect 7098 17320 7104 17332
rect 6871 17292 7104 17320
rect 6871 17289 6883 17292
rect 6825 17283 6883 17289
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 7190 17280 7196 17332
rect 7248 17280 7254 17332
rect 7282 17280 7288 17332
rect 7340 17280 7346 17332
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7892 17292 8033 17320
rect 7892 17280 7898 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 8021 17283 8079 17289
rect 9490 17280 9496 17332
rect 9548 17320 9554 17332
rect 9677 17323 9735 17329
rect 9677 17320 9689 17323
rect 9548 17292 9689 17320
rect 9548 17280 9554 17292
rect 9677 17289 9689 17292
rect 9723 17320 9735 17323
rect 10781 17323 10839 17329
rect 9723 17292 10732 17320
rect 9723 17289 9735 17292
rect 9677 17283 9735 17289
rect 2314 17212 2320 17264
rect 2372 17252 2378 17264
rect 5166 17252 5172 17264
rect 2372 17224 5172 17252
rect 2372 17212 2378 17224
rect 5166 17212 5172 17224
rect 5224 17212 5230 17264
rect 5721 17255 5779 17261
rect 5721 17221 5733 17255
rect 5767 17252 5779 17255
rect 5994 17252 6000 17264
rect 5767 17224 6000 17252
rect 5767 17221 5779 17224
rect 5721 17215 5779 17221
rect 5994 17212 6000 17224
rect 6052 17212 6058 17264
rect 8478 17212 8484 17264
rect 8536 17212 8542 17264
rect 9585 17255 9643 17261
rect 9585 17221 9597 17255
rect 9631 17252 9643 17255
rect 10042 17252 10048 17264
rect 9631 17224 10048 17252
rect 9631 17221 9643 17224
rect 9585 17215 9643 17221
rect 10042 17212 10048 17224
rect 10100 17212 10106 17264
rect 10704 17252 10732 17292
rect 10781 17289 10793 17323
rect 10827 17320 10839 17323
rect 11330 17320 11336 17332
rect 10827 17292 11336 17320
rect 10827 17289 10839 17292
rect 10781 17283 10839 17289
rect 11330 17280 11336 17292
rect 11388 17280 11394 17332
rect 11882 17280 11888 17332
rect 11940 17320 11946 17332
rect 12529 17323 12587 17329
rect 12529 17320 12541 17323
rect 11940 17292 12541 17320
rect 11940 17280 11946 17292
rect 12529 17289 12541 17292
rect 12575 17289 12587 17323
rect 12529 17283 12587 17289
rect 12989 17323 13047 17329
rect 12989 17289 13001 17323
rect 13035 17320 13047 17323
rect 20162 17320 20168 17332
rect 13035 17292 20168 17320
rect 13035 17289 13047 17292
rect 12989 17283 13047 17289
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 20717 17323 20775 17329
rect 20717 17289 20729 17323
rect 20763 17289 20775 17323
rect 20717 17283 20775 17289
rect 21085 17323 21143 17329
rect 21085 17289 21097 17323
rect 21131 17320 21143 17323
rect 21450 17320 21456 17332
rect 21131 17292 21456 17320
rect 21131 17289 21143 17292
rect 21085 17283 21143 17289
rect 10704 17224 12434 17252
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 3326 17184 3332 17196
rect 1811 17156 3332 17184
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 3418 17144 3424 17196
rect 3476 17144 3482 17196
rect 5629 17187 5687 17193
rect 5629 17184 5641 17187
rect 5368 17156 5641 17184
rect 5368 17128 5396 17156
rect 5629 17153 5641 17156
rect 5675 17153 5687 17187
rect 5629 17147 5687 17153
rect 8294 17144 8300 17196
rect 8352 17184 8358 17196
rect 8389 17187 8447 17193
rect 8389 17184 8401 17187
rect 8352 17156 8401 17184
rect 8352 17144 8358 17156
rect 8389 17153 8401 17156
rect 8435 17153 8447 17187
rect 9398 17184 9404 17196
rect 8389 17147 8447 17153
rect 8496 17156 9404 17184
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1360 17088 2053 17116
rect 1360 17076 1366 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 3786 17076 3792 17128
rect 3844 17116 3850 17128
rect 3881 17119 3939 17125
rect 3881 17116 3893 17119
rect 3844 17088 3893 17116
rect 3844 17076 3850 17088
rect 3881 17085 3893 17088
rect 3927 17085 3939 17119
rect 3881 17079 3939 17085
rect 5350 17076 5356 17128
rect 5408 17076 5414 17128
rect 5902 17076 5908 17128
rect 5960 17076 5966 17128
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7469 17119 7527 17125
rect 7469 17116 7481 17119
rect 7248 17088 7481 17116
rect 7248 17076 7254 17088
rect 7469 17085 7481 17088
rect 7515 17116 7527 17119
rect 7650 17116 7656 17128
rect 7515 17088 7656 17116
rect 7515 17085 7527 17088
rect 7469 17079 7527 17085
rect 7650 17076 7656 17088
rect 7708 17116 7714 17128
rect 8496 17116 8524 17156
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10318 17184 10324 17196
rect 10008 17156 10324 17184
rect 10008 17144 10014 17156
rect 10318 17144 10324 17156
rect 10376 17184 10382 17196
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 10376 17156 11805 17184
rect 10376 17144 10382 17156
rect 11793 17153 11805 17156
rect 11839 17153 11851 17187
rect 12406 17184 12434 17224
rect 13906 17212 13912 17264
rect 13964 17252 13970 17264
rect 14737 17255 14795 17261
rect 14737 17252 14749 17255
rect 13964 17224 14749 17252
rect 13964 17212 13970 17224
rect 14737 17221 14749 17224
rect 14783 17221 14795 17255
rect 14737 17215 14795 17221
rect 17678 17212 17684 17264
rect 17736 17252 17742 17264
rect 20732 17252 20760 17283
rect 21450 17280 21456 17292
rect 21508 17280 21514 17332
rect 21542 17280 21548 17332
rect 21600 17320 21606 17332
rect 21913 17323 21971 17329
rect 21913 17320 21925 17323
rect 21600 17292 21925 17320
rect 21600 17280 21606 17292
rect 21913 17289 21925 17292
rect 21959 17289 21971 17323
rect 21913 17283 21971 17289
rect 22066 17292 22324 17320
rect 17736 17224 18906 17252
rect 19996 17224 20760 17252
rect 21177 17255 21235 17261
rect 17736 17212 17742 17224
rect 12897 17187 12955 17193
rect 12897 17184 12909 17187
rect 12406 17156 12909 17184
rect 11793 17147 11851 17153
rect 12897 17153 12909 17156
rect 12943 17153 12955 17187
rect 14645 17187 14703 17193
rect 14645 17184 14657 17187
rect 12897 17147 12955 17153
rect 13004 17156 14657 17184
rect 7708 17088 8524 17116
rect 7708 17076 7714 17088
rect 8570 17076 8576 17128
rect 8628 17076 8634 17128
rect 8754 17076 8760 17128
rect 8812 17116 8818 17128
rect 9490 17116 9496 17128
rect 8812 17088 9496 17116
rect 8812 17076 8818 17088
rect 9490 17076 9496 17088
rect 9548 17076 9554 17128
rect 9582 17076 9588 17128
rect 9640 17116 9646 17128
rect 9769 17119 9827 17125
rect 9769 17116 9781 17119
rect 9640 17088 9781 17116
rect 9640 17076 9646 17088
rect 9769 17085 9781 17088
rect 9815 17085 9827 17119
rect 9769 17079 9827 17085
rect 10870 17076 10876 17128
rect 10928 17076 10934 17128
rect 10962 17076 10968 17128
rect 11020 17076 11026 17128
rect 13004 17116 13032 17156
rect 14645 17153 14657 17156
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 16850 17144 16856 17196
rect 16908 17184 16914 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 16908 17156 17233 17184
rect 16908 17144 16914 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 12084 17088 13032 17116
rect 13173 17119 13231 17125
rect 6454 17008 6460 17060
rect 6512 17048 6518 17060
rect 11977 17051 12035 17057
rect 11977 17048 11989 17051
rect 6512 17020 11989 17048
rect 6512 17008 6518 17020
rect 11977 17017 11989 17020
rect 12023 17017 12035 17051
rect 11977 17011 12035 17017
rect 5258 16940 5264 16992
rect 5316 16940 5322 16992
rect 5626 16940 5632 16992
rect 5684 16980 5690 16992
rect 5994 16980 6000 16992
rect 5684 16952 6000 16980
rect 5684 16940 5690 16952
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 8570 16940 8576 16992
rect 8628 16980 8634 16992
rect 9217 16983 9275 16989
rect 9217 16980 9229 16983
rect 8628 16952 9229 16980
rect 8628 16940 8634 16952
rect 9217 16949 9229 16952
rect 9263 16949 9275 16983
rect 9217 16943 9275 16949
rect 9306 16940 9312 16992
rect 9364 16980 9370 16992
rect 10413 16983 10471 16989
rect 10413 16980 10425 16983
rect 9364 16952 10425 16980
rect 9364 16940 9370 16952
rect 10413 16949 10425 16952
rect 10459 16949 10471 16983
rect 10413 16943 10471 16949
rect 10686 16940 10692 16992
rect 10744 16980 10750 16992
rect 12084 16980 12112 17088
rect 13173 17085 13185 17119
rect 13219 17116 13231 17119
rect 13630 17116 13636 17128
rect 13219 17088 13636 17116
rect 13219 17085 13231 17088
rect 13173 17079 13231 17085
rect 13630 17076 13636 17088
rect 13688 17076 13694 17128
rect 14829 17119 14887 17125
rect 13740 17088 14228 17116
rect 12618 17008 12624 17060
rect 12676 17048 12682 17060
rect 13740 17048 13768 17088
rect 12676 17020 13768 17048
rect 14200 17048 14228 17088
rect 14829 17085 14841 17119
rect 14875 17085 14887 17119
rect 14829 17079 14887 17085
rect 14844 17048 14872 17079
rect 16022 17076 16028 17128
rect 16080 17116 16086 17128
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 16080 17088 17325 17116
rect 16080 17076 16086 17088
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17494 17076 17500 17128
rect 17552 17076 17558 17128
rect 18141 17119 18199 17125
rect 18141 17085 18153 17119
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 14200 17020 14872 17048
rect 12676 17008 12682 17020
rect 14918 17008 14924 17060
rect 14976 17048 14982 17060
rect 16942 17048 16948 17060
rect 14976 17020 16948 17048
rect 14976 17008 14982 17020
rect 16942 17008 16948 17020
rect 17000 17008 17006 17060
rect 17034 17008 17040 17060
rect 17092 17048 17098 17060
rect 18156 17048 18184 17079
rect 18414 17076 18420 17128
rect 18472 17076 18478 17128
rect 18874 17076 18880 17128
rect 18932 17116 18938 17128
rect 19889 17119 19947 17125
rect 19889 17116 19901 17119
rect 18932 17088 19901 17116
rect 18932 17076 18938 17088
rect 19889 17085 19901 17088
rect 19935 17085 19947 17119
rect 19889 17079 19947 17085
rect 19996 17048 20024 17224
rect 21177 17221 21189 17255
rect 21223 17252 21235 17255
rect 22066 17252 22094 17292
rect 21223 17224 22094 17252
rect 22296 17252 22324 17292
rect 22738 17280 22744 17332
rect 22796 17320 22802 17332
rect 26513 17323 26571 17329
rect 26513 17320 26525 17323
rect 22796 17292 26525 17320
rect 22796 17280 22802 17292
rect 26513 17289 26525 17292
rect 26559 17289 26571 17323
rect 30190 17320 30196 17332
rect 26513 17283 26571 17289
rect 27724 17292 30196 17320
rect 25130 17252 25136 17264
rect 22296 17224 25136 17252
rect 21223 17221 21235 17224
rect 21177 17215 21235 17221
rect 25130 17212 25136 17224
rect 25188 17212 25194 17264
rect 26418 17252 26424 17264
rect 26266 17224 26424 17252
rect 26418 17212 26424 17224
rect 26476 17252 26482 17264
rect 27154 17252 27160 17264
rect 26476 17224 27160 17252
rect 26476 17212 26482 17224
rect 27154 17212 27160 17224
rect 27212 17212 27218 17264
rect 17092 17020 18184 17048
rect 19444 17020 20024 17048
rect 20180 17156 22232 17184
rect 17092 17008 17098 17020
rect 10744 16952 12112 16980
rect 10744 16940 10750 16952
rect 14182 16940 14188 16992
rect 14240 16980 14246 16992
rect 14277 16983 14335 16989
rect 14277 16980 14289 16983
rect 14240 16952 14289 16980
rect 14240 16940 14246 16952
rect 14277 16949 14289 16952
rect 14323 16949 14335 16983
rect 14277 16943 14335 16949
rect 14826 16940 14832 16992
rect 14884 16980 14890 16992
rect 15841 16983 15899 16989
rect 15841 16980 15853 16983
rect 14884 16952 15853 16980
rect 14884 16940 14890 16952
rect 15841 16949 15853 16952
rect 15887 16949 15899 16983
rect 15841 16943 15899 16949
rect 15930 16940 15936 16992
rect 15988 16980 15994 16992
rect 16853 16983 16911 16989
rect 16853 16980 16865 16983
rect 15988 16952 16865 16980
rect 15988 16940 15994 16952
rect 16853 16949 16865 16952
rect 16899 16949 16911 16983
rect 16853 16943 16911 16949
rect 17126 16940 17132 16992
rect 17184 16980 17190 16992
rect 19444 16980 19472 17020
rect 17184 16952 19472 16980
rect 17184 16940 17190 16952
rect 19518 16940 19524 16992
rect 19576 16980 19582 16992
rect 20180 16980 20208 17156
rect 20254 17076 20260 17128
rect 20312 17116 20318 17128
rect 20312 17088 21220 17116
rect 20312 17076 20318 17088
rect 21192 17048 21220 17088
rect 21266 17076 21272 17128
rect 21324 17116 21330 17128
rect 22204 17116 22232 17156
rect 22278 17144 22284 17196
rect 22336 17144 22342 17196
rect 22373 17187 22431 17193
rect 22373 17153 22385 17187
rect 22419 17184 22431 17187
rect 22830 17184 22836 17196
rect 22419 17156 22836 17184
rect 22419 17153 22431 17156
rect 22373 17147 22431 17153
rect 22830 17144 22836 17156
rect 22888 17144 22894 17196
rect 23566 17144 23572 17196
rect 23624 17184 23630 17196
rect 23661 17187 23719 17193
rect 23661 17184 23673 17187
rect 23624 17156 23673 17184
rect 23624 17144 23630 17156
rect 23661 17153 23673 17156
rect 23707 17153 23719 17187
rect 23661 17147 23719 17153
rect 24486 17144 24492 17196
rect 24544 17144 24550 17196
rect 24762 17144 24768 17196
rect 24820 17144 24826 17196
rect 22465 17119 22523 17125
rect 22465 17116 22477 17119
rect 21324 17088 22094 17116
rect 22204 17088 22477 17116
rect 21324 17076 21330 17088
rect 22066 17048 22094 17088
rect 22465 17085 22477 17088
rect 22511 17085 22523 17119
rect 22465 17079 22523 17085
rect 23753 17119 23811 17125
rect 23753 17085 23765 17119
rect 23799 17085 23811 17119
rect 23753 17079 23811 17085
rect 22738 17048 22744 17060
rect 21192 17020 21956 17048
rect 22066 17020 22744 17048
rect 19576 16952 20208 16980
rect 21928 16980 21956 17020
rect 22738 17008 22744 17020
rect 22796 17008 22802 17060
rect 22830 17008 22836 17060
rect 22888 17048 22894 17060
rect 23293 17051 23351 17057
rect 23293 17048 23305 17051
rect 22888 17020 23305 17048
rect 22888 17008 22894 17020
rect 23293 17017 23305 17020
rect 23339 17017 23351 17051
rect 23768 17048 23796 17079
rect 23842 17076 23848 17128
rect 23900 17076 23906 17128
rect 25041 17119 25099 17125
rect 25041 17085 25053 17119
rect 25087 17116 25099 17119
rect 26694 17116 26700 17128
rect 25087 17088 26700 17116
rect 25087 17085 25099 17088
rect 25041 17079 25099 17085
rect 26694 17076 26700 17088
rect 26752 17076 26758 17128
rect 27724 17048 27752 17292
rect 30190 17280 30196 17292
rect 30248 17280 30254 17332
rect 29454 17252 29460 17264
rect 29394 17224 29460 17252
rect 29454 17212 29460 17224
rect 29512 17252 29518 17264
rect 30098 17252 30104 17264
rect 29512 17224 30104 17252
rect 29512 17212 29518 17224
rect 30098 17212 30104 17224
rect 30156 17212 30162 17264
rect 27798 17144 27804 17196
rect 27856 17184 27862 17196
rect 27893 17187 27951 17193
rect 27893 17184 27905 17187
rect 27856 17156 27905 17184
rect 27856 17144 27862 17156
rect 27893 17153 27905 17156
rect 27939 17153 27951 17187
rect 27893 17147 27951 17153
rect 28169 17119 28227 17125
rect 28169 17085 28181 17119
rect 28215 17116 28227 17119
rect 30006 17116 30012 17128
rect 28215 17088 30012 17116
rect 28215 17085 28227 17088
rect 28169 17079 28227 17085
rect 30006 17076 30012 17088
rect 30064 17076 30070 17128
rect 23293 17011 23351 17017
rect 23676 17020 23796 17048
rect 27356 17020 27752 17048
rect 23109 16983 23167 16989
rect 23109 16980 23121 16983
rect 21928 16952 23121 16980
rect 19576 16940 19582 16952
rect 23109 16949 23121 16952
rect 23155 16980 23167 16983
rect 23676 16980 23704 17020
rect 27356 16980 27384 17020
rect 23155 16952 27384 16980
rect 27433 16983 27491 16989
rect 23155 16949 23167 16952
rect 23109 16943 23167 16949
rect 27433 16949 27445 16983
rect 27479 16980 27491 16983
rect 28166 16980 28172 16992
rect 27479 16952 28172 16980
rect 27479 16949 27491 16952
rect 27433 16943 27491 16949
rect 28166 16940 28172 16952
rect 28224 16940 28230 16992
rect 28258 16940 28264 16992
rect 28316 16980 28322 16992
rect 29641 16983 29699 16989
rect 29641 16980 29653 16983
rect 28316 16952 29653 16980
rect 28316 16940 28322 16952
rect 29641 16949 29653 16952
rect 29687 16949 29699 16983
rect 29641 16943 29699 16949
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 8110 16776 8116 16788
rect 2746 16748 8116 16776
rect 2222 16600 2228 16652
rect 2280 16640 2286 16652
rect 2746 16640 2774 16748
rect 8110 16736 8116 16748
rect 8168 16776 8174 16788
rect 8168 16748 11652 16776
rect 8168 16736 8174 16748
rect 10045 16711 10103 16717
rect 10045 16708 10057 16711
rect 4172 16680 10057 16708
rect 4172 16640 4200 16680
rect 10045 16677 10057 16680
rect 10091 16677 10103 16711
rect 10045 16671 10103 16677
rect 10137 16711 10195 16717
rect 10137 16677 10149 16711
rect 10183 16708 10195 16711
rect 10226 16708 10232 16720
rect 10183 16680 10232 16708
rect 10183 16677 10195 16680
rect 10137 16671 10195 16677
rect 10226 16668 10232 16680
rect 10284 16668 10290 16720
rect 10318 16668 10324 16720
rect 10376 16708 10382 16720
rect 10870 16708 10876 16720
rect 10376 16680 10876 16708
rect 10376 16668 10382 16680
rect 10870 16668 10876 16680
rect 10928 16668 10934 16720
rect 2280 16612 2774 16640
rect 3988 16612 4200 16640
rect 2280 16600 2286 16612
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 3988 16572 4016 16612
rect 5258 16600 5264 16652
rect 5316 16640 5322 16652
rect 7101 16643 7159 16649
rect 7101 16640 7113 16643
rect 5316 16612 7113 16640
rect 5316 16600 5322 16612
rect 7101 16609 7113 16612
rect 7147 16609 7159 16643
rect 7101 16603 7159 16609
rect 7190 16600 7196 16652
rect 7248 16600 7254 16652
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 7300 16612 8401 16640
rect 1811 16544 4016 16572
rect 4065 16575 4123 16581
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 4065 16541 4077 16575
rect 4111 16572 4123 16575
rect 6089 16575 6147 16581
rect 6089 16572 6101 16575
rect 4111 16544 5120 16572
rect 4111 16541 4123 16544
rect 4065 16535 4123 16541
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 2501 16467 2559 16473
rect 3970 16464 3976 16516
rect 4028 16504 4034 16516
rect 4893 16507 4951 16513
rect 4893 16504 4905 16507
rect 4028 16476 4905 16504
rect 4028 16464 4034 16476
rect 4893 16473 4905 16476
rect 4939 16473 4951 16507
rect 4893 16467 4951 16473
rect 5092 16436 5120 16544
rect 5644 16544 6101 16572
rect 5166 16464 5172 16516
rect 5224 16504 5230 16516
rect 5644 16504 5672 16544
rect 6089 16541 6101 16544
rect 6135 16541 6147 16575
rect 6089 16535 6147 16541
rect 6546 16532 6552 16584
rect 6604 16572 6610 16584
rect 7300 16572 7328 16612
rect 8389 16609 8401 16612
rect 8435 16640 8447 16643
rect 10689 16643 10747 16649
rect 10689 16640 10701 16643
rect 8435 16612 10701 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 10689 16609 10701 16612
rect 10735 16640 10747 16643
rect 10962 16640 10968 16652
rect 10735 16612 10968 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 10962 16600 10968 16612
rect 11020 16640 11026 16652
rect 11514 16640 11520 16652
rect 11020 16612 11520 16640
rect 11020 16600 11026 16612
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 11624 16640 11652 16748
rect 12342 16736 12348 16788
rect 12400 16776 12406 16788
rect 15930 16776 15936 16788
rect 12400 16748 15936 16776
rect 12400 16736 12406 16748
rect 15930 16736 15936 16748
rect 15988 16736 15994 16788
rect 16850 16736 16856 16788
rect 16908 16736 16914 16788
rect 16942 16736 16948 16788
rect 17000 16776 17006 16788
rect 17000 16748 18736 16776
rect 17000 16736 17006 16748
rect 12989 16711 13047 16717
rect 12989 16677 13001 16711
rect 13035 16677 13047 16711
rect 18414 16708 18420 16720
rect 12989 16671 13047 16677
rect 13648 16680 18420 16708
rect 12253 16643 12311 16649
rect 12253 16640 12265 16643
rect 11624 16612 12265 16640
rect 12253 16609 12265 16612
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 12434 16600 12440 16652
rect 12492 16600 12498 16652
rect 6604 16544 7328 16572
rect 6604 16532 6610 16544
rect 8202 16532 8208 16584
rect 8260 16532 8266 16584
rect 9677 16575 9735 16581
rect 9677 16541 9689 16575
rect 9723 16572 9735 16575
rect 9766 16572 9772 16584
rect 9723 16544 9772 16572
rect 9723 16541 9735 16544
rect 9677 16535 9735 16541
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 9861 16575 9919 16581
rect 9861 16541 9873 16575
rect 9907 16572 9919 16575
rect 10134 16572 10140 16584
rect 9907 16544 10140 16572
rect 9907 16541 9919 16544
rect 9861 16535 9919 16541
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 10594 16532 10600 16584
rect 10652 16532 10658 16584
rect 12066 16572 12072 16584
rect 11164 16544 12072 16572
rect 11164 16516 11192 16544
rect 12066 16532 12072 16544
rect 12124 16532 12130 16584
rect 13004 16572 13032 16671
rect 13446 16600 13452 16652
rect 13504 16600 13510 16652
rect 13648 16649 13676 16680
rect 18414 16668 18420 16680
rect 18472 16668 18478 16720
rect 18708 16708 18736 16748
rect 18782 16736 18788 16788
rect 18840 16736 18846 16788
rect 18874 16736 18880 16788
rect 18932 16776 18938 16788
rect 19426 16776 19432 16788
rect 18932 16748 19432 16776
rect 18932 16736 18938 16748
rect 19426 16736 19432 16748
rect 19484 16736 19490 16788
rect 20254 16776 20260 16788
rect 19536 16748 20260 16776
rect 19536 16708 19564 16748
rect 20254 16736 20260 16748
rect 20312 16736 20318 16788
rect 21174 16736 21180 16788
rect 21232 16776 21238 16788
rect 25774 16776 25780 16788
rect 21232 16748 25780 16776
rect 21232 16736 21238 16748
rect 25774 16736 25780 16748
rect 25832 16736 25838 16788
rect 18708 16680 19564 16708
rect 20806 16668 20812 16720
rect 20864 16708 20870 16720
rect 21542 16708 21548 16720
rect 20864 16680 21548 16708
rect 20864 16668 20870 16680
rect 21542 16668 21548 16680
rect 21600 16668 21606 16720
rect 22649 16711 22707 16717
rect 22649 16677 22661 16711
rect 22695 16708 22707 16711
rect 22922 16708 22928 16720
rect 22695 16680 22928 16708
rect 22695 16677 22707 16680
rect 22649 16671 22707 16677
rect 22922 16668 22928 16680
rect 22980 16708 22986 16720
rect 23382 16708 23388 16720
rect 22980 16680 23388 16708
rect 22980 16668 22986 16680
rect 23382 16668 23388 16680
rect 23440 16668 23446 16720
rect 25222 16668 25228 16720
rect 25280 16708 25286 16720
rect 25280 16680 28488 16708
rect 25280 16668 25286 16680
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16609 13691 16643
rect 13633 16603 13691 16609
rect 14553 16643 14611 16649
rect 14553 16609 14565 16643
rect 14599 16640 14611 16643
rect 15378 16640 15384 16652
rect 14599 16612 15384 16640
rect 14599 16609 14611 16612
rect 14553 16603 14611 16609
rect 15378 16600 15384 16612
rect 15436 16600 15442 16652
rect 15657 16643 15715 16649
rect 15657 16609 15669 16643
rect 15703 16640 15715 16643
rect 15838 16640 15844 16652
rect 15703 16612 15844 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 21266 16640 21272 16652
rect 19751 16612 21272 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 22738 16600 22744 16652
rect 22796 16640 22802 16652
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 22796 16612 23765 16640
rect 22796 16600 22802 16612
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 25130 16600 25136 16652
rect 25188 16600 25194 16652
rect 25317 16643 25375 16649
rect 25317 16609 25329 16643
rect 25363 16640 25375 16643
rect 25682 16640 25688 16652
rect 25363 16612 25688 16640
rect 25363 16609 25375 16612
rect 25317 16603 25375 16609
rect 25682 16600 25688 16612
rect 25740 16600 25746 16652
rect 27062 16600 27068 16652
rect 27120 16600 27126 16652
rect 27246 16600 27252 16652
rect 27304 16640 27310 16652
rect 28258 16640 28264 16652
rect 27304 16612 28264 16640
rect 27304 16600 27310 16612
rect 28258 16600 28264 16612
rect 28316 16600 28322 16652
rect 28460 16649 28488 16680
rect 28445 16643 28503 16649
rect 28445 16609 28457 16643
rect 28491 16640 28503 16643
rect 31570 16640 31576 16652
rect 28491 16612 31576 16640
rect 28491 16609 28503 16612
rect 28445 16603 28503 16609
rect 31570 16600 31576 16612
rect 31628 16600 31634 16652
rect 16758 16572 16764 16584
rect 13004 16544 16764 16572
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16572 17555 16575
rect 17862 16572 17868 16584
rect 17543 16544 17868 16572
rect 17543 16541 17555 16544
rect 17497 16535 17555 16541
rect 17862 16532 17868 16544
rect 17920 16532 17926 16584
rect 18141 16575 18199 16581
rect 18141 16541 18153 16575
rect 18187 16572 18199 16575
rect 18414 16572 18420 16584
rect 18187 16544 18420 16572
rect 18187 16541 18199 16544
rect 18141 16535 18199 16541
rect 18414 16532 18420 16544
rect 18472 16532 18478 16584
rect 19426 16532 19432 16584
rect 19484 16532 19490 16584
rect 23474 16532 23480 16584
rect 23532 16572 23538 16584
rect 23569 16575 23627 16581
rect 23569 16572 23581 16575
rect 23532 16544 23581 16572
rect 23532 16532 23538 16544
rect 23569 16541 23581 16544
rect 23615 16541 23627 16575
rect 23569 16535 23627 16541
rect 24118 16532 24124 16584
rect 24176 16572 24182 16584
rect 26973 16575 27031 16581
rect 24176 16544 25452 16572
rect 24176 16532 24182 16544
rect 5224 16476 5672 16504
rect 5905 16507 5963 16513
rect 5224 16464 5230 16476
rect 5905 16473 5917 16507
rect 5951 16504 5963 16507
rect 5994 16504 6000 16516
rect 5951 16476 6000 16504
rect 5951 16473 5963 16476
rect 5905 16467 5963 16473
rect 5994 16464 6000 16476
rect 6052 16464 6058 16516
rect 7374 16504 7380 16516
rect 6656 16476 7380 16504
rect 6454 16436 6460 16448
rect 5092 16408 6460 16436
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 6656 16445 6684 16476
rect 7374 16464 7380 16476
rect 7432 16464 7438 16516
rect 8110 16464 8116 16516
rect 8168 16504 8174 16516
rect 8297 16507 8355 16513
rect 8297 16504 8309 16507
rect 8168 16476 8309 16504
rect 8168 16464 8174 16476
rect 8297 16473 8309 16476
rect 8343 16473 8355 16507
rect 8297 16467 8355 16473
rect 8478 16464 8484 16516
rect 8536 16504 8542 16516
rect 10226 16504 10232 16516
rect 8536 16476 10232 16504
rect 8536 16464 8542 16476
rect 10226 16464 10232 16476
rect 10284 16464 10290 16516
rect 11146 16464 11152 16516
rect 11204 16464 11210 16516
rect 13538 16504 13544 16516
rect 11808 16476 13544 16504
rect 6641 16439 6699 16445
rect 6641 16405 6653 16439
rect 6687 16405 6699 16439
rect 6641 16399 6699 16405
rect 7006 16396 7012 16448
rect 7064 16396 7070 16448
rect 7834 16396 7840 16448
rect 7892 16396 7898 16448
rect 9398 16396 9404 16448
rect 9456 16436 9462 16448
rect 10134 16436 10140 16448
rect 9456 16408 10140 16436
rect 9456 16396 9462 16408
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 10502 16396 10508 16448
rect 10560 16396 10566 16448
rect 11808 16445 11836 16476
rect 13538 16464 13544 16476
rect 13596 16464 13602 16516
rect 19334 16504 19340 16516
rect 15028 16476 19340 16504
rect 11793 16439 11851 16445
rect 11793 16405 11805 16439
rect 11839 16405 11851 16439
rect 11793 16399 11851 16405
rect 11882 16396 11888 16448
rect 11940 16436 11946 16448
rect 12161 16439 12219 16445
rect 12161 16436 12173 16439
rect 11940 16408 12173 16436
rect 11940 16396 11946 16408
rect 12161 16405 12173 16408
rect 12207 16405 12219 16439
rect 12161 16399 12219 16405
rect 13262 16396 13268 16448
rect 13320 16436 13326 16448
rect 15028 16445 15056 16476
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 20990 16504 20996 16516
rect 20930 16476 20996 16504
rect 20990 16464 20996 16476
rect 21048 16464 21054 16516
rect 21450 16464 21456 16516
rect 21508 16464 21514 16516
rect 22066 16476 23244 16504
rect 13357 16439 13415 16445
rect 13357 16436 13369 16439
rect 13320 16408 13369 16436
rect 13320 16396 13326 16408
rect 13357 16405 13369 16408
rect 13403 16405 13415 16439
rect 13357 16399 13415 16405
rect 15013 16439 15071 16445
rect 15013 16405 15025 16439
rect 15059 16405 15071 16439
rect 15013 16399 15071 16405
rect 15378 16396 15384 16448
rect 15436 16396 15442 16448
rect 15470 16396 15476 16448
rect 15528 16396 15534 16448
rect 15654 16396 15660 16448
rect 15712 16436 15718 16448
rect 17313 16439 17371 16445
rect 17313 16436 17325 16439
rect 15712 16408 17325 16436
rect 15712 16396 15718 16408
rect 17313 16405 17325 16408
rect 17359 16405 17371 16439
rect 17313 16399 17371 16405
rect 17957 16439 18015 16445
rect 17957 16405 17969 16439
rect 18003 16436 18015 16439
rect 19150 16436 19156 16448
rect 18003 16408 19156 16436
rect 18003 16405 18015 16408
rect 17957 16399 18015 16405
rect 19150 16396 19156 16408
rect 19208 16396 19214 16448
rect 20714 16396 20720 16448
rect 20772 16436 20778 16448
rect 22066 16436 22094 16476
rect 23216 16445 23244 16476
rect 23382 16464 23388 16516
rect 23440 16504 23446 16516
rect 25041 16507 25099 16513
rect 23440 16476 24716 16504
rect 23440 16464 23446 16476
rect 20772 16408 22094 16436
rect 23201 16439 23259 16445
rect 20772 16396 20778 16408
rect 23201 16405 23213 16439
rect 23247 16405 23259 16439
rect 23201 16399 23259 16405
rect 23661 16439 23719 16445
rect 23661 16405 23673 16439
rect 23707 16436 23719 16439
rect 23750 16436 23756 16448
rect 23707 16408 23756 16436
rect 23707 16405 23719 16408
rect 23661 16399 23719 16405
rect 23750 16396 23756 16408
rect 23808 16436 23814 16448
rect 24210 16436 24216 16448
rect 23808 16408 24216 16436
rect 23808 16396 23814 16408
rect 24210 16396 24216 16408
rect 24268 16396 24274 16448
rect 24688 16445 24716 16476
rect 25041 16473 25053 16507
rect 25087 16504 25099 16507
rect 25222 16504 25228 16516
rect 25087 16476 25228 16504
rect 25087 16473 25099 16476
rect 25041 16467 25099 16473
rect 25222 16464 25228 16476
rect 25280 16464 25286 16516
rect 24673 16439 24731 16445
rect 24673 16405 24685 16439
rect 24719 16405 24731 16439
rect 25424 16436 25452 16544
rect 26973 16541 26985 16575
rect 27019 16572 27031 16575
rect 27614 16572 27620 16584
rect 27019 16544 27620 16572
rect 27019 16541 27031 16544
rect 26973 16535 27031 16541
rect 27614 16532 27620 16544
rect 27672 16532 27678 16584
rect 28166 16532 28172 16584
rect 28224 16532 28230 16584
rect 25498 16464 25504 16516
rect 25556 16504 25562 16516
rect 25556 16476 27844 16504
rect 25556 16464 25562 16476
rect 27816 16445 27844 16476
rect 27890 16464 27896 16516
rect 27948 16504 27954 16516
rect 28261 16507 28319 16513
rect 28261 16504 28273 16507
rect 27948 16476 28273 16504
rect 27948 16464 27954 16476
rect 28261 16473 28273 16476
rect 28307 16504 28319 16507
rect 28442 16504 28448 16516
rect 28307 16476 28448 16504
rect 28307 16473 28319 16476
rect 28261 16467 28319 16473
rect 28442 16464 28448 16476
rect 28500 16464 28506 16516
rect 26605 16439 26663 16445
rect 26605 16436 26617 16439
rect 25424 16408 26617 16436
rect 24673 16399 24731 16405
rect 26605 16405 26617 16408
rect 26651 16405 26663 16439
rect 26605 16399 26663 16405
rect 27801 16439 27859 16445
rect 27801 16405 27813 16439
rect 27847 16405 27859 16439
rect 27801 16399 27859 16405
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 5629 16235 5687 16241
rect 5629 16201 5641 16235
rect 5675 16232 5687 16235
rect 6086 16232 6092 16244
rect 5675 16204 6092 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 6086 16192 6092 16204
rect 6144 16192 6150 16244
rect 7285 16235 7343 16241
rect 7285 16201 7297 16235
rect 7331 16232 7343 16235
rect 7558 16232 7564 16244
rect 7331 16204 7564 16232
rect 7331 16201 7343 16204
rect 7285 16195 7343 16201
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 7742 16192 7748 16244
rect 7800 16232 7806 16244
rect 7926 16232 7932 16244
rect 7800 16204 7932 16232
rect 7800 16192 7806 16204
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 12710 16232 12716 16244
rect 10060 16204 12716 16232
rect 10060 16176 10088 16204
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 13354 16192 13360 16244
rect 13412 16232 13418 16244
rect 13817 16235 13875 16241
rect 13817 16232 13829 16235
rect 13412 16204 13829 16232
rect 13412 16192 13418 16204
rect 13817 16201 13829 16204
rect 13863 16201 13875 16235
rect 13817 16195 13875 16201
rect 14826 16192 14832 16244
rect 14884 16192 14890 16244
rect 15378 16192 15384 16244
rect 15436 16232 15442 16244
rect 17773 16235 17831 16241
rect 17773 16232 17785 16235
rect 15436 16204 17785 16232
rect 15436 16192 15442 16204
rect 17773 16201 17785 16204
rect 17819 16201 17831 16235
rect 17773 16195 17831 16201
rect 17865 16235 17923 16241
rect 17865 16201 17877 16235
rect 17911 16232 17923 16235
rect 20806 16232 20812 16244
rect 17911 16204 20812 16232
rect 17911 16201 17923 16204
rect 17865 16195 17923 16201
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 21082 16192 21088 16244
rect 21140 16192 21146 16244
rect 22186 16192 22192 16244
rect 22244 16192 22250 16244
rect 22646 16192 22652 16244
rect 22704 16232 22710 16244
rect 22833 16235 22891 16241
rect 22833 16232 22845 16235
rect 22704 16204 22845 16232
rect 22704 16192 22710 16204
rect 22833 16201 22845 16204
rect 22879 16232 22891 16235
rect 22922 16232 22928 16244
rect 22879 16204 22928 16232
rect 22879 16201 22891 16204
rect 22833 16195 22891 16201
rect 22922 16192 22928 16204
rect 22980 16232 22986 16244
rect 23661 16235 23719 16241
rect 23661 16232 23673 16235
rect 22980 16204 23673 16232
rect 22980 16192 22986 16204
rect 23661 16201 23673 16204
rect 23707 16201 23719 16235
rect 23661 16195 23719 16201
rect 23750 16192 23756 16244
rect 23808 16192 23814 16244
rect 24946 16192 24952 16244
rect 25004 16232 25010 16244
rect 26605 16235 26663 16241
rect 26605 16232 26617 16235
rect 25004 16204 26617 16232
rect 25004 16192 25010 16204
rect 26605 16201 26617 16204
rect 26651 16201 26663 16235
rect 26605 16195 26663 16201
rect 4338 16124 4344 16176
rect 4396 16124 4402 16176
rect 6825 16167 6883 16173
rect 5644 16136 6776 16164
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 3605 16099 3663 16105
rect 1811 16068 2774 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2746 16028 2774 16068
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 5644 16096 5672 16136
rect 3651 16068 5672 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 6454 16096 6460 16108
rect 5776 16068 6460 16096
rect 5776 16056 5782 16068
rect 6454 16056 6460 16068
rect 6512 16056 6518 16108
rect 6641 16099 6699 16105
rect 6641 16065 6653 16099
rect 6687 16065 6699 16099
rect 6641 16059 6699 16065
rect 4798 16028 4804 16040
rect 2746 16000 4804 16028
rect 2041 15991 2099 15997
rect 4798 15988 4804 16000
rect 4856 15988 4862 16040
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 16028 5963 16031
rect 6546 16028 6552 16040
rect 5951 16000 6552 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 6546 15988 6552 16000
rect 6604 15988 6610 16040
rect 5261 15895 5319 15901
rect 5261 15861 5273 15895
rect 5307 15892 5319 15895
rect 6546 15892 6552 15904
rect 5307 15864 6552 15892
rect 5307 15861 5319 15864
rect 5261 15855 5319 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 6656 15892 6684 16059
rect 6748 15960 6776 16136
rect 6825 16133 6837 16167
rect 6871 16164 6883 16167
rect 8662 16164 8668 16176
rect 6871 16136 8668 16164
rect 6871 16133 6883 16136
rect 6825 16127 6883 16133
rect 8662 16124 8668 16136
rect 8720 16124 8726 16176
rect 8757 16167 8815 16173
rect 8757 16133 8769 16167
rect 8803 16164 8815 16167
rect 8846 16164 8852 16176
rect 8803 16136 8852 16164
rect 8803 16133 8815 16136
rect 8757 16127 8815 16133
rect 8846 16124 8852 16136
rect 8904 16124 8910 16176
rect 10042 16164 10048 16176
rect 9982 16136 10048 16164
rect 10042 16124 10048 16136
rect 10100 16124 10106 16176
rect 12618 16164 12624 16176
rect 10152 16136 12624 16164
rect 7650 16056 7656 16108
rect 7708 16056 7714 16108
rect 7926 16096 7932 16108
rect 7852 16068 7932 16096
rect 7742 15988 7748 16040
rect 7800 15988 7806 16040
rect 7852 16037 7880 16068
rect 7926 16056 7932 16068
rect 7984 16056 7990 16108
rect 8386 16056 8392 16108
rect 8444 16096 8450 16108
rect 8481 16099 8539 16105
rect 8481 16096 8493 16099
rect 8444 16068 8493 16096
rect 8444 16056 8450 16068
rect 8481 16065 8493 16068
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 7837 16031 7895 16037
rect 7837 15997 7849 16031
rect 7883 15997 7895 16031
rect 7837 15991 7895 15997
rect 8018 15988 8024 16040
rect 8076 16028 8082 16040
rect 10152 16028 10180 16136
rect 12618 16124 12624 16136
rect 12676 16124 12682 16176
rect 12728 16164 12756 16192
rect 21450 16164 21456 16176
rect 12728 16136 12834 16164
rect 13832 16136 21456 16164
rect 11146 16056 11152 16108
rect 11204 16056 11210 16108
rect 11974 16056 11980 16108
rect 12032 16096 12038 16108
rect 12069 16099 12127 16105
rect 12069 16096 12081 16099
rect 12032 16068 12081 16096
rect 12032 16056 12038 16068
rect 12069 16065 12081 16068
rect 12115 16065 12127 16099
rect 12069 16059 12127 16065
rect 8076 16000 10180 16028
rect 8076 15988 8082 16000
rect 10226 15988 10232 16040
rect 10284 16028 10290 16040
rect 10410 16028 10416 16040
rect 10284 16000 10416 16028
rect 10284 15988 10290 16000
rect 10410 15988 10416 16000
rect 10468 15988 10474 16040
rect 12345 16031 12403 16037
rect 12345 15997 12357 16031
rect 12391 16028 12403 16031
rect 13538 16028 13544 16040
rect 12391 16000 13544 16028
rect 12391 15997 12403 16000
rect 12345 15991 12403 15997
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 7926 15960 7932 15972
rect 6748 15932 7932 15960
rect 7926 15920 7932 15932
rect 7984 15920 7990 15972
rect 10502 15960 10508 15972
rect 10152 15932 10508 15960
rect 10152 15892 10180 15932
rect 10502 15920 10508 15932
rect 10560 15920 10566 15972
rect 6656 15864 10180 15892
rect 10594 15852 10600 15904
rect 10652 15892 10658 15904
rect 10965 15895 11023 15901
rect 10965 15892 10977 15895
rect 10652 15864 10977 15892
rect 10652 15852 10658 15864
rect 10965 15861 10977 15864
rect 11011 15861 11023 15895
rect 10965 15855 11023 15861
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 12158 15892 12164 15904
rect 11572 15864 12164 15892
rect 11572 15852 11578 15864
rect 12158 15852 12164 15864
rect 12216 15892 12222 15904
rect 13832 15892 13860 16136
rect 21450 16124 21456 16136
rect 21508 16124 21514 16176
rect 27154 16164 27160 16176
rect 26358 16136 27160 16164
rect 27154 16124 27160 16136
rect 27212 16124 27218 16176
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16065 16359 16099
rect 16301 16059 16359 16065
rect 14458 15988 14464 16040
rect 14516 16028 14522 16040
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 14516 16000 14933 16028
rect 14516 15988 14522 16000
rect 14921 15997 14933 16000
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 15010 15988 15016 16040
rect 15068 15988 15074 16040
rect 16316 15960 16344 16059
rect 18506 16056 18512 16108
rect 18564 16096 18570 16108
rect 18785 16099 18843 16105
rect 18785 16096 18797 16099
rect 18564 16068 18797 16096
rect 18564 16056 18570 16068
rect 18785 16065 18797 16068
rect 18831 16065 18843 16099
rect 18785 16059 18843 16065
rect 18966 16056 18972 16108
rect 19024 16096 19030 16108
rect 19153 16099 19211 16105
rect 19153 16096 19165 16099
rect 19024 16068 19165 16096
rect 19024 16056 19030 16068
rect 19153 16065 19165 16068
rect 19199 16065 19211 16099
rect 19153 16059 19211 16065
rect 20162 16056 20168 16108
rect 20220 16096 20226 16108
rect 21177 16099 21235 16105
rect 21177 16096 21189 16099
rect 20220 16068 21189 16096
rect 20220 16056 20226 16068
rect 21177 16065 21189 16068
rect 21223 16065 21235 16099
rect 21177 16059 21235 16065
rect 23768 16068 24348 16096
rect 17402 15988 17408 16040
rect 17460 16028 17466 16040
rect 17957 16031 18015 16037
rect 17957 16028 17969 16031
rect 17460 16000 17969 16028
rect 17460 15988 17466 16000
rect 17957 15997 17969 16000
rect 18003 15997 18015 16031
rect 17957 15991 18015 15997
rect 18322 15988 18328 16040
rect 18380 16028 18386 16040
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 18380 16000 18889 16028
rect 18380 15988 18386 16000
rect 18877 15997 18889 16000
rect 18923 15997 18935 16031
rect 18877 15991 18935 15997
rect 21361 16031 21419 16037
rect 21361 15997 21373 16031
rect 21407 16028 21419 16031
rect 23768 16028 23796 16068
rect 21407 16000 23796 16028
rect 21407 15997 21419 16000
rect 21361 15991 21419 15997
rect 23842 15988 23848 16040
rect 23900 15988 23906 16040
rect 24320 16028 24348 16068
rect 24854 16056 24860 16108
rect 24912 16056 24918 16108
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24320 16000 25145 16028
rect 25133 15997 25145 16000
rect 25179 16028 25191 16031
rect 27246 16028 27252 16040
rect 25179 16000 27252 16028
rect 25179 15997 25191 16000
rect 25133 15991 25191 15997
rect 27246 15988 27252 16000
rect 27304 15988 27310 16040
rect 16316 15932 17816 15960
rect 12216 15864 13860 15892
rect 12216 15852 12222 15864
rect 13906 15852 13912 15904
rect 13964 15892 13970 15904
rect 14461 15895 14519 15901
rect 14461 15892 14473 15895
rect 13964 15864 14473 15892
rect 13964 15852 13970 15864
rect 14461 15861 14473 15864
rect 14507 15861 14519 15895
rect 14461 15855 14519 15861
rect 16114 15852 16120 15904
rect 16172 15852 16178 15904
rect 16666 15852 16672 15904
rect 16724 15892 16730 15904
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 16724 15864 17417 15892
rect 16724 15852 16730 15864
rect 17405 15861 17417 15864
rect 17451 15861 17463 15895
rect 17788 15892 17816 15932
rect 17862 15920 17868 15972
rect 17920 15960 17926 15972
rect 17920 15932 22094 15960
rect 17920 15920 17926 15932
rect 20622 15892 20628 15904
rect 17788 15864 20628 15892
rect 17405 15855 17463 15861
rect 20622 15852 20628 15864
rect 20680 15852 20686 15904
rect 20717 15895 20775 15901
rect 20717 15861 20729 15895
rect 20763 15892 20775 15895
rect 21358 15892 21364 15904
rect 20763 15864 21364 15892
rect 20763 15861 20775 15864
rect 20717 15855 20775 15861
rect 21358 15852 21364 15864
rect 21416 15852 21422 15904
rect 22066 15892 22094 15932
rect 22554 15920 22560 15972
rect 22612 15960 22618 15972
rect 23293 15963 23351 15969
rect 23293 15960 23305 15963
rect 22612 15932 23305 15960
rect 22612 15920 22618 15932
rect 23293 15929 23305 15932
rect 23339 15929 23351 15963
rect 23293 15923 23351 15929
rect 24670 15892 24676 15904
rect 22066 15864 24676 15892
rect 24670 15852 24676 15864
rect 24728 15852 24734 15904
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 3973 15691 4031 15697
rect 3973 15657 3985 15691
rect 4019 15688 4031 15691
rect 4019 15660 6960 15688
rect 4019 15657 4031 15660
rect 3973 15651 4031 15657
rect 6932 15620 6960 15660
rect 7006 15648 7012 15700
rect 7064 15688 7070 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7064 15660 7849 15688
rect 7064 15648 7070 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 7926 15648 7932 15700
rect 7984 15688 7990 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 7984 15660 9321 15688
rect 7984 15648 7990 15660
rect 9309 15657 9321 15660
rect 9355 15657 9367 15691
rect 9309 15651 9367 15657
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 10686 15688 10692 15700
rect 9548 15660 10692 15688
rect 9548 15648 9554 15660
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 10778 15648 10784 15700
rect 10836 15688 10842 15700
rect 10836 15660 11008 15688
rect 10836 15648 10842 15660
rect 8662 15620 8668 15632
rect 6932 15592 8668 15620
rect 8662 15580 8668 15592
rect 8720 15580 8726 15632
rect 10226 15580 10232 15632
rect 10284 15580 10290 15632
rect 10870 15580 10876 15632
rect 10928 15580 10934 15632
rect 10980 15620 11008 15660
rect 12066 15648 12072 15700
rect 12124 15648 12130 15700
rect 12250 15648 12256 15700
rect 12308 15688 12314 15700
rect 16114 15688 16120 15700
rect 12308 15660 16120 15688
rect 12308 15648 12314 15660
rect 16114 15648 16120 15660
rect 16172 15648 16178 15700
rect 19429 15691 19487 15697
rect 19429 15657 19441 15691
rect 19475 15688 19487 15691
rect 19518 15688 19524 15700
rect 19475 15660 19524 15688
rect 19475 15657 19487 15660
rect 19429 15651 19487 15657
rect 19518 15648 19524 15660
rect 19576 15648 19582 15700
rect 19978 15648 19984 15700
rect 20036 15688 20042 15700
rect 20036 15660 23152 15688
rect 20036 15648 20042 15660
rect 13541 15623 13599 15629
rect 13541 15620 13553 15623
rect 10980 15592 13553 15620
rect 13541 15589 13553 15592
rect 13587 15589 13599 15623
rect 13541 15583 13599 15589
rect 14737 15623 14795 15629
rect 14737 15589 14749 15623
rect 14783 15620 14795 15623
rect 15470 15620 15476 15632
rect 14783 15592 15476 15620
rect 14783 15589 14795 15592
rect 14737 15583 14795 15589
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 15933 15623 15991 15629
rect 15933 15589 15945 15623
rect 15979 15620 15991 15623
rect 16022 15620 16028 15632
rect 15979 15592 16028 15620
rect 15979 15589 15991 15592
rect 15933 15583 15991 15589
rect 16022 15580 16028 15592
rect 16080 15580 16086 15632
rect 22186 15580 22192 15632
rect 22244 15620 22250 15632
rect 23017 15623 23075 15629
rect 23017 15620 23029 15623
rect 22244 15592 23029 15620
rect 22244 15580 22250 15592
rect 23017 15589 23029 15592
rect 23063 15589 23075 15623
rect 23017 15583 23075 15589
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 1360 15524 2053 15552
rect 1360 15512 1366 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 4430 15512 4436 15564
rect 4488 15512 4494 15564
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15552 4675 15555
rect 4706 15552 4712 15564
rect 4663 15524 4712 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 5721 15555 5779 15561
rect 5721 15552 5733 15555
rect 5592 15524 5733 15552
rect 5592 15512 5598 15524
rect 5721 15521 5733 15524
rect 5767 15552 5779 15555
rect 6730 15552 6736 15564
rect 5767 15524 6736 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 6730 15512 6736 15524
rect 6788 15512 6794 15564
rect 7006 15512 7012 15564
rect 7064 15512 7070 15564
rect 7374 15512 7380 15564
rect 7432 15552 7438 15564
rect 8018 15552 8024 15564
rect 7432 15524 8024 15552
rect 7432 15512 7438 15524
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 8481 15555 8539 15561
rect 8481 15521 8493 15555
rect 8527 15552 8539 15555
rect 8846 15552 8852 15564
rect 8527 15524 8852 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 8846 15512 8852 15524
rect 8904 15552 8910 15564
rect 8904 15524 9674 15552
rect 8904 15512 8910 15524
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 2498 15484 2504 15496
rect 1811 15456 2504 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 6362 15444 6368 15496
rect 6420 15484 6426 15496
rect 6420 15456 6776 15484
rect 6420 15444 6426 15456
rect 5629 15419 5687 15425
rect 5629 15385 5641 15419
rect 5675 15416 5687 15419
rect 5810 15416 5816 15428
rect 5675 15388 5816 15416
rect 5675 15385 5687 15388
rect 5629 15379 5687 15385
rect 5810 15376 5816 15388
rect 5868 15416 5874 15428
rect 6086 15416 6092 15428
rect 5868 15388 6092 15416
rect 5868 15376 5874 15388
rect 6086 15376 6092 15388
rect 6144 15376 6150 15428
rect 6638 15416 6644 15428
rect 6288 15388 6644 15416
rect 4062 15308 4068 15360
rect 4120 15348 4126 15360
rect 4341 15351 4399 15357
rect 4341 15348 4353 15351
rect 4120 15320 4353 15348
rect 4120 15308 4126 15320
rect 4341 15317 4353 15320
rect 4387 15317 4399 15351
rect 4341 15311 4399 15317
rect 5166 15308 5172 15360
rect 5224 15308 5230 15360
rect 5537 15351 5595 15357
rect 5537 15317 5549 15351
rect 5583 15348 5595 15351
rect 6288 15348 6316 15388
rect 6638 15376 6644 15388
rect 6696 15376 6702 15428
rect 6748 15416 6776 15456
rect 7190 15444 7196 15496
rect 7248 15484 7254 15496
rect 8297 15487 8355 15493
rect 8297 15484 8309 15487
rect 7248 15456 8309 15484
rect 7248 15444 7254 15456
rect 8297 15453 8309 15456
rect 8343 15453 8355 15487
rect 8297 15447 8355 15453
rect 9030 15444 9036 15496
rect 9088 15484 9094 15496
rect 9646 15484 9674 15524
rect 11422 15512 11428 15564
rect 11480 15512 11486 15564
rect 12710 15512 12716 15564
rect 12768 15512 12774 15564
rect 14918 15512 14924 15564
rect 14976 15552 14982 15564
rect 15289 15555 15347 15561
rect 15289 15552 15301 15555
rect 14976 15524 15301 15552
rect 14976 15512 14982 15524
rect 15289 15521 15301 15524
rect 15335 15521 15347 15555
rect 15289 15515 15347 15521
rect 16393 15555 16451 15561
rect 16393 15521 16405 15555
rect 16439 15552 16451 15555
rect 16482 15552 16488 15564
rect 16439 15524 16488 15552
rect 16439 15521 16451 15524
rect 16393 15515 16451 15521
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 16577 15555 16635 15561
rect 16577 15521 16589 15555
rect 16623 15552 16635 15555
rect 17405 15555 17463 15561
rect 17405 15552 17417 15555
rect 16623 15524 17417 15552
rect 16623 15521 16635 15524
rect 16577 15515 16635 15521
rect 17405 15521 17417 15524
rect 17451 15552 17463 15555
rect 18414 15552 18420 15564
rect 17451 15524 18420 15552
rect 17451 15521 17463 15524
rect 17405 15515 17463 15521
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 19426 15512 19432 15564
rect 19484 15552 19490 15564
rect 19705 15555 19763 15561
rect 19705 15552 19717 15555
rect 19484 15524 19717 15552
rect 19484 15512 19490 15524
rect 19705 15521 19717 15524
rect 19751 15552 19763 15555
rect 20622 15552 20628 15564
rect 19751 15524 20628 15552
rect 19751 15521 19763 15524
rect 19705 15515 19763 15521
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 22094 15512 22100 15564
rect 22152 15552 22158 15564
rect 22465 15555 22523 15561
rect 22465 15552 22477 15555
rect 22152 15524 22477 15552
rect 22152 15512 22158 15524
rect 22465 15521 22477 15524
rect 22511 15521 22523 15555
rect 22465 15515 22523 15521
rect 22649 15555 22707 15561
rect 22649 15521 22661 15555
rect 22695 15552 22707 15555
rect 23124 15552 23152 15660
rect 23750 15552 23756 15564
rect 22695 15524 23756 15552
rect 22695 15521 22707 15524
rect 22649 15515 22707 15521
rect 23750 15512 23756 15524
rect 23808 15512 23814 15564
rect 25682 15512 25688 15564
rect 25740 15552 25746 15564
rect 25777 15555 25835 15561
rect 25777 15552 25789 15555
rect 25740 15524 25789 15552
rect 25740 15512 25746 15524
rect 25777 15521 25789 15524
rect 25823 15521 25835 15555
rect 25777 15515 25835 15521
rect 10226 15484 10232 15496
rect 9088 15456 9352 15484
rect 9646 15456 10232 15484
rect 9088 15444 9094 15456
rect 6825 15419 6883 15425
rect 6825 15416 6837 15419
rect 6748 15388 6837 15416
rect 6825 15385 6837 15388
rect 6871 15385 6883 15419
rect 8570 15416 8576 15428
rect 6825 15379 6883 15385
rect 6932 15388 8576 15416
rect 5583 15320 6316 15348
rect 5583 15317 5595 15320
rect 5537 15311 5595 15317
rect 6362 15308 6368 15360
rect 6420 15308 6426 15360
rect 6733 15351 6791 15357
rect 6733 15317 6745 15351
rect 6779 15348 6791 15351
rect 6932 15348 6960 15388
rect 8570 15376 8576 15388
rect 8628 15376 8634 15428
rect 9214 15376 9220 15428
rect 9272 15376 9278 15428
rect 9324 15416 9352 15456
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 10413 15487 10471 15493
rect 10413 15453 10425 15487
rect 10459 15484 10471 15487
rect 10962 15484 10968 15496
rect 10459 15456 10968 15484
rect 10459 15453 10471 15456
rect 10413 15447 10471 15453
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 11241 15487 11299 15493
rect 11241 15484 11253 15487
rect 11204 15456 11253 15484
rect 11204 15444 11210 15456
rect 11241 15453 11253 15456
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 12066 15444 12072 15496
rect 12124 15484 12130 15496
rect 12529 15487 12587 15493
rect 12529 15484 12541 15487
rect 12124 15456 12541 15484
rect 12124 15444 12130 15456
rect 12529 15453 12541 15456
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 16942 15484 16948 15496
rect 13771 15456 16948 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 17034 15444 17040 15496
rect 17092 15484 17098 15496
rect 17129 15487 17187 15493
rect 17129 15484 17141 15487
rect 17092 15456 17141 15484
rect 17092 15444 17098 15456
rect 17129 15453 17141 15456
rect 17175 15453 17187 15487
rect 17129 15447 17187 15453
rect 19334 15444 19340 15496
rect 19392 15484 19398 15496
rect 19613 15487 19671 15493
rect 19613 15484 19625 15487
rect 19392 15456 19625 15484
rect 19392 15444 19398 15456
rect 19613 15453 19625 15456
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 20990 15444 20996 15496
rect 21048 15484 21054 15496
rect 22002 15484 22008 15496
rect 21048 15456 22008 15484
rect 21048 15444 21054 15456
rect 22002 15444 22008 15456
rect 22060 15444 22066 15496
rect 22373 15487 22431 15493
rect 22373 15453 22385 15487
rect 22419 15484 22431 15487
rect 22830 15484 22836 15496
rect 22419 15456 22836 15484
rect 22419 15453 22431 15456
rect 22373 15447 22431 15453
rect 22830 15444 22836 15456
rect 22888 15444 22894 15496
rect 23109 15487 23167 15493
rect 23109 15453 23121 15487
rect 23155 15484 23167 15487
rect 24578 15484 24584 15496
rect 23155 15456 24584 15484
rect 23155 15453 23167 15456
rect 23109 15447 23167 15453
rect 10778 15416 10784 15428
rect 9324 15388 10784 15416
rect 10778 15376 10784 15388
rect 10836 15376 10842 15428
rect 11330 15376 11336 15428
rect 11388 15376 11394 15428
rect 15194 15376 15200 15428
rect 15252 15376 15258 15428
rect 17678 15376 17684 15428
rect 17736 15416 17742 15428
rect 17736 15388 17894 15416
rect 17736 15376 17742 15388
rect 19978 15376 19984 15428
rect 20036 15376 20042 15428
rect 23124 15416 23152 15447
rect 24578 15444 24584 15456
rect 24636 15484 24642 15496
rect 25038 15484 25044 15496
rect 24636 15456 25044 15484
rect 24636 15444 24642 15456
rect 25038 15444 25044 15456
rect 25096 15444 25102 15496
rect 25406 15444 25412 15496
rect 25464 15484 25470 15496
rect 25593 15487 25651 15493
rect 25593 15484 25605 15487
rect 25464 15456 25605 15484
rect 25464 15444 25470 15456
rect 25593 15453 25605 15456
rect 25639 15484 25651 15487
rect 26142 15484 26148 15496
rect 25639 15456 26148 15484
rect 25639 15453 25651 15456
rect 25593 15447 25651 15453
rect 26142 15444 26148 15456
rect 26200 15444 26206 15496
rect 21284 15388 23152 15416
rect 6779 15320 6960 15348
rect 6779 15317 6791 15320
rect 6733 15311 6791 15317
rect 8202 15308 8208 15360
rect 8260 15348 8266 15360
rect 12250 15348 12256 15360
rect 8260 15320 12256 15348
rect 8260 15308 8266 15320
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 12434 15308 12440 15360
rect 12492 15308 12498 15360
rect 14734 15308 14740 15360
rect 14792 15348 14798 15360
rect 15105 15351 15163 15357
rect 15105 15348 15117 15351
rect 14792 15320 15117 15348
rect 14792 15308 14798 15320
rect 15105 15317 15117 15320
rect 15151 15317 15163 15351
rect 15105 15311 15163 15317
rect 16298 15308 16304 15360
rect 16356 15308 16362 15360
rect 17218 15308 17224 15360
rect 17276 15348 17282 15360
rect 17494 15348 17500 15360
rect 17276 15320 17500 15348
rect 17276 15308 17282 15320
rect 17494 15308 17500 15320
rect 17552 15348 17558 15360
rect 18877 15351 18935 15357
rect 18877 15348 18889 15351
rect 17552 15320 18889 15348
rect 17552 15308 17558 15320
rect 18877 15317 18889 15320
rect 18923 15317 18935 15351
rect 18877 15311 18935 15317
rect 19702 15308 19708 15360
rect 19760 15348 19766 15360
rect 21284 15348 21312 15388
rect 23934 15376 23940 15428
rect 23992 15376 23998 15428
rect 24854 15376 24860 15428
rect 24912 15416 24918 15428
rect 25424 15416 25452 15444
rect 24912 15388 25452 15416
rect 25685 15419 25743 15425
rect 24912 15376 24918 15388
rect 25685 15385 25697 15419
rect 25731 15416 25743 15419
rect 25774 15416 25780 15428
rect 25731 15388 25780 15416
rect 25731 15385 25743 15388
rect 25685 15379 25743 15385
rect 25774 15376 25780 15388
rect 25832 15376 25838 15428
rect 19760 15320 21312 15348
rect 19760 15308 19766 15320
rect 21450 15308 21456 15360
rect 21508 15308 21514 15360
rect 21542 15308 21548 15360
rect 21600 15348 21606 15360
rect 22005 15351 22063 15357
rect 22005 15348 22017 15351
rect 21600 15320 22017 15348
rect 21600 15308 21606 15320
rect 22005 15317 22017 15320
rect 22051 15317 22063 15351
rect 22005 15311 22063 15317
rect 22094 15308 22100 15360
rect 22152 15348 22158 15360
rect 23566 15348 23572 15360
rect 22152 15320 23572 15348
rect 22152 15308 22158 15320
rect 23566 15308 23572 15320
rect 23624 15308 23630 15360
rect 24118 15308 24124 15360
rect 24176 15348 24182 15360
rect 25225 15351 25283 15357
rect 25225 15348 25237 15351
rect 24176 15320 25237 15348
rect 24176 15308 24182 15320
rect 25225 15317 25237 15320
rect 25271 15317 25283 15351
rect 25225 15311 25283 15317
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 4798 15104 4804 15156
rect 4856 15144 4862 15156
rect 6733 15147 6791 15153
rect 6733 15144 6745 15147
rect 4856 15116 6745 15144
rect 4856 15104 4862 15116
rect 6733 15113 6745 15116
rect 6779 15113 6791 15147
rect 6733 15107 6791 15113
rect 7745 15147 7803 15153
rect 7745 15113 7757 15147
rect 7791 15144 7803 15147
rect 8570 15144 8576 15156
rect 7791 15116 8576 15144
rect 7791 15113 7803 15116
rect 7745 15107 7803 15113
rect 4433 15079 4491 15085
rect 4433 15045 4445 15079
rect 4479 15076 4491 15079
rect 4706 15076 4712 15088
rect 4479 15048 4712 15076
rect 4479 15045 4491 15048
rect 4433 15039 4491 15045
rect 4706 15036 4712 15048
rect 4764 15036 4770 15088
rect 5994 15036 6000 15088
rect 6052 15076 6058 15088
rect 7760 15076 7788 15107
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 8846 15104 8852 15156
rect 8904 15144 8910 15156
rect 9217 15147 9275 15153
rect 9217 15144 9229 15147
rect 8904 15116 9229 15144
rect 8904 15104 8910 15116
rect 9217 15113 9229 15116
rect 9263 15113 9275 15147
rect 9217 15107 9275 15113
rect 9398 15104 9404 15156
rect 9456 15144 9462 15156
rect 11882 15144 11888 15156
rect 9456 15116 11888 15144
rect 9456 15104 9462 15116
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12860 15116 13001 15144
rect 12860 15104 12866 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 13872 15116 16160 15144
rect 13872 15104 13878 15116
rect 6052 15048 7788 15076
rect 6052 15036 6058 15048
rect 7834 15036 7840 15088
rect 7892 15076 7898 15088
rect 7892 15048 8294 15076
rect 7892 15036 7898 15048
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 1854 15008 1860 15020
rect 1811 14980 1860 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 4154 14968 4160 15020
rect 4212 14968 4218 15020
rect 6270 15008 6276 15020
rect 5566 14980 6276 15008
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 6638 14968 6644 15020
rect 6696 14968 6702 15020
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 6788 14980 7972 15008
rect 6788 14968 6794 14980
rect 7944 14952 7972 14980
rect 1302 14900 1308 14952
rect 1360 14940 1366 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 1360 14912 2053 14940
rect 1360 14900 1366 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 2314 14900 2320 14952
rect 2372 14940 2378 14952
rect 3602 14940 3608 14952
rect 2372 14912 3608 14940
rect 2372 14900 2378 14912
rect 3602 14900 3608 14912
rect 3660 14900 3666 14952
rect 7742 14940 7748 14952
rect 4264 14912 7748 14940
rect 1486 14832 1492 14884
rect 1544 14872 1550 14884
rect 4264 14872 4292 14912
rect 7742 14900 7748 14912
rect 7800 14940 7806 14952
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 7800 14912 7849 14940
rect 7800 14900 7806 14912
rect 7837 14909 7849 14912
rect 7883 14909 7895 14943
rect 7837 14903 7895 14909
rect 7926 14900 7932 14952
rect 7984 14900 7990 14952
rect 1544 14844 4292 14872
rect 1544 14832 1550 14844
rect 5810 14832 5816 14884
rect 5868 14872 5874 14884
rect 5905 14875 5963 14881
rect 5905 14872 5917 14875
rect 5868 14844 5917 14872
rect 5868 14832 5874 14844
rect 5905 14841 5917 14844
rect 5951 14872 5963 14875
rect 7098 14872 7104 14884
rect 5951 14844 7104 14872
rect 5951 14841 5963 14844
rect 5905 14835 5963 14841
rect 7098 14832 7104 14844
rect 7156 14832 7162 14884
rect 7558 14872 7564 14884
rect 7208 14844 7564 14872
rect 3697 14807 3755 14813
rect 3697 14773 3709 14807
rect 3743 14804 3755 14807
rect 7208 14804 7236 14844
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 8266 14872 8294 15048
rect 9306 15036 9312 15088
rect 9364 15076 9370 15088
rect 9364 15048 9444 15076
rect 9364 15036 9370 15048
rect 9416 15008 9444 15048
rect 10778 15036 10784 15088
rect 10836 15036 10842 15088
rect 10873 15079 10931 15085
rect 10873 15045 10885 15079
rect 10919 15076 10931 15079
rect 10919 15048 11100 15076
rect 10919 15045 10931 15048
rect 10873 15039 10931 15045
rect 9585 15011 9643 15017
rect 9585 15008 9597 15011
rect 9416 14980 9597 15008
rect 9585 14977 9597 14980
rect 9631 14977 9643 15011
rect 11072 15008 11100 15048
rect 11514 15036 11520 15088
rect 11572 15076 11578 15088
rect 13357 15079 13415 15085
rect 13357 15076 13369 15079
rect 11572 15048 13369 15076
rect 11572 15036 11578 15048
rect 13357 15045 13369 15048
rect 13403 15045 13415 15079
rect 13357 15039 13415 15045
rect 15102 15036 15108 15088
rect 15160 15076 15166 15088
rect 16132 15076 16160 15116
rect 16942 15104 16948 15156
rect 17000 15144 17006 15156
rect 19429 15147 19487 15153
rect 19429 15144 19441 15147
rect 17000 15116 19441 15144
rect 17000 15104 17006 15116
rect 19429 15113 19441 15116
rect 19475 15113 19487 15147
rect 19429 15107 19487 15113
rect 20622 15104 20628 15156
rect 20680 15144 20686 15156
rect 21910 15144 21916 15156
rect 20680 15116 21916 15144
rect 20680 15104 20686 15116
rect 21910 15104 21916 15116
rect 21968 15144 21974 15156
rect 22278 15144 22284 15156
rect 21968 15116 22284 15144
rect 21968 15104 21974 15116
rect 19797 15079 19855 15085
rect 19797 15076 19809 15079
rect 15160 15048 15318 15076
rect 16132 15048 19809 15076
rect 15160 15036 15166 15048
rect 19797 15045 19809 15048
rect 19843 15045 19855 15079
rect 19797 15039 19855 15045
rect 19889 15079 19947 15085
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 21542 15076 21548 15088
rect 19935 15048 21548 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 21542 15036 21548 15048
rect 21600 15036 21606 15088
rect 11422 15008 11428 15020
rect 11072 14980 11428 15008
rect 9585 14971 9643 14977
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 11974 14968 11980 15020
rect 12032 14968 12038 15020
rect 17126 14968 17132 15020
rect 17184 14968 17190 15020
rect 20625 15011 20683 15017
rect 20625 15008 20637 15011
rect 19904 14980 20637 15008
rect 8757 14943 8815 14949
rect 8757 14909 8769 14943
rect 8803 14940 8815 14943
rect 9490 14940 9496 14952
rect 8803 14912 9496 14940
rect 8803 14909 8815 14912
rect 8757 14903 8815 14909
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 9677 14943 9735 14949
rect 9677 14940 9689 14943
rect 9600 14912 9689 14940
rect 9600 14872 9628 14912
rect 9677 14909 9689 14912
rect 9723 14909 9735 14943
rect 9677 14903 9735 14909
rect 9766 14900 9772 14952
rect 9824 14900 9830 14952
rect 10965 14943 11023 14949
rect 10965 14909 10977 14943
rect 11011 14909 11023 14943
rect 10965 14903 11023 14909
rect 11701 14943 11759 14949
rect 11701 14909 11713 14943
rect 11747 14940 11759 14943
rect 12342 14940 12348 14952
rect 11747 14912 12348 14940
rect 11747 14909 11759 14912
rect 11701 14903 11759 14909
rect 8266 14844 9628 14872
rect 10410 14832 10416 14884
rect 10468 14832 10474 14884
rect 3743 14776 7236 14804
rect 3743 14773 3755 14776
rect 3697 14767 3755 14773
rect 7282 14764 7288 14816
rect 7340 14804 7346 14816
rect 7377 14807 7435 14813
rect 7377 14804 7389 14807
rect 7340 14776 7389 14804
rect 7340 14764 7346 14776
rect 7377 14773 7389 14776
rect 7423 14773 7435 14807
rect 7377 14767 7435 14773
rect 7926 14764 7932 14816
rect 7984 14804 7990 14816
rect 10980 14804 11008 14903
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 13446 14900 13452 14952
rect 13504 14900 13510 14952
rect 13538 14900 13544 14952
rect 13596 14900 13602 14952
rect 14550 14900 14556 14952
rect 14608 14900 14614 14952
rect 14829 14943 14887 14949
rect 14829 14909 14841 14943
rect 14875 14940 14887 14943
rect 14918 14940 14924 14952
rect 14875 14912 14924 14940
rect 14875 14909 14887 14912
rect 14829 14903 14887 14909
rect 14918 14900 14924 14912
rect 14976 14940 14982 14952
rect 15286 14940 15292 14952
rect 14976 14912 15292 14940
rect 14976 14900 14982 14912
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 15838 14940 15844 14952
rect 15528 14912 15844 14940
rect 15528 14900 15534 14912
rect 15838 14900 15844 14912
rect 15896 14940 15902 14952
rect 16301 14943 16359 14949
rect 16301 14940 16313 14943
rect 15896 14912 16313 14940
rect 15896 14900 15902 14912
rect 16301 14909 16313 14912
rect 16347 14909 16359 14943
rect 16301 14903 16359 14909
rect 18874 14900 18880 14952
rect 18932 14900 18938 14952
rect 19058 14900 19064 14952
rect 19116 14940 19122 14952
rect 19904 14940 19932 14980
rect 20625 14977 20637 14980
rect 20671 14977 20683 15011
rect 20625 14971 20683 14977
rect 20898 14968 20904 15020
rect 20956 14968 20962 15020
rect 22020 15017 22048 15116
rect 22278 15104 22284 15116
rect 22336 15144 22342 15156
rect 23934 15144 23940 15156
rect 22336 15116 23940 15144
rect 22336 15104 22342 15116
rect 23934 15104 23940 15116
rect 23992 15104 23998 15156
rect 24946 15104 24952 15156
rect 25004 15104 25010 15156
rect 23566 15076 23572 15088
rect 23506 15048 23572 15076
rect 23566 15036 23572 15048
rect 23624 15076 23630 15088
rect 24394 15076 24400 15088
rect 23624 15048 24400 15076
rect 23624 15036 23630 15048
rect 24394 15036 24400 15048
rect 24452 15036 24458 15088
rect 24964 15076 24992 15104
rect 25133 15079 25191 15085
rect 25133 15076 25145 15079
rect 24964 15048 25145 15076
rect 25133 15045 25145 15048
rect 25179 15045 25191 15079
rect 27154 15076 27160 15088
rect 26358 15048 27160 15076
rect 25133 15039 25191 15045
rect 27154 15036 27160 15048
rect 27212 15036 27218 15088
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 23934 14968 23940 15020
rect 23992 15008 23998 15020
rect 24857 15011 24915 15017
rect 24857 15008 24869 15011
rect 23992 14980 24869 15008
rect 23992 14968 23998 14980
rect 24857 14977 24869 14980
rect 24903 14977 24915 15011
rect 24857 14971 24915 14977
rect 19116 14912 19932 14940
rect 20073 14943 20131 14949
rect 19116 14900 19122 14912
rect 20073 14909 20085 14943
rect 20119 14909 20131 14943
rect 20073 14903 20131 14909
rect 20088 14872 20116 14903
rect 23750 14900 23756 14952
rect 23808 14900 23814 14952
rect 21450 14872 21456 14884
rect 20088 14844 21456 14872
rect 21450 14832 21456 14844
rect 21508 14832 21514 14884
rect 7984 14776 11008 14804
rect 7984 14764 7990 14776
rect 11606 14764 11612 14816
rect 11664 14804 11670 14816
rect 16114 14804 16120 14816
rect 11664 14776 16120 14804
rect 11664 14764 11670 14776
rect 16114 14764 16120 14776
rect 16172 14764 16178 14816
rect 22268 14807 22326 14813
rect 22268 14773 22280 14807
rect 22314 14804 22326 14807
rect 22462 14804 22468 14816
rect 22314 14776 22468 14804
rect 22314 14773 22326 14776
rect 22268 14767 22326 14773
rect 22462 14764 22468 14776
rect 22520 14764 22526 14816
rect 26602 14764 26608 14816
rect 26660 14764 26666 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 3973 14603 4031 14609
rect 3973 14569 3985 14603
rect 4019 14600 4031 14603
rect 4062 14600 4068 14612
rect 4019 14572 4068 14600
rect 4019 14569 4031 14572
rect 3973 14563 4031 14569
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 9401 14603 9459 14609
rect 9401 14569 9413 14603
rect 9447 14600 9459 14603
rect 9447 14572 9904 14600
rect 9447 14569 9459 14572
rect 9401 14563 9459 14569
rect 9876 14544 9904 14572
rect 12250 14560 12256 14612
rect 12308 14600 12314 14612
rect 14734 14600 14740 14612
rect 12308 14572 14740 14600
rect 12308 14560 12314 14572
rect 14734 14560 14740 14572
rect 14792 14560 14798 14612
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 18601 14603 18659 14609
rect 18601 14600 18613 14603
rect 15344 14572 18613 14600
rect 15344 14560 15350 14572
rect 18601 14569 18613 14572
rect 18647 14569 18659 14603
rect 22922 14600 22928 14612
rect 18601 14563 18659 14569
rect 21192 14572 22928 14600
rect 6638 14492 6644 14544
rect 6696 14532 6702 14544
rect 6696 14504 9720 14532
rect 6696 14492 6702 14504
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1360 14436 2053 14464
rect 1360 14424 1366 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14464 4583 14467
rect 5534 14464 5540 14476
rect 4571 14436 5540 14464
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 5626 14424 5632 14476
rect 5684 14464 5690 14476
rect 5994 14464 6000 14476
rect 5684 14436 6000 14464
rect 5684 14424 5690 14436
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6546 14424 6552 14476
rect 6604 14464 6610 14476
rect 8389 14467 8447 14473
rect 6604 14436 8248 14464
rect 6604 14424 6610 14436
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 2866 14396 2872 14408
rect 1811 14368 2872 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 4062 14356 4068 14408
rect 4120 14396 4126 14408
rect 4614 14396 4620 14408
rect 4120 14368 4620 14396
rect 4120 14356 4126 14368
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 5261 14399 5319 14405
rect 5261 14396 5273 14399
rect 4856 14368 5273 14396
rect 4856 14356 4862 14368
rect 5261 14365 5273 14368
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 7285 14399 7343 14405
rect 7285 14365 7297 14399
rect 7331 14396 7343 14399
rect 7374 14396 7380 14408
rect 7331 14368 7380 14396
rect 7331 14365 7343 14368
rect 7285 14359 7343 14365
rect 7374 14356 7380 14368
rect 7432 14396 7438 14408
rect 7558 14396 7564 14408
rect 7432 14368 7564 14396
rect 7432 14356 7438 14368
rect 7558 14356 7564 14368
rect 7616 14356 7622 14408
rect 8220 14405 8248 14436
rect 8389 14433 8401 14467
rect 8435 14464 8447 14467
rect 9490 14464 9496 14476
rect 8435 14436 9496 14464
rect 8435 14433 8447 14436
rect 8389 14427 8447 14433
rect 9490 14424 9496 14436
rect 9548 14424 9554 14476
rect 9692 14464 9720 14504
rect 9858 14492 9864 14544
rect 9916 14492 9922 14544
rect 10502 14532 10508 14544
rect 9968 14504 10508 14532
rect 9968 14464 9996 14504
rect 10502 14492 10508 14504
rect 10560 14532 10566 14544
rect 11054 14532 11060 14544
rect 10560 14504 11060 14532
rect 10560 14492 10566 14504
rect 11054 14492 11060 14504
rect 11112 14492 11118 14544
rect 13538 14492 13544 14544
rect 13596 14532 13602 14544
rect 13725 14535 13783 14541
rect 13725 14532 13737 14535
rect 13596 14504 13737 14532
rect 13596 14492 13602 14504
rect 13725 14501 13737 14504
rect 13771 14501 13783 14535
rect 13725 14495 13783 14501
rect 18782 14492 18788 14544
rect 18840 14532 18846 14544
rect 19058 14532 19064 14544
rect 18840 14504 19064 14532
rect 18840 14492 18846 14504
rect 19058 14492 19064 14504
rect 19116 14532 19122 14544
rect 21192 14532 21220 14572
rect 22922 14560 22928 14572
rect 22980 14560 22986 14612
rect 19116 14504 21220 14532
rect 19116 14492 19122 14504
rect 9692 14436 9996 14464
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 10134 14464 10140 14476
rect 10091 14436 10140 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 10318 14424 10324 14476
rect 10376 14464 10382 14476
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 10376 14436 11161 14464
rect 10376 14424 10382 14436
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 11149 14427 11207 14433
rect 12253 14467 12311 14473
rect 12253 14433 12265 14467
rect 12299 14464 12311 14467
rect 12710 14464 12716 14476
rect 12299 14436 12716 14464
rect 12299 14433 12311 14436
rect 12253 14427 12311 14433
rect 12710 14424 12716 14436
rect 12768 14464 12774 14476
rect 13446 14464 13452 14476
rect 12768 14436 13452 14464
rect 12768 14424 12774 14436
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 15470 14464 15476 14476
rect 14967 14436 15476 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 16114 14424 16120 14476
rect 16172 14464 16178 14476
rect 19705 14467 19763 14473
rect 19705 14464 19717 14467
rect 16172 14436 19717 14464
rect 16172 14424 16178 14436
rect 19705 14433 19717 14436
rect 19751 14433 19763 14467
rect 19705 14427 19763 14433
rect 8205 14399 8263 14405
rect 8205 14365 8217 14399
rect 8251 14365 8263 14399
rect 8205 14359 8263 14365
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 8478 14396 8484 14408
rect 8343 14368 8484 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 9030 14356 9036 14408
rect 9088 14396 9094 14408
rect 9398 14396 9404 14408
rect 9088 14368 9404 14396
rect 9088 14356 9094 14368
rect 9398 14356 9404 14368
rect 9456 14396 9462 14408
rect 9766 14396 9772 14408
rect 9456 14368 9772 14396
rect 9456 14356 9462 14368
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14396 9919 14399
rect 10870 14396 10876 14408
rect 9907 14368 10876 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11790 14396 11796 14408
rect 11011 14368 11796 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 11974 14356 11980 14408
rect 12032 14356 12038 14408
rect 14642 14356 14648 14408
rect 14700 14356 14706 14408
rect 16853 14399 16911 14405
rect 16853 14365 16865 14399
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14396 19487 14399
rect 20806 14396 20812 14408
rect 19475 14368 20812 14396
rect 19475 14365 19487 14368
rect 19429 14359 19487 14365
rect 4154 14288 4160 14340
rect 4212 14328 4218 14340
rect 4433 14331 4491 14337
rect 4433 14328 4445 14331
rect 4212 14300 4445 14328
rect 4212 14288 4218 14300
rect 4433 14297 4445 14300
rect 4479 14328 4491 14331
rect 4890 14328 4896 14340
rect 4479 14300 4896 14328
rect 4479 14297 4491 14300
rect 4433 14291 4491 14297
rect 4890 14288 4896 14300
rect 4948 14288 4954 14340
rect 6270 14288 6276 14340
rect 6328 14288 6334 14340
rect 7392 14300 12388 14328
rect 4338 14220 4344 14272
rect 4396 14220 4402 14272
rect 4522 14220 4528 14272
rect 4580 14260 4586 14272
rect 7392 14260 7420 14300
rect 4580 14232 7420 14260
rect 4580 14220 4586 14232
rect 7834 14220 7840 14272
rect 7892 14220 7898 14272
rect 9769 14263 9827 14269
rect 9769 14229 9781 14263
rect 9815 14260 9827 14263
rect 9858 14260 9864 14272
rect 9815 14232 9864 14260
rect 9815 14229 9827 14232
rect 9769 14223 9827 14229
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 10134 14220 10140 14272
rect 10192 14260 10198 14272
rect 10597 14263 10655 14269
rect 10597 14260 10609 14263
rect 10192 14232 10609 14260
rect 10192 14220 10198 14232
rect 10597 14229 10609 14232
rect 10643 14229 10655 14263
rect 10597 14223 10655 14229
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 10744 14232 11069 14260
rect 10744 14220 10750 14232
rect 11057 14229 11069 14232
rect 11103 14260 11115 14263
rect 12250 14260 12256 14272
rect 11103 14232 12256 14260
rect 11103 14229 11115 14232
rect 11057 14223 11115 14229
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 12360 14260 12388 14300
rect 12710 14288 12716 14340
rect 12768 14288 12774 14340
rect 16868 14328 16896 14359
rect 20806 14356 20812 14368
rect 20864 14356 20870 14408
rect 21085 14399 21143 14405
rect 21085 14365 21097 14399
rect 21131 14396 21143 14399
rect 21192 14396 21220 14504
rect 21269 14467 21327 14473
rect 21269 14433 21281 14467
rect 21315 14433 21327 14467
rect 21269 14427 21327 14433
rect 21131 14368 21220 14396
rect 21131 14365 21143 14368
rect 21085 14359 21143 14365
rect 17034 14328 17040 14340
rect 15120 14300 15410 14328
rect 16868 14300 17040 14328
rect 15120 14272 15148 14300
rect 17034 14288 17040 14300
rect 17092 14288 17098 14340
rect 17129 14331 17187 14337
rect 17129 14297 17141 14331
rect 17175 14328 17187 14331
rect 17218 14328 17224 14340
rect 17175 14300 17224 14328
rect 17175 14297 17187 14300
rect 17129 14291 17187 14297
rect 17218 14288 17224 14300
rect 17276 14288 17282 14340
rect 17586 14288 17592 14340
rect 17644 14288 17650 14340
rect 19150 14288 19156 14340
rect 19208 14328 19214 14340
rect 21284 14328 21312 14427
rect 22278 14424 22284 14476
rect 22336 14424 22342 14476
rect 22646 14424 22652 14476
rect 22704 14464 22710 14476
rect 25133 14467 25191 14473
rect 25133 14464 25145 14467
rect 22704 14436 25145 14464
rect 22704 14424 22710 14436
rect 25133 14433 25145 14436
rect 25179 14464 25191 14467
rect 26329 14467 26387 14473
rect 26329 14464 26341 14467
rect 25179 14436 26341 14464
rect 25179 14433 25191 14436
rect 25133 14427 25191 14433
rect 26329 14433 26341 14436
rect 26375 14464 26387 14467
rect 26602 14464 26608 14476
rect 26375 14436 26608 14464
rect 26375 14433 26387 14436
rect 26329 14427 26387 14433
rect 26602 14424 26608 14436
rect 26660 14424 26666 14476
rect 24854 14396 24860 14408
rect 23860 14368 24860 14396
rect 19208 14300 21312 14328
rect 19208 14288 19214 14300
rect 21450 14288 21456 14340
rect 21508 14328 21514 14340
rect 22557 14331 22615 14337
rect 22557 14328 22569 14331
rect 21508 14300 22569 14328
rect 21508 14288 21514 14300
rect 22557 14297 22569 14300
rect 22603 14297 22615 14331
rect 22557 14291 22615 14297
rect 23566 14288 23572 14340
rect 23624 14288 23630 14340
rect 13906 14260 13912 14272
rect 12360 14232 13912 14260
rect 13906 14220 13912 14232
rect 13964 14220 13970 14272
rect 15102 14220 15108 14272
rect 15160 14220 15166 14272
rect 15194 14220 15200 14272
rect 15252 14260 15258 14272
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 15252 14232 16405 14260
rect 15252 14220 15258 14232
rect 16393 14229 16405 14232
rect 16439 14229 16451 14263
rect 16393 14223 16451 14229
rect 19426 14220 19432 14272
rect 19484 14260 19490 14272
rect 20717 14263 20775 14269
rect 20717 14260 20729 14263
rect 19484 14232 20729 14260
rect 19484 14220 19490 14232
rect 20717 14229 20729 14232
rect 20763 14229 20775 14263
rect 20717 14223 20775 14229
rect 21177 14263 21235 14269
rect 21177 14229 21189 14263
rect 21223 14260 21235 14263
rect 21634 14260 21640 14272
rect 21223 14232 21640 14260
rect 21223 14229 21235 14232
rect 21177 14223 21235 14229
rect 21634 14220 21640 14232
rect 21692 14220 21698 14272
rect 22094 14220 22100 14272
rect 22152 14260 22158 14272
rect 23860 14260 23888 14368
rect 24854 14356 24860 14368
rect 24912 14356 24918 14408
rect 24949 14399 25007 14405
rect 24949 14365 24961 14399
rect 24995 14396 25007 14399
rect 25222 14396 25228 14408
rect 24995 14368 25228 14396
rect 24995 14365 25007 14368
rect 24949 14359 25007 14365
rect 25222 14356 25228 14368
rect 25280 14356 25286 14408
rect 25774 14356 25780 14408
rect 25832 14396 25838 14408
rect 26237 14399 26295 14405
rect 26237 14396 26249 14399
rect 25832 14368 26249 14396
rect 25832 14356 25838 14368
rect 26237 14365 26249 14368
rect 26283 14365 26295 14399
rect 26237 14359 26295 14365
rect 27522 14356 27528 14408
rect 27580 14396 27586 14408
rect 35802 14396 35808 14408
rect 27580 14368 35808 14396
rect 27580 14356 27586 14368
rect 35802 14356 35808 14368
rect 35860 14356 35866 14408
rect 25682 14328 25688 14340
rect 24044 14300 25688 14328
rect 22152 14232 23888 14260
rect 22152 14220 22158 14232
rect 23934 14220 23940 14272
rect 23992 14260 23998 14272
rect 24044 14269 24072 14300
rect 25682 14288 25688 14300
rect 25740 14288 25746 14340
rect 26142 14288 26148 14340
rect 26200 14288 26206 14340
rect 24029 14263 24087 14269
rect 24029 14260 24041 14263
rect 23992 14232 24041 14260
rect 23992 14220 23998 14232
rect 24029 14229 24041 14232
rect 24075 14229 24087 14263
rect 24029 14223 24087 14229
rect 24581 14263 24639 14269
rect 24581 14229 24593 14263
rect 24627 14260 24639 14263
rect 24854 14260 24860 14272
rect 24627 14232 24860 14260
rect 24627 14229 24639 14232
rect 24581 14223 24639 14229
rect 24854 14220 24860 14232
rect 24912 14220 24918 14272
rect 25041 14263 25099 14269
rect 25041 14229 25053 14263
rect 25087 14260 25099 14263
rect 25130 14260 25136 14272
rect 25087 14232 25136 14260
rect 25087 14229 25099 14232
rect 25041 14223 25099 14229
rect 25130 14220 25136 14232
rect 25188 14220 25194 14272
rect 25774 14220 25780 14272
rect 25832 14220 25838 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 4614 14016 4620 14068
rect 4672 14056 4678 14068
rect 5261 14059 5319 14065
rect 5261 14056 5273 14059
rect 4672 14028 5273 14056
rect 4672 14016 4678 14028
rect 5261 14025 5273 14028
rect 5307 14025 5319 14059
rect 5261 14019 5319 14025
rect 5629 14059 5687 14065
rect 5629 14025 5641 14059
rect 5675 14056 5687 14059
rect 6362 14056 6368 14068
rect 5675 14028 6368 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 6917 14059 6975 14065
rect 6917 14025 6929 14059
rect 6963 14025 6975 14059
rect 6917 14019 6975 14025
rect 4522 13988 4528 14000
rect 3436 13960 4528 13988
rect 3436 13929 3464 13960
rect 4522 13948 4528 13960
rect 4580 13948 4586 14000
rect 6932 13988 6960 14019
rect 7282 14016 7288 14068
rect 7340 14016 7346 14068
rect 8573 14059 8631 14065
rect 8573 14025 8585 14059
rect 8619 14056 8631 14059
rect 8662 14056 8668 14068
rect 8619 14028 8668 14056
rect 8619 14025 8631 14028
rect 8573 14019 8631 14025
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 9600 14028 10916 14056
rect 9600 13997 9628 14028
rect 8481 13991 8539 13997
rect 8481 13988 8493 13991
rect 6932 13960 8493 13988
rect 8481 13957 8493 13960
rect 8527 13957 8539 13991
rect 8481 13951 8539 13957
rect 9585 13991 9643 13997
rect 9585 13957 9597 13991
rect 9631 13957 9643 13991
rect 9585 13951 9643 13957
rect 10042 13948 10048 14000
rect 10100 13948 10106 14000
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13920 3019 13923
rect 3421 13923 3479 13929
rect 3421 13920 3433 13923
rect 3007 13892 3433 13920
rect 3007 13889 3019 13892
rect 2961 13883 3019 13889
rect 3421 13889 3433 13892
rect 3467 13889 3479 13923
rect 3421 13883 3479 13889
rect 3694 13880 3700 13932
rect 3752 13880 3758 13932
rect 5166 13880 5172 13932
rect 5224 13920 5230 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 5224 13892 7389 13920
rect 5224 13880 5230 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 10888 13920 10916 14028
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11112 14028 11989 14056
rect 11112 14016 11118 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 11977 14019 12035 14025
rect 12452 14028 14749 14056
rect 11146 13948 11152 14000
rect 11204 13988 11210 14000
rect 12345 13991 12403 13997
rect 12345 13988 12357 13991
rect 11204 13960 12357 13988
rect 11204 13948 11210 13960
rect 12345 13957 12357 13960
rect 12391 13957 12403 13991
rect 12345 13951 12403 13957
rect 10888 13892 11192 13920
rect 7377 13883 7435 13889
rect 5718 13812 5724 13864
rect 5776 13812 5782 13864
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13821 5871 13855
rect 5813 13815 5871 13821
rect 5828 13784 5856 13815
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7558 13852 7564 13864
rect 7156 13824 7564 13852
rect 7156 13812 7162 13824
rect 7558 13812 7564 13824
rect 7616 13852 7622 13864
rect 8478 13852 8484 13864
rect 7616 13824 8484 13852
rect 7616 13812 7622 13824
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 5902 13784 5908 13796
rect 5828 13756 5908 13784
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 7282 13744 7288 13796
rect 7340 13784 7346 13796
rect 8202 13784 8208 13796
rect 7340 13756 8208 13784
rect 7340 13744 7346 13756
rect 8202 13744 8208 13756
rect 8260 13784 8266 13796
rect 8680 13784 8708 13815
rect 9306 13812 9312 13864
rect 9364 13812 9370 13864
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 11057 13855 11115 13861
rect 11057 13852 11069 13855
rect 9640 13824 11069 13852
rect 9640 13812 9646 13824
rect 11057 13821 11069 13824
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 8260 13756 8708 13784
rect 11164 13784 11192 13892
rect 11238 13880 11244 13932
rect 11296 13920 11302 13932
rect 11606 13920 11612 13932
rect 11296 13892 11612 13920
rect 11296 13880 11302 13892
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 11698 13880 11704 13932
rect 11756 13920 11762 13932
rect 12452 13929 12480 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 14737 14019 14795 14025
rect 14826 14016 14832 14068
rect 14884 14016 14890 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 18322 14056 18328 14068
rect 15611 14028 18328 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 18414 14016 18420 14068
rect 18472 14056 18478 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 18472 14028 18889 14056
rect 18472 14016 18478 14028
rect 18877 14025 18889 14028
rect 18923 14025 18935 14059
rect 18877 14019 18935 14025
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 20165 14059 20223 14065
rect 20165 14056 20177 14059
rect 19300 14028 20177 14056
rect 19300 14016 19306 14028
rect 20165 14025 20177 14028
rect 20211 14025 20223 14059
rect 20165 14019 20223 14025
rect 21082 14016 21088 14068
rect 21140 14056 21146 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 21140 14028 23397 14056
rect 21140 14016 21146 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 23566 14016 23572 14068
rect 23624 14056 23630 14068
rect 24581 14059 24639 14065
rect 24581 14056 24593 14059
rect 23624 14028 24593 14056
rect 23624 14016 23630 14028
rect 24581 14025 24593 14028
rect 24627 14025 24639 14059
rect 24581 14019 24639 14025
rect 24949 14059 25007 14065
rect 24949 14025 24961 14059
rect 24995 14056 25007 14059
rect 25774 14056 25780 14068
rect 24995 14028 25780 14056
rect 24995 14025 25007 14028
rect 24949 14019 25007 14025
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 13633 13991 13691 13997
rect 13633 13988 13645 13991
rect 12544 13960 13645 13988
rect 12437 13923 12495 13929
rect 12437 13920 12449 13923
rect 11756 13892 12449 13920
rect 11756 13880 11762 13892
rect 12437 13889 12449 13892
rect 12483 13889 12495 13923
rect 12437 13883 12495 13889
rect 11624 13852 11652 13880
rect 12544 13852 12572 13960
rect 13633 13957 13645 13960
rect 13679 13957 13691 13991
rect 13633 13951 13691 13957
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 16390 13988 16396 14000
rect 15344 13960 16396 13988
rect 15344 13948 15350 13960
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 17402 13948 17408 14000
rect 17460 13948 17466 14000
rect 17678 13948 17684 14000
rect 17736 13988 17742 14000
rect 17736 13960 17894 13988
rect 17736 13948 17742 13960
rect 18690 13948 18696 14000
rect 18748 13988 18754 14000
rect 22094 13988 22100 14000
rect 18748 13960 22100 13988
rect 18748 13948 18754 13960
rect 22094 13948 22100 13960
rect 22152 13948 22158 14000
rect 22186 13948 22192 14000
rect 22244 13988 22250 14000
rect 22557 13991 22615 13997
rect 22557 13988 22569 13991
rect 22244 13960 22569 13988
rect 22244 13948 22250 13960
rect 22557 13957 22569 13960
rect 22603 13957 22615 13991
rect 22557 13951 22615 13957
rect 22649 13991 22707 13997
rect 22649 13957 22661 13991
rect 22695 13988 22707 13991
rect 22922 13988 22928 14000
rect 22695 13960 22928 13988
rect 22695 13957 22707 13960
rect 22649 13951 22707 13957
rect 12802 13880 12808 13932
rect 12860 13920 12866 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 12860 13892 13553 13920
rect 12860 13880 12866 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 15378 13920 15384 13932
rect 13541 13883 13599 13889
rect 13648 13892 15384 13920
rect 11624 13824 12572 13852
rect 12621 13855 12679 13861
rect 12621 13821 12633 13855
rect 12667 13821 12679 13855
rect 13648 13852 13676 13892
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13920 15991 13923
rect 16206 13920 16212 13932
rect 15979 13892 16212 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 18782 13880 18788 13932
rect 18840 13920 18846 13932
rect 18966 13920 18972 13932
rect 18840 13892 18972 13920
rect 18840 13880 18846 13892
rect 18966 13880 18972 13892
rect 19024 13880 19030 13932
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13920 19671 13923
rect 20070 13920 20076 13932
rect 19659 13892 20076 13920
rect 19659 13889 19671 13892
rect 19613 13883 19671 13889
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13889 20591 13923
rect 20533 13883 20591 13889
rect 20625 13923 20683 13929
rect 20625 13889 20637 13923
rect 20671 13920 20683 13923
rect 21358 13920 21364 13932
rect 20671 13892 21364 13920
rect 20671 13889 20683 13892
rect 20625 13883 20683 13889
rect 12621 13815 12679 13821
rect 13188 13824 13676 13852
rect 13817 13855 13875 13861
rect 12158 13784 12164 13796
rect 11164 13756 12164 13784
rect 8260 13744 8266 13756
rect 12158 13744 12164 13756
rect 12216 13784 12222 13796
rect 12636 13784 12664 13815
rect 13188 13793 13216 13824
rect 13817 13821 13829 13855
rect 13863 13821 13875 13855
rect 14458 13852 14464 13864
rect 13817 13815 13875 13821
rect 14384 13824 14464 13852
rect 12216 13756 12664 13784
rect 13173 13787 13231 13793
rect 12216 13744 12222 13756
rect 13173 13753 13185 13787
rect 13219 13753 13231 13787
rect 13832 13784 13860 13815
rect 14384 13793 14412 13824
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 15013 13855 15071 13861
rect 15013 13821 15025 13855
rect 15059 13852 15071 13855
rect 15194 13852 15200 13864
rect 15059 13824 15200 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 16022 13812 16028 13864
rect 16080 13812 16086 13864
rect 16117 13855 16175 13861
rect 16117 13821 16129 13855
rect 16163 13821 16175 13855
rect 16117 13815 16175 13821
rect 14369 13787 14427 13793
rect 13832 13756 13952 13784
rect 13173 13747 13231 13753
rect 7558 13676 7564 13728
rect 7616 13716 7622 13728
rect 8113 13719 8171 13725
rect 8113 13716 8125 13719
rect 7616 13688 8125 13716
rect 7616 13676 7622 13688
rect 8113 13685 8125 13688
rect 8159 13685 8171 13719
rect 8113 13679 8171 13685
rect 8294 13676 8300 13728
rect 8352 13716 8358 13728
rect 10594 13716 10600 13728
rect 8352 13688 10600 13716
rect 8352 13676 8358 13688
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 11146 13676 11152 13728
rect 11204 13716 11210 13728
rect 12434 13716 12440 13728
rect 11204 13688 12440 13716
rect 11204 13676 11210 13688
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 13924 13716 13952 13756
rect 14369 13753 14381 13787
rect 14415 13753 14427 13787
rect 14369 13747 14427 13753
rect 15378 13716 15384 13728
rect 13924 13688 15384 13716
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 16132 13716 16160 13815
rect 16298 13812 16304 13864
rect 16356 13852 16362 13864
rect 16356 13824 16988 13852
rect 16356 13812 16362 13824
rect 16960 13784 16988 13824
rect 17034 13812 17040 13864
rect 17092 13852 17098 13864
rect 17129 13855 17187 13861
rect 17129 13852 17141 13855
rect 17092 13824 17141 13852
rect 17092 13812 17098 13824
rect 17129 13821 17141 13824
rect 17175 13821 17187 13855
rect 20548 13852 20576 13883
rect 21358 13880 21364 13892
rect 21416 13880 21422 13932
rect 22572 13920 22600 13951
rect 22922 13948 22928 13960
rect 22980 13988 22986 14000
rect 22980 13960 23888 13988
rect 22980 13948 22986 13960
rect 23860 13929 23888 13960
rect 24854 13948 24860 14000
rect 24912 13988 24918 14000
rect 25041 13991 25099 13997
rect 25041 13988 25053 13991
rect 24912 13960 25053 13988
rect 24912 13948 24918 13960
rect 25041 13957 25053 13960
rect 25087 13957 25099 13991
rect 25041 13951 25099 13957
rect 23753 13923 23811 13929
rect 23753 13920 23765 13923
rect 22572 13892 23765 13920
rect 23753 13889 23765 13892
rect 23799 13889 23811 13923
rect 23753 13883 23811 13889
rect 23845 13923 23903 13929
rect 23845 13889 23857 13923
rect 23891 13920 23903 13923
rect 23891 13892 31754 13920
rect 23891 13889 23903 13892
rect 23845 13883 23903 13889
rect 17129 13815 17187 13821
rect 17236 13824 20576 13852
rect 20809 13855 20867 13861
rect 17236 13784 17264 13824
rect 20809 13821 20821 13855
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 16960 13756 17264 13784
rect 19429 13787 19487 13793
rect 19429 13753 19441 13787
rect 19475 13784 19487 13787
rect 19794 13784 19800 13796
rect 19475 13756 19800 13784
rect 19475 13753 19487 13756
rect 19429 13747 19487 13753
rect 19794 13744 19800 13756
rect 19852 13744 19858 13796
rect 20824 13784 20852 13815
rect 22738 13812 22744 13864
rect 22796 13812 22802 13864
rect 23937 13855 23995 13861
rect 23937 13821 23949 13855
rect 23983 13821 23995 13855
rect 23937 13815 23995 13821
rect 25133 13855 25191 13861
rect 25133 13821 25145 13855
rect 25179 13821 25191 13855
rect 31726 13852 31754 13892
rect 49234 13852 49240 13864
rect 31726 13824 49240 13852
rect 25133 13815 25191 13821
rect 21818 13784 21824 13796
rect 20824 13756 21824 13784
rect 21818 13744 21824 13756
rect 21876 13744 21882 13796
rect 23842 13744 23848 13796
rect 23900 13784 23906 13796
rect 23952 13784 23980 13815
rect 24026 13784 24032 13796
rect 23900 13756 24032 13784
rect 23900 13744 23906 13756
rect 24026 13744 24032 13756
rect 24084 13744 24090 13796
rect 25148 13728 25176 13815
rect 49234 13812 49240 13824
rect 49292 13812 49298 13864
rect 18966 13716 18972 13728
rect 16132 13688 18972 13716
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 21174 13716 21180 13728
rect 19576 13688 21180 13716
rect 19576 13676 19582 13688
rect 21174 13676 21180 13688
rect 21232 13676 21238 13728
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 22189 13719 22247 13725
rect 22189 13716 22201 13719
rect 22152 13688 22201 13716
rect 22152 13676 22158 13688
rect 22189 13685 22201 13688
rect 22235 13685 22247 13719
rect 22189 13679 22247 13685
rect 25130 13676 25136 13728
rect 25188 13676 25194 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 3988 13484 13400 13512
rect 2774 13336 2780 13388
rect 2832 13336 2838 13388
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13308 1823 13311
rect 3988 13308 4016 13484
rect 8202 13404 8208 13456
rect 8260 13444 8266 13456
rect 8481 13447 8539 13453
rect 8481 13444 8493 13447
rect 8260 13416 8493 13444
rect 8260 13404 8266 13416
rect 8481 13413 8493 13416
rect 8527 13444 8539 13447
rect 13372 13444 13400 13484
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 13725 13515 13783 13521
rect 13725 13512 13737 13515
rect 13504 13484 13737 13512
rect 13504 13472 13510 13484
rect 13725 13481 13737 13484
rect 13771 13481 13783 13515
rect 13725 13475 13783 13481
rect 15010 13472 15016 13524
rect 15068 13512 15074 13524
rect 15068 13484 15700 13512
rect 15068 13472 15074 13484
rect 15672 13456 15700 13484
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 17460 13484 18889 13512
rect 17460 13472 17466 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 21358 13472 21364 13524
rect 21416 13512 21422 13524
rect 22833 13515 22891 13521
rect 22833 13512 22845 13515
rect 21416 13484 22845 13512
rect 21416 13472 21422 13484
rect 22833 13481 22845 13484
rect 22879 13481 22891 13515
rect 22833 13475 22891 13481
rect 14090 13444 14096 13456
rect 8527 13416 10824 13444
rect 13372 13416 14096 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 4157 13379 4215 13385
rect 4157 13345 4169 13379
rect 4203 13376 4215 13379
rect 4798 13376 4804 13388
rect 4203 13348 4804 13376
rect 4203 13345 4215 13348
rect 4157 13339 4215 13345
rect 4798 13336 4804 13348
rect 4856 13376 4862 13388
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 4856 13348 6745 13376
rect 4856 13336 4862 13348
rect 6733 13345 6745 13348
rect 6779 13376 6791 13379
rect 8294 13376 8300 13388
rect 6779 13348 8300 13376
rect 6779 13345 6791 13348
rect 6733 13339 6791 13345
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 10796 13385 10824 13416
rect 14090 13404 14096 13416
rect 14148 13404 14154 13456
rect 15654 13404 15660 13456
rect 15712 13444 15718 13456
rect 16025 13447 16083 13453
rect 16025 13444 16037 13447
rect 15712 13416 16037 13444
rect 15712 13404 15718 13416
rect 16025 13413 16037 13416
rect 16071 13413 16083 13447
rect 16025 13407 16083 13413
rect 22097 13447 22155 13453
rect 22097 13413 22109 13447
rect 22143 13444 22155 13447
rect 22462 13444 22468 13456
rect 22143 13416 22468 13444
rect 22143 13413 22155 13416
rect 22097 13407 22155 13413
rect 22462 13404 22468 13416
rect 22520 13404 22526 13456
rect 10781 13379 10839 13385
rect 10781 13345 10793 13379
rect 10827 13345 10839 13379
rect 10781 13339 10839 13345
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 12032 13348 14289 13376
rect 12032 13336 12038 13348
rect 14277 13345 14289 13348
rect 14323 13376 14335 13379
rect 14642 13376 14648 13388
rect 14323 13348 14648 13376
rect 14323 13345 14335 13348
rect 14277 13339 14335 13345
rect 14642 13336 14648 13348
rect 14700 13376 14706 13388
rect 15838 13376 15844 13388
rect 14700 13348 15844 13376
rect 14700 13336 14706 13348
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 17034 13336 17040 13388
rect 17092 13376 17098 13388
rect 17129 13379 17187 13385
rect 17129 13376 17141 13379
rect 17092 13348 17141 13376
rect 17092 13336 17098 13348
rect 17129 13345 17141 13348
rect 17175 13376 17187 13379
rect 17494 13376 17500 13388
rect 17175 13348 17500 13376
rect 17175 13345 17187 13348
rect 17129 13339 17187 13345
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 20349 13379 20407 13385
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 22186 13376 22192 13388
rect 20395 13348 22192 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 22186 13336 22192 13348
rect 22244 13336 22250 13388
rect 23293 13379 23351 13385
rect 23293 13345 23305 13379
rect 23339 13376 23351 13379
rect 23382 13376 23388 13388
rect 23339 13348 23388 13376
rect 23339 13345 23351 13348
rect 23293 13339 23351 13345
rect 23382 13336 23388 13348
rect 23440 13336 23446 13388
rect 23474 13336 23480 13388
rect 23532 13336 23538 13388
rect 1811 13280 4016 13308
rect 1811 13277 1823 13280
rect 1765 13271 1823 13277
rect 9766 13268 9772 13320
rect 9824 13268 9830 13320
rect 16666 13268 16672 13320
rect 16724 13268 16730 13320
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 19613 13311 19671 13317
rect 19613 13308 19625 13311
rect 19392 13280 19625 13308
rect 19392 13268 19398 13280
rect 19613 13277 19625 13280
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 23014 13268 23020 13320
rect 23072 13308 23078 13320
rect 23072 13280 25452 13308
rect 23072 13268 23078 13280
rect 4433 13243 4491 13249
rect 4433 13209 4445 13243
rect 4479 13240 4491 13243
rect 4522 13240 4528 13252
rect 4479 13212 4528 13240
rect 4479 13209 4491 13212
rect 4433 13203 4491 13209
rect 4522 13200 4528 13212
rect 4580 13200 4586 13252
rect 6270 13240 6276 13252
rect 5658 13212 6276 13240
rect 6270 13200 6276 13212
rect 6328 13240 6334 13252
rect 6638 13240 6644 13252
rect 6328 13212 6644 13240
rect 6328 13200 6334 13212
rect 6638 13200 6644 13212
rect 6696 13200 6702 13252
rect 7009 13243 7067 13249
rect 7009 13209 7021 13243
rect 7055 13240 7067 13243
rect 7098 13240 7104 13252
rect 7055 13212 7104 13240
rect 7055 13209 7067 13212
rect 7009 13203 7067 13209
rect 7098 13200 7104 13212
rect 7156 13200 7162 13252
rect 10597 13243 10655 13249
rect 7208 13212 7498 13240
rect 8312 13212 10272 13240
rect 5902 13132 5908 13184
rect 5960 13132 5966 13184
rect 6656 13172 6684 13200
rect 7208 13172 7236 13212
rect 6656 13144 7236 13172
rect 7374 13132 7380 13184
rect 7432 13172 7438 13184
rect 8312 13172 8340 13212
rect 7432 13144 8340 13172
rect 7432 13132 7438 13144
rect 8570 13132 8576 13184
rect 8628 13172 8634 13184
rect 10244 13181 10272 13212
rect 10597 13209 10609 13243
rect 10643 13240 10655 13243
rect 12253 13243 12311 13249
rect 10643 13212 11560 13240
rect 10643 13209 10655 13212
rect 10597 13203 10655 13209
rect 9585 13175 9643 13181
rect 9585 13172 9597 13175
rect 8628 13144 9597 13172
rect 8628 13132 8634 13144
rect 9585 13141 9597 13144
rect 9631 13141 9643 13175
rect 9585 13135 9643 13141
rect 10229 13175 10287 13181
rect 10229 13141 10241 13175
rect 10275 13141 10287 13175
rect 10229 13135 10287 13141
rect 10686 13132 10692 13184
rect 10744 13132 10750 13184
rect 11532 13172 11560 13212
rect 12253 13209 12265 13243
rect 12299 13240 12311 13243
rect 12342 13240 12348 13252
rect 12299 13212 12348 13240
rect 12299 13209 12311 13212
rect 12253 13203 12311 13209
rect 12342 13200 12348 13212
rect 12400 13200 12406 13252
rect 12526 13200 12532 13252
rect 12584 13240 12590 13252
rect 12710 13240 12716 13252
rect 12584 13212 12716 13240
rect 12584 13200 12590 13212
rect 12710 13200 12716 13212
rect 12768 13200 12774 13252
rect 14553 13243 14611 13249
rect 14553 13209 14565 13243
rect 14599 13209 14611 13243
rect 14553 13203 14611 13209
rect 13630 13172 13636 13184
rect 11532 13144 13636 13172
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 14568 13172 14596 13203
rect 15010 13200 15016 13252
rect 15068 13200 15074 13252
rect 17405 13243 17463 13249
rect 17405 13240 17417 13243
rect 16040 13212 17417 13240
rect 15194 13172 15200 13184
rect 14568 13144 15200 13172
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 15378 13132 15384 13184
rect 15436 13172 15442 13184
rect 16040 13172 16068 13212
rect 17405 13209 17417 13212
rect 17451 13209 17463 13243
rect 17405 13203 17463 13209
rect 15436 13144 16068 13172
rect 15436 13132 15442 13144
rect 16482 13132 16488 13184
rect 16540 13132 16546 13184
rect 17420 13172 17448 13203
rect 17678 13200 17684 13252
rect 17736 13240 17742 13252
rect 17736 13212 17894 13240
rect 17736 13200 17742 13212
rect 18966 13200 18972 13252
rect 19024 13240 19030 13252
rect 20625 13243 20683 13249
rect 20625 13240 20637 13243
rect 19024 13212 20637 13240
rect 19024 13200 19030 13212
rect 20625 13209 20637 13212
rect 20671 13209 20683 13243
rect 20625 13203 20683 13209
rect 21634 13200 21640 13252
rect 21692 13200 21698 13252
rect 23201 13243 23259 13249
rect 23201 13209 23213 13243
rect 23247 13240 23259 13243
rect 24118 13240 24124 13252
rect 23247 13212 24124 13240
rect 23247 13209 23259 13212
rect 23201 13203 23259 13209
rect 24118 13200 24124 13212
rect 24176 13200 24182 13252
rect 24578 13200 24584 13252
rect 24636 13200 24642 13252
rect 25424 13249 25452 13280
rect 25409 13243 25467 13249
rect 25409 13209 25421 13243
rect 25455 13240 25467 13243
rect 26878 13240 26884 13252
rect 25455 13212 26884 13240
rect 25455 13209 25467 13212
rect 25409 13203 25467 13209
rect 26878 13200 26884 13212
rect 26936 13200 26942 13252
rect 18414 13172 18420 13184
rect 17420 13144 18420 13172
rect 18414 13132 18420 13144
rect 18472 13172 18478 13184
rect 18782 13172 18788 13184
rect 18472 13144 18788 13172
rect 18472 13132 18478 13144
rect 18782 13132 18788 13144
rect 18840 13132 18846 13184
rect 19429 13175 19487 13181
rect 19429 13141 19441 13175
rect 19475 13172 19487 13175
rect 28534 13172 28540 13184
rect 19475 13144 28540 13172
rect 19475 13141 19487 13144
rect 19429 13135 19487 13141
rect 28534 13132 28540 13144
rect 28592 13132 28598 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 3510 12928 3516 12980
rect 3568 12928 3574 12980
rect 4065 12971 4123 12977
rect 4065 12937 4077 12971
rect 4111 12968 4123 12971
rect 5718 12968 5724 12980
rect 4111 12940 5724 12968
rect 4111 12937 4123 12940
rect 4065 12931 4123 12937
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 7374 12928 7380 12980
rect 7432 12928 7438 12980
rect 7469 12971 7527 12977
rect 7469 12937 7481 12971
rect 7515 12968 7527 12971
rect 7558 12968 7564 12980
rect 7515 12940 7564 12968
rect 7515 12937 7527 12940
rect 7469 12931 7527 12937
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 9306 12968 9312 12980
rect 8352 12940 9312 12968
rect 8352 12928 8358 12940
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 12621 12971 12679 12977
rect 12621 12968 12633 12971
rect 11020 12940 12633 12968
rect 11020 12928 11026 12940
rect 12621 12937 12633 12940
rect 12667 12937 12679 12971
rect 12989 12971 13047 12977
rect 12989 12968 13001 12971
rect 12621 12931 12679 12937
rect 12715 12940 13001 12968
rect 2774 12860 2780 12912
rect 2832 12860 2838 12912
rect 3421 12903 3479 12909
rect 3421 12869 3433 12903
rect 3467 12900 3479 12903
rect 3786 12900 3792 12912
rect 3467 12872 3792 12900
rect 3467 12869 3479 12872
rect 3421 12863 3479 12869
rect 3786 12860 3792 12872
rect 3844 12860 3850 12912
rect 4430 12860 4436 12912
rect 4488 12860 4494 12912
rect 4522 12860 4528 12912
rect 4580 12900 4586 12912
rect 8312 12900 8340 12928
rect 4580 12872 4752 12900
rect 4580 12860 4586 12872
rect 1762 12792 1768 12844
rect 1820 12792 1826 12844
rect 4522 12724 4528 12776
rect 4580 12724 4586 12776
rect 4724 12773 4752 12872
rect 8220 12872 8340 12900
rect 5626 12792 5632 12844
rect 5684 12792 5690 12844
rect 5721 12835 5779 12841
rect 5721 12801 5733 12835
rect 5767 12832 5779 12835
rect 6730 12832 6736 12844
rect 5767 12804 6736 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 4709 12767 4767 12773
rect 4709 12733 4721 12767
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 4724 12696 4752 12727
rect 5534 12724 5540 12776
rect 5592 12764 5598 12776
rect 5736 12764 5764 12795
rect 6730 12792 6736 12804
rect 6788 12792 6794 12844
rect 8220 12841 8248 12872
rect 8478 12860 8484 12912
rect 8536 12860 8542 12912
rect 8754 12860 8760 12912
rect 8812 12900 8818 12912
rect 8812 12872 8970 12900
rect 8812 12860 8818 12872
rect 10226 12860 10232 12912
rect 10284 12860 10290 12912
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 12715 12900 12743 12940
rect 12989 12937 13001 12940
rect 13035 12937 13047 12971
rect 12989 12931 13047 12937
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 13127 12940 14964 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 14277 12903 14335 12909
rect 14277 12900 14289 12903
rect 12124 12872 12743 12900
rect 12912 12872 14289 12900
rect 12124 12860 12130 12872
rect 8205 12835 8263 12841
rect 7024 12804 8156 12832
rect 5592 12736 5764 12764
rect 5905 12767 5963 12773
rect 5592 12724 5598 12736
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 6270 12764 6276 12776
rect 5951 12736 6276 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 5810 12696 5816 12708
rect 4724 12668 5816 12696
rect 5810 12656 5816 12668
rect 5868 12696 5874 12708
rect 5920 12696 5948 12727
rect 6270 12724 6276 12736
rect 6328 12724 6334 12776
rect 7024 12705 7052 12804
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12733 7711 12767
rect 8128 12764 8156 12804
rect 8205 12801 8217 12835
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 11149 12835 11207 12841
rect 9916 12804 10732 12832
rect 9916 12792 9922 12804
rect 10704 12764 10732 12804
rect 11149 12801 11161 12835
rect 11195 12832 11207 12835
rect 12802 12832 12808 12844
rect 11195 12804 12808 12832
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 12912 12764 12940 12872
rect 14277 12869 14289 12872
rect 14323 12869 14335 12903
rect 14277 12863 14335 12869
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12832 14243 12835
rect 14734 12832 14740 12844
rect 14231 12804 14740 12832
rect 14231 12801 14243 12804
rect 14185 12795 14243 12801
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 14936 12832 14964 12940
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 17957 12971 18015 12977
rect 17957 12968 17969 12971
rect 16080 12940 17969 12968
rect 16080 12928 16086 12940
rect 17957 12937 17969 12940
rect 18003 12937 18015 12971
rect 17957 12931 18015 12937
rect 18325 12971 18383 12977
rect 18325 12937 18337 12971
rect 18371 12968 18383 12971
rect 18371 12940 21220 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 15010 12860 15016 12912
rect 15068 12900 15074 12912
rect 18874 12900 18880 12912
rect 15068 12872 18880 12900
rect 15068 12860 15074 12872
rect 18874 12860 18880 12872
rect 18932 12900 18938 12912
rect 19150 12900 19156 12912
rect 18932 12872 19156 12900
rect 18932 12860 18938 12872
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 21082 12860 21088 12912
rect 21140 12860 21146 12912
rect 17862 12832 17868 12844
rect 14936 12804 17868 12832
rect 17862 12792 17868 12804
rect 17920 12792 17926 12844
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12832 18475 12835
rect 20714 12832 20720 12844
rect 18463 12804 20720 12832
rect 18463 12801 18475 12804
rect 18417 12795 18475 12801
rect 20714 12792 20720 12804
rect 20772 12792 20778 12844
rect 21192 12832 21220 12940
rect 22002 12928 22008 12980
rect 22060 12968 22066 12980
rect 23474 12968 23480 12980
rect 22060 12940 23480 12968
rect 22060 12928 22066 12940
rect 23474 12928 23480 12940
rect 23532 12968 23538 12980
rect 24765 12971 24823 12977
rect 24765 12968 24777 12971
rect 23532 12940 24777 12968
rect 23532 12928 23538 12940
rect 24765 12937 24777 12940
rect 24811 12937 24823 12971
rect 24765 12931 24823 12937
rect 22094 12832 22100 12844
rect 21192 12804 22100 12832
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 23014 12832 23020 12844
rect 22244 12804 23020 12832
rect 22244 12792 22250 12804
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 24394 12792 24400 12844
rect 24452 12792 24458 12844
rect 8128 12736 9812 12764
rect 10704 12736 12940 12764
rect 13265 12767 13323 12773
rect 7653 12727 7711 12733
rect 5868 12668 5948 12696
rect 7009 12699 7067 12705
rect 5868 12656 5874 12668
rect 7009 12665 7021 12699
rect 7055 12665 7067 12699
rect 7009 12659 7067 12665
rect 5258 12588 5264 12640
rect 5316 12588 5322 12640
rect 7668 12628 7696 12727
rect 8478 12628 8484 12640
rect 7668 12600 8484 12628
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 9674 12628 9680 12640
rect 9180 12600 9680 12628
rect 9180 12588 9186 12600
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 9784 12628 9812 12736
rect 13265 12733 13277 12767
rect 13311 12733 13323 12767
rect 13265 12727 13323 12733
rect 12161 12699 12219 12705
rect 12161 12665 12173 12699
rect 12207 12696 12219 12699
rect 13280 12696 13308 12727
rect 14458 12724 14464 12776
rect 14516 12724 14522 12776
rect 15838 12724 15844 12776
rect 15896 12724 15902 12776
rect 15930 12724 15936 12776
rect 15988 12764 15994 12776
rect 16298 12764 16304 12776
rect 15988 12736 16304 12764
rect 15988 12724 15994 12736
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 18601 12767 18659 12773
rect 18601 12733 18613 12767
rect 18647 12764 18659 12767
rect 18782 12764 18788 12776
rect 18647 12736 18788 12764
rect 18647 12733 18659 12736
rect 18601 12727 18659 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12764 20039 12767
rect 20070 12764 20076 12776
rect 20027 12736 20076 12764
rect 20027 12733 20039 12736
rect 19981 12727 20039 12733
rect 15378 12696 15384 12708
rect 12207 12668 12940 12696
rect 13280 12668 15384 12696
rect 12207 12665 12219 12668
rect 12161 12659 12219 12665
rect 12618 12628 12624 12640
rect 9784 12600 12624 12628
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 12912 12628 12940 12668
rect 15378 12656 15384 12668
rect 15436 12656 15442 12708
rect 17494 12656 17500 12708
rect 17552 12696 17558 12708
rect 19996 12696 20024 12727
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 21177 12767 21235 12773
rect 21177 12733 21189 12767
rect 21223 12733 21235 12767
rect 21177 12727 21235 12733
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 21450 12764 21456 12776
rect 21407 12736 21456 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 17552 12668 20024 12696
rect 21192 12696 21220 12727
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 23293 12767 23351 12773
rect 23293 12733 23305 12767
rect 23339 12764 23351 12767
rect 23934 12764 23940 12776
rect 23339 12736 23940 12764
rect 23339 12733 23351 12736
rect 23293 12727 23351 12733
rect 23934 12724 23940 12736
rect 23992 12724 23998 12776
rect 22554 12696 22560 12708
rect 21192 12668 22560 12696
rect 17552 12656 17558 12668
rect 22554 12656 22560 12668
rect 22612 12656 22618 12708
rect 13354 12628 13360 12640
rect 12912 12600 13360 12628
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 13814 12588 13820 12640
rect 13872 12588 13878 12640
rect 15470 12588 15476 12640
rect 15528 12628 15534 12640
rect 17037 12631 17095 12637
rect 17037 12628 17049 12631
rect 15528 12600 17049 12628
rect 15528 12588 15534 12600
rect 17037 12597 17049 12600
rect 17083 12597 17095 12631
rect 17037 12591 17095 12597
rect 20714 12588 20720 12640
rect 20772 12588 20778 12640
rect 23934 12588 23940 12640
rect 23992 12628 23998 12640
rect 24394 12628 24400 12640
rect 23992 12600 24400 12628
rect 23992 12588 23998 12600
rect 24394 12588 24400 12600
rect 24452 12588 24458 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 4065 12427 4123 12433
rect 4065 12393 4077 12427
rect 4111 12424 4123 12427
rect 4522 12424 4528 12436
rect 4111 12396 4528 12424
rect 4111 12393 4123 12396
rect 4065 12387 4123 12393
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 6086 12384 6092 12436
rect 6144 12424 6150 12436
rect 6362 12424 6368 12436
rect 6144 12396 6368 12424
rect 6144 12384 6150 12396
rect 6362 12384 6368 12396
rect 6420 12384 6426 12436
rect 7374 12384 7380 12436
rect 7432 12384 7438 12436
rect 7466 12384 7472 12436
rect 7524 12424 7530 12436
rect 7742 12424 7748 12436
rect 7524 12396 7748 12424
rect 7524 12384 7530 12396
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 7837 12427 7895 12433
rect 7837 12393 7849 12427
rect 7883 12424 7895 12427
rect 10686 12424 10692 12436
rect 7883 12396 10692 12424
rect 7883 12393 7895 12396
rect 7837 12387 7895 12393
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 11793 12427 11851 12433
rect 11793 12393 11805 12427
rect 11839 12424 11851 12427
rect 11974 12424 11980 12436
rect 11839 12396 11980 12424
rect 11839 12393 11851 12396
rect 11793 12387 11851 12393
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 15746 12424 15752 12436
rect 13035 12396 15752 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 18049 12427 18107 12433
rect 18049 12393 18061 12427
rect 18095 12424 18107 12427
rect 18414 12424 18420 12436
rect 18095 12396 18420 12424
rect 18095 12393 18107 12396
rect 18049 12387 18107 12393
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 21818 12384 21824 12436
rect 21876 12424 21882 12436
rect 21876 12396 22094 12424
rect 21876 12384 21882 12396
rect 3418 12316 3424 12368
rect 3476 12316 3482 12368
rect 5350 12356 5356 12368
rect 4080 12328 5356 12356
rect 1578 12248 1584 12300
rect 1636 12248 1642 12300
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12288 1915 12291
rect 4080 12288 4108 12328
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 7392 12356 7420 12384
rect 10410 12356 10416 12368
rect 7392 12328 8248 12356
rect 1903 12260 4108 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 4706 12248 4712 12300
rect 4764 12248 4770 12300
rect 7377 12291 7435 12297
rect 7377 12257 7389 12291
rect 7423 12288 7435 12291
rect 7650 12288 7656 12300
rect 7423 12260 7656 12288
rect 7423 12257 7435 12260
rect 7377 12251 7435 12257
rect 7650 12248 7656 12260
rect 7708 12248 7714 12300
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12220 2651 12223
rect 2866 12220 2872 12232
rect 2639 12192 2872 12220
rect 2639 12189 2651 12192
rect 2593 12183 2651 12189
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 3142 12180 3148 12232
rect 3200 12220 3206 12232
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 3200 12192 3249 12220
rect 3200 12180 3206 12192
rect 3237 12189 3249 12192
rect 3283 12220 3295 12223
rect 4338 12220 4344 12232
rect 3283 12192 4344 12220
rect 3283 12189 3295 12192
rect 3237 12183 3295 12189
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 4430 12180 4436 12232
rect 4488 12180 4494 12232
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 8220 12229 8248 12328
rect 8312 12328 10416 12356
rect 8312 12297 8340 12328
rect 10410 12316 10416 12328
rect 10468 12316 10474 12368
rect 15286 12356 15292 12368
rect 10520 12328 15292 12356
rect 8297 12291 8355 12297
rect 8297 12257 8309 12291
rect 8343 12257 8355 12291
rect 8297 12251 8355 12257
rect 8481 12291 8539 12297
rect 8481 12257 8493 12291
rect 8527 12288 8539 12291
rect 8570 12288 8576 12300
rect 8527 12260 8576 12288
rect 8527 12257 8539 12260
rect 8481 12251 8539 12257
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 9364 12260 9873 12288
rect 9364 12248 9370 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 10520 12288 10548 12328
rect 15286 12316 15292 12328
rect 15344 12316 15350 12368
rect 19996 12328 20208 12356
rect 9861 12251 9919 12257
rect 9968 12260 10548 12288
rect 5353 12223 5411 12229
rect 5353 12220 5365 12223
rect 4856 12192 5365 12220
rect 4856 12180 4862 12192
rect 5353 12189 5365 12192
rect 5399 12189 5411 12223
rect 5353 12183 5411 12189
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12189 8263 12223
rect 8205 12183 8263 12189
rect 8386 12180 8392 12232
rect 8444 12220 8450 12232
rect 8846 12220 8852 12232
rect 8444 12192 8852 12220
rect 8444 12180 8450 12192
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9968 12220 9996 12260
rect 10778 12248 10784 12300
rect 10836 12248 10842 12300
rect 12342 12248 12348 12300
rect 12400 12248 12406 12300
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 14826 12288 14832 12300
rect 13679 12260 14832 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 15838 12248 15844 12300
rect 15896 12288 15902 12300
rect 16301 12291 16359 12297
rect 16301 12288 16313 12291
rect 15896 12260 16313 12288
rect 15896 12248 15902 12260
rect 16301 12257 16313 12260
rect 16347 12257 16359 12291
rect 16301 12251 16359 12257
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 17310 12288 17316 12300
rect 16724 12260 17316 12288
rect 16724 12248 16730 12260
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 9232 12192 9996 12220
rect 10505 12223 10563 12229
rect 2774 12112 2780 12164
rect 2832 12112 2838 12164
rect 4525 12155 4583 12161
rect 4525 12152 4537 12155
rect 3620 12124 4537 12152
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 3620 12084 3648 12124
rect 4525 12121 4537 12124
rect 4571 12121 4583 12155
rect 4525 12115 4583 12121
rect 5629 12155 5687 12161
rect 5629 12121 5641 12155
rect 5675 12152 5687 12155
rect 5718 12152 5724 12164
rect 5675 12124 5724 12152
rect 5675 12121 5687 12124
rect 5629 12115 5687 12121
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 6638 12112 6644 12164
rect 6696 12112 6702 12164
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 9232 12152 9260 12192
rect 10505 12189 10517 12223
rect 10551 12220 10563 12223
rect 11974 12220 11980 12232
rect 10551 12192 11980 12220
rect 10551 12189 10563 12192
rect 10505 12183 10563 12189
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 12253 12223 12311 12229
rect 12253 12189 12265 12223
rect 12299 12220 12311 12223
rect 16114 12220 16120 12232
rect 12299 12192 16120 12220
rect 12299 12189 12311 12192
rect 12253 12183 12311 12189
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 6972 12124 9260 12152
rect 6972 12112 6978 12124
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 14369 12155 14427 12161
rect 14369 12152 14381 12155
rect 9732 12124 14381 12152
rect 9732 12112 9738 12124
rect 14369 12121 14381 12124
rect 14415 12152 14427 12155
rect 15010 12152 15016 12164
rect 14415 12124 15016 12152
rect 14415 12121 14427 12124
rect 14369 12115 14427 12121
rect 15010 12112 15016 12124
rect 15068 12112 15074 12164
rect 15102 12112 15108 12164
rect 15160 12112 15166 12164
rect 15378 12112 15384 12164
rect 15436 12152 15442 12164
rect 16482 12152 16488 12164
rect 15436 12124 16488 12152
rect 15436 12112 15442 12124
rect 16482 12112 16488 12124
rect 16540 12152 16546 12164
rect 16577 12155 16635 12161
rect 16577 12152 16589 12155
rect 16540 12124 16589 12152
rect 16540 12112 16546 12124
rect 16577 12121 16589 12124
rect 16623 12121 16635 12155
rect 16577 12115 16635 12121
rect 17034 12112 17040 12164
rect 17092 12112 17098 12164
rect 19996 12152 20024 12328
rect 20070 12248 20076 12300
rect 20128 12248 20134 12300
rect 20180 12288 20208 12328
rect 21910 12288 21916 12300
rect 20180 12260 21916 12288
rect 21910 12248 21916 12260
rect 21968 12248 21974 12300
rect 22066 12288 22094 12396
rect 22557 12291 22615 12297
rect 22557 12288 22569 12291
rect 22066 12260 22569 12288
rect 22557 12257 22569 12260
rect 22603 12257 22615 12291
rect 22557 12251 22615 12257
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 22281 12223 22339 12229
rect 22281 12220 22293 12223
rect 22244 12192 22293 12220
rect 22244 12180 22250 12192
rect 22281 12189 22293 12192
rect 22327 12189 22339 12223
rect 22281 12183 22339 12189
rect 20349 12155 20407 12161
rect 20349 12152 20361 12155
rect 18156 12124 20361 12152
rect 2096 12056 3648 12084
rect 2096 12044 2102 12056
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 12161 12087 12219 12093
rect 12161 12084 12173 12087
rect 7248 12056 12173 12084
rect 7248 12044 7254 12056
rect 12161 12053 12173 12056
rect 12207 12053 12219 12087
rect 12161 12047 12219 12053
rect 12434 12044 12440 12096
rect 12492 12084 12498 12096
rect 12618 12084 12624 12096
rect 12492 12056 12624 12084
rect 12492 12044 12498 12056
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 13354 12044 13360 12096
rect 13412 12044 13418 12096
rect 13449 12087 13507 12093
rect 13449 12053 13461 12087
rect 13495 12084 13507 12087
rect 16850 12084 16856 12096
rect 13495 12056 16856 12084
rect 13495 12053 13507 12056
rect 13449 12047 13507 12053
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 18156 12084 18184 12124
rect 20349 12121 20361 12124
rect 20395 12121 20407 12155
rect 23934 12152 23940 12164
rect 20349 12115 20407 12121
rect 20732 12124 20838 12152
rect 21652 12124 22140 12152
rect 23782 12124 23940 12152
rect 20732 12096 20760 12124
rect 21652 12096 21680 12124
rect 17368 12056 18184 12084
rect 17368 12044 17374 12056
rect 20714 12044 20720 12096
rect 20772 12084 20778 12096
rect 21634 12084 21640 12096
rect 20772 12056 21640 12084
rect 20772 12044 20778 12056
rect 21634 12044 21640 12056
rect 21692 12044 21698 12096
rect 22112 12084 22140 12124
rect 23860 12084 23888 12124
rect 23934 12112 23940 12124
rect 23992 12112 23998 12164
rect 22112 12056 23888 12084
rect 24026 12044 24032 12096
rect 24084 12044 24090 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 1765 11883 1823 11889
rect 1765 11849 1777 11883
rect 1811 11880 1823 11883
rect 3142 11880 3148 11892
rect 1811 11852 3148 11880
rect 1811 11849 1823 11852
rect 1765 11843 1823 11849
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 4433 11883 4491 11889
rect 4433 11849 4445 11883
rect 4479 11880 4491 11883
rect 4614 11880 4620 11892
rect 4479 11852 4620 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 6549 11883 6607 11889
rect 6549 11849 6561 11883
rect 6595 11880 6607 11883
rect 6914 11880 6920 11892
rect 6595 11852 6920 11880
rect 6595 11849 6607 11852
rect 6549 11843 6607 11849
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 7374 11840 7380 11892
rect 7432 11880 7438 11892
rect 7926 11880 7932 11892
rect 7432 11852 7932 11880
rect 7432 11840 7438 11852
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 8478 11840 8484 11892
rect 8536 11880 8542 11892
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 8536 11852 9137 11880
rect 8536 11840 8542 11852
rect 9125 11849 9137 11852
rect 9171 11849 9183 11883
rect 9125 11843 9183 11849
rect 11974 11840 11980 11892
rect 12032 11840 12038 11892
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 14921 11883 14979 11889
rect 14921 11880 14933 11883
rect 12216 11852 14933 11880
rect 12216 11840 12222 11852
rect 14921 11849 14933 11852
rect 14967 11849 14979 11883
rect 14921 11843 14979 11849
rect 15562 11840 15568 11892
rect 15620 11840 15626 11892
rect 16942 11840 16948 11892
rect 17000 11880 17006 11892
rect 17405 11883 17463 11889
rect 17405 11880 17417 11883
rect 17000 11852 17417 11880
rect 17000 11840 17006 11852
rect 17405 11849 17417 11852
rect 17451 11849 17463 11883
rect 17405 11843 17463 11849
rect 17862 11840 17868 11892
rect 17920 11880 17926 11892
rect 18141 11883 18199 11889
rect 18141 11880 18153 11883
rect 17920 11852 18153 11880
rect 17920 11840 17926 11852
rect 18141 11849 18153 11852
rect 18187 11849 18199 11883
rect 18141 11843 18199 11849
rect 18506 11840 18512 11892
rect 18564 11840 18570 11892
rect 18601 11883 18659 11889
rect 18601 11849 18613 11883
rect 18647 11880 18659 11883
rect 20254 11880 20260 11892
rect 18647 11852 20260 11880
rect 18647 11849 18659 11852
rect 18601 11843 18659 11849
rect 20254 11840 20260 11852
rect 20312 11840 20318 11892
rect 20806 11880 20812 11892
rect 20364 11852 20812 11880
rect 7282 11772 7288 11824
rect 7340 11812 7346 11824
rect 7653 11815 7711 11821
rect 7653 11812 7665 11815
rect 7340 11784 7665 11812
rect 7340 11772 7346 11784
rect 7653 11781 7665 11784
rect 7699 11781 7711 11815
rect 7653 11775 7711 11781
rect 9585 11815 9643 11821
rect 9585 11781 9597 11815
rect 9631 11812 9643 11815
rect 9674 11812 9680 11824
rect 9631 11784 9680 11812
rect 9631 11781 9643 11784
rect 9585 11775 9643 11781
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 12526 11772 12532 11824
rect 12584 11812 12590 11824
rect 16025 11815 16083 11821
rect 12584 11784 13938 11812
rect 12584 11772 12590 11784
rect 16025 11781 16037 11815
rect 16071 11812 16083 11815
rect 20364 11812 20392 11852
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 24026 11880 24032 11892
rect 22112 11852 24032 11880
rect 16071 11784 20392 11812
rect 16071 11781 16083 11784
rect 16025 11775 16083 11781
rect 20714 11772 20720 11824
rect 20772 11772 20778 11824
rect 1946 11704 1952 11756
rect 2004 11704 2010 11756
rect 2130 11704 2136 11756
rect 2188 11704 2194 11756
rect 2406 11704 2412 11756
rect 2464 11704 2470 11756
rect 4338 11704 4344 11756
rect 4396 11704 4402 11756
rect 5442 11704 5448 11756
rect 5500 11704 5506 11756
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 4617 11679 4675 11685
rect 4617 11645 4629 11679
rect 4663 11645 4675 11679
rect 4617 11639 4675 11645
rect 5169 11679 5227 11685
rect 5169 11645 5181 11679
rect 5215 11676 5227 11679
rect 6748 11676 6776 11707
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7190 11744 7196 11756
rect 6972 11716 7196 11744
rect 6972 11704 6978 11716
rect 7190 11704 7196 11716
rect 7248 11704 7254 11756
rect 8754 11704 8760 11756
rect 8812 11704 8818 11756
rect 11146 11704 11152 11756
rect 11204 11704 11210 11756
rect 11974 11704 11980 11756
rect 12032 11744 12038 11756
rect 12158 11744 12164 11756
rect 12032 11716 12164 11744
rect 12032 11704 12038 11716
rect 12158 11704 12164 11716
rect 12216 11704 12222 11756
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11744 12403 11747
rect 12802 11744 12808 11756
rect 12391 11716 12808 11744
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 15930 11704 15936 11756
rect 15988 11704 15994 11756
rect 16114 11704 16120 11756
rect 16172 11744 16178 11756
rect 17313 11747 17371 11753
rect 17313 11744 17325 11747
rect 16172 11716 17325 11744
rect 16172 11704 16178 11716
rect 17313 11713 17325 11716
rect 17359 11744 17371 11747
rect 19058 11744 19064 11756
rect 17359 11716 19064 11744
rect 17359 11713 17371 11716
rect 17313 11707 17371 11713
rect 19058 11704 19064 11716
rect 19116 11704 19122 11756
rect 7282 11676 7288 11688
rect 5215 11648 6684 11676
rect 6748 11648 7288 11676
rect 5215 11645 5227 11648
rect 5169 11639 5227 11645
rect 4632 11608 4660 11639
rect 5718 11608 5724 11620
rect 4632 11580 5724 11608
rect 5718 11568 5724 11580
rect 5776 11568 5782 11620
rect 6656 11608 6684 11648
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 7374 11636 7380 11688
rect 7432 11636 7438 11688
rect 8772 11676 8800 11704
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 7484 11648 8800 11676
rect 9508 11648 10333 11676
rect 7190 11608 7196 11620
rect 6656 11580 7196 11608
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 7484 11608 7512 11648
rect 7300 11580 7512 11608
rect 3694 11500 3700 11552
rect 3752 11540 3758 11552
rect 3973 11543 4031 11549
rect 3973 11540 3985 11543
rect 3752 11512 3985 11540
rect 3752 11500 3758 11512
rect 3973 11509 3985 11512
rect 4019 11509 4031 11543
rect 3973 11503 4031 11509
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 7300 11540 7328 11580
rect 6696 11512 7328 11540
rect 6696 11500 6702 11512
rect 7374 11500 7380 11552
rect 7432 11540 7438 11552
rect 9508 11540 9536 11648
rect 10321 11645 10333 11648
rect 10367 11676 10379 11679
rect 11514 11676 11520 11688
rect 10367 11648 11520 11676
rect 10367 11645 10379 11648
rect 10321 11639 10379 11645
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 11940 11648 12449 11676
rect 11940 11636 11946 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 12529 11679 12587 11685
rect 12529 11645 12541 11679
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11676 13507 11679
rect 15654 11676 15660 11688
rect 13495 11648 15660 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 12544 11608 12572 11639
rect 12216 11580 12572 11608
rect 12216 11568 12222 11580
rect 7432 11512 9536 11540
rect 7432 11500 7438 11512
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 10134 11540 10140 11552
rect 9916 11512 10140 11540
rect 9916 11500 9922 11512
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 12342 11500 12348 11552
rect 12400 11540 12406 11552
rect 13188 11540 13216 11639
rect 15654 11636 15660 11648
rect 15712 11636 15718 11688
rect 16209 11679 16267 11685
rect 16209 11645 16221 11679
rect 16255 11676 16267 11679
rect 17402 11676 17408 11688
rect 16255 11648 17408 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 17402 11636 17408 11648
rect 17460 11636 17466 11688
rect 17497 11679 17555 11685
rect 17497 11645 17509 11679
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 16850 11568 16856 11620
rect 16908 11608 16914 11620
rect 16945 11611 17003 11617
rect 16945 11608 16957 11611
rect 16908 11580 16957 11608
rect 16908 11568 16914 11580
rect 16945 11577 16957 11580
rect 16991 11577 17003 11611
rect 16945 11571 17003 11577
rect 17218 11568 17224 11620
rect 17276 11608 17282 11620
rect 17512 11608 17540 11639
rect 17586 11636 17592 11688
rect 17644 11676 17650 11688
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 17644 11648 18705 11676
rect 17644 11636 17650 11648
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 19702 11636 19708 11688
rect 19760 11636 19766 11688
rect 19981 11679 20039 11685
rect 19981 11645 19993 11679
rect 20027 11676 20039 11679
rect 22112 11676 22140 11852
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 24121 11883 24179 11889
rect 24121 11849 24133 11883
rect 24167 11880 24179 11883
rect 25130 11880 25136 11892
rect 24167 11852 25136 11880
rect 24167 11849 24179 11852
rect 24121 11843 24179 11849
rect 22646 11772 22652 11824
rect 22704 11772 22710 11824
rect 23934 11812 23940 11824
rect 23874 11784 23940 11812
rect 23934 11772 23940 11784
rect 23992 11772 23998 11824
rect 20027 11648 22140 11676
rect 20027 11645 20039 11648
rect 19981 11639 20039 11645
rect 22186 11636 22192 11688
rect 22244 11676 22250 11688
rect 22373 11679 22431 11685
rect 22373 11676 22385 11679
rect 22244 11648 22385 11676
rect 22244 11636 22250 11648
rect 22373 11645 22385 11648
rect 22419 11645 22431 11679
rect 22373 11639 22431 11645
rect 23290 11636 23296 11688
rect 23348 11676 23354 11688
rect 24136 11676 24164 11843
rect 25130 11840 25136 11852
rect 25188 11840 25194 11892
rect 23348 11648 24164 11676
rect 23348 11636 23354 11648
rect 17276 11580 17540 11608
rect 17276 11568 17282 11580
rect 14550 11540 14556 11552
rect 12400 11512 14556 11540
rect 12400 11500 12406 11512
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 14734 11500 14740 11552
rect 14792 11540 14798 11552
rect 17034 11540 17040 11552
rect 14792 11512 17040 11540
rect 14792 11500 14798 11512
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 21450 11500 21456 11552
rect 21508 11500 21514 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 2590 11336 2596 11348
rect 2179 11308 2596 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 5534 11336 5540 11348
rect 4172 11308 5540 11336
rect 2498 11228 2504 11280
rect 2556 11268 2562 11280
rect 3973 11271 4031 11277
rect 3973 11268 3985 11271
rect 2556 11240 3985 11268
rect 2556 11228 2562 11240
rect 3973 11237 3985 11240
rect 4019 11237 4031 11271
rect 3973 11231 4031 11237
rect 2774 11160 2780 11212
rect 2832 11160 2838 11212
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3970 11132 3976 11144
rect 3099 11104 3976 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 4172 11141 4200 11308
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 5776 11308 6561 11336
rect 5776 11296 5782 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 7377 11339 7435 11345
rect 7377 11305 7389 11339
rect 7423 11336 7435 11339
rect 7742 11336 7748 11348
rect 7423 11308 7748 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 7837 11339 7895 11345
rect 7837 11305 7849 11339
rect 7883 11336 7895 11339
rect 10226 11336 10232 11348
rect 7883 11308 10232 11336
rect 7883 11305 7895 11308
rect 7837 11299 7895 11305
rect 10226 11296 10232 11308
rect 10284 11296 10290 11348
rect 10321 11339 10379 11345
rect 10321 11305 10333 11339
rect 10367 11336 10379 11339
rect 11882 11336 11888 11348
rect 10367 11308 11888 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 12250 11296 12256 11348
rect 12308 11336 12314 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 12308 11308 13277 11336
rect 12308 11296 12314 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 14792 11308 16436 11336
rect 14792 11296 14798 11308
rect 6638 11228 6644 11280
rect 6696 11268 6702 11280
rect 9125 11271 9183 11277
rect 6696 11240 8616 11268
rect 6696 11228 6702 11240
rect 4798 11160 4804 11212
rect 4856 11160 4862 11212
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5810 11200 5816 11212
rect 5123 11172 5816 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 7834 11160 7840 11212
rect 7892 11200 7898 11212
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 7892 11172 8309 11200
rect 7892 11160 7898 11172
rect 8297 11169 8309 11172
rect 8343 11169 8355 11203
rect 8297 11163 8355 11169
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11169 8539 11203
rect 8588 11200 8616 11240
rect 9125 11237 9137 11271
rect 9171 11268 9183 11271
rect 9306 11268 9312 11280
rect 9171 11240 9312 11268
rect 9171 11237 9183 11240
rect 9125 11231 9183 11237
rect 9306 11228 9312 11240
rect 9364 11228 9370 11280
rect 9416 11240 10732 11268
rect 9416 11200 9444 11240
rect 8588 11172 9444 11200
rect 8481 11163 8539 11169
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 8386 11132 8392 11144
rect 8251 11104 8392 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 6546 11064 6552 11076
rect 6302 11036 6552 11064
rect 6546 11024 6552 11036
rect 6604 11024 6610 11076
rect 7282 10956 7288 11008
rect 7340 10996 7346 11008
rect 8496 10996 8524 11163
rect 9674 11160 9680 11212
rect 9732 11160 9738 11212
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9493 11135 9551 11141
rect 9493 11132 9505 11135
rect 9272 11104 9505 11132
rect 9272 11092 9278 11104
rect 9493 11101 9505 11104
rect 9539 11101 9551 11135
rect 9493 11095 9551 11101
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11132 9643 11135
rect 9631 11104 10640 11132
rect 9631 11101 9643 11104
rect 9585 11095 9643 11101
rect 10134 10996 10140 11008
rect 7340 10968 10140 10996
rect 7340 10956 7346 10968
rect 10134 10956 10140 10968
rect 10192 10956 10198 11008
rect 10612 10996 10640 11104
rect 10704 11073 10732 11240
rect 11146 11228 11152 11280
rect 11204 11268 11210 11280
rect 16408 11268 16436 11308
rect 16482 11296 16488 11348
rect 16540 11296 16546 11348
rect 17386 11339 17444 11345
rect 17386 11336 17398 11339
rect 17236 11308 17398 11336
rect 17236 11268 17264 11308
rect 17386 11305 17398 11308
rect 17432 11336 17444 11339
rect 18782 11336 18788 11348
rect 17432 11308 18788 11336
rect 17432 11305 17444 11308
rect 17386 11299 17444 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 18874 11296 18880 11348
rect 18932 11296 18938 11348
rect 11204 11240 11652 11268
rect 16408 11240 17264 11268
rect 11204 11228 11210 11240
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 11011 11172 11468 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 10689 11067 10747 11073
rect 10689 11033 10701 11067
rect 10735 11033 10747 11067
rect 10689 11027 10747 11033
rect 10778 11024 10784 11076
rect 10836 11024 10842 11076
rect 11054 11064 11060 11076
rect 10888 11036 11060 11064
rect 10888 10996 10916 11036
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 10612 10968 10916 10996
rect 11440 10996 11468 11172
rect 11514 11160 11520 11212
rect 11572 11160 11578 11212
rect 11624 11200 11652 11240
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 11624 11172 11805 11200
rect 11793 11169 11805 11172
rect 11839 11200 11851 11203
rect 12250 11200 12256 11212
rect 11839 11172 12256 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 14550 11160 14556 11212
rect 14608 11200 14614 11212
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 14608 11172 14749 11200
rect 14608 11160 14614 11172
rect 14737 11169 14749 11172
rect 14783 11200 14795 11203
rect 15102 11200 15108 11212
rect 14783 11172 15108 11200
rect 14783 11169 14795 11172
rect 14737 11163 14795 11169
rect 15102 11160 15108 11172
rect 15160 11160 15166 11212
rect 22646 11160 22652 11212
rect 22704 11160 22710 11212
rect 26878 11160 26884 11212
rect 26936 11200 26942 11212
rect 29733 11203 29791 11209
rect 29733 11200 29745 11203
rect 26936 11172 29745 11200
rect 26936 11160 26942 11172
rect 29733 11169 29745 11172
rect 29779 11169 29791 11203
rect 29733 11163 29791 11169
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 16908 11104 17141 11132
rect 16908 11092 16914 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 19150 11092 19156 11144
rect 19208 11132 19214 11144
rect 19521 11135 19579 11141
rect 19521 11132 19533 11135
rect 19208 11104 19533 11132
rect 19208 11092 19214 11104
rect 19521 11101 19533 11104
rect 19567 11101 19579 11135
rect 20901 11135 20959 11141
rect 20901 11132 20913 11135
rect 19521 11095 19579 11101
rect 20272 11104 20913 11132
rect 11882 11024 11888 11076
rect 11940 11064 11946 11076
rect 11940 11036 12112 11064
rect 11940 11024 11946 11036
rect 11974 10996 11980 11008
rect 11440 10968 11980 10996
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 12084 10996 12112 11036
rect 12526 11024 12532 11076
rect 12584 11024 12590 11076
rect 15010 11024 15016 11076
rect 15068 11024 15074 11076
rect 15286 11024 15292 11076
rect 15344 11064 15350 11076
rect 15344 11036 15502 11064
rect 15344 11024 15350 11036
rect 17862 11024 17868 11076
rect 17920 11024 17926 11076
rect 19702 11024 19708 11076
rect 19760 11064 19766 11076
rect 20272 11073 20300 11104
rect 20901 11101 20913 11104
rect 20947 11101 20959 11135
rect 20901 11095 20959 11101
rect 20257 11067 20315 11073
rect 20257 11064 20269 11067
rect 19760 11036 20269 11064
rect 19760 11024 19766 11036
rect 20257 11033 20269 11036
rect 20303 11033 20315 11067
rect 20257 11027 20315 11033
rect 21174 11024 21180 11076
rect 21232 11024 21238 11076
rect 21284 11036 21666 11064
rect 15194 10996 15200 11008
rect 12084 10968 15200 10996
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 15654 10956 15660 11008
rect 15712 10996 15718 11008
rect 19334 10996 19340 11008
rect 15712 10968 19340 10996
rect 15712 10956 15718 10968
rect 19334 10956 19340 10968
rect 19392 10956 19398 11008
rect 20714 10956 20720 11008
rect 20772 10996 20778 11008
rect 21284 10996 21312 11036
rect 28350 11024 28356 11076
rect 28408 11064 28414 11076
rect 30009 11067 30067 11073
rect 30009 11064 30021 11067
rect 28408 11036 30021 11064
rect 28408 11024 28414 11036
rect 30009 11033 30021 11036
rect 30055 11033 30067 11067
rect 30009 11027 30067 11033
rect 30098 11024 30104 11076
rect 30156 11064 30162 11076
rect 30156 11036 30498 11064
rect 30156 11024 30162 11036
rect 31662 11024 31668 11076
rect 31720 11064 31726 11076
rect 31757 11067 31815 11073
rect 31757 11064 31769 11067
rect 31720 11036 31769 11064
rect 31720 11024 31726 11036
rect 31757 11033 31769 11036
rect 31803 11064 31815 11067
rect 47854 11064 47860 11076
rect 31803 11036 47860 11064
rect 31803 11033 31815 11036
rect 31757 11027 31815 11033
rect 47854 11024 47860 11036
rect 47912 11024 47918 11076
rect 20772 10968 21312 10996
rect 20772 10956 20778 10968
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 3878 10752 3884 10804
rect 3936 10752 3942 10804
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 5261 10795 5319 10801
rect 5261 10792 5273 10795
rect 4396 10764 5273 10792
rect 4396 10752 4402 10764
rect 5261 10761 5273 10764
rect 5307 10761 5319 10795
rect 5261 10755 5319 10761
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 6972 10764 7144 10792
rect 6972 10752 6978 10764
rect 4246 10684 4252 10736
rect 4304 10724 4310 10736
rect 4304 10696 4660 10724
rect 4304 10684 4310 10696
rect 2038 10616 2044 10668
rect 2096 10616 2102 10668
rect 2314 10616 2320 10668
rect 2372 10616 2378 10668
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10656 3847 10659
rect 4430 10656 4436 10668
rect 3835 10628 4436 10656
rect 3835 10625 3847 10628
rect 3789 10619 3847 10625
rect 4430 10616 4436 10628
rect 4488 10616 4494 10668
rect 4522 10616 4528 10668
rect 4580 10616 4586 10668
rect 4632 10656 4660 10696
rect 4706 10684 4712 10736
rect 4764 10684 4770 10736
rect 7116 10724 7144 10764
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 7248 10764 10333 10792
rect 7248 10752 7254 10764
rect 10321 10761 10333 10764
rect 10367 10761 10379 10795
rect 10321 10755 10379 10761
rect 11514 10752 11520 10804
rect 11572 10792 11578 10804
rect 12158 10792 12164 10804
rect 11572 10764 12164 10792
rect 11572 10752 11578 10764
rect 12158 10752 12164 10764
rect 12216 10792 12222 10804
rect 13817 10795 13875 10801
rect 13817 10792 13829 10795
rect 12216 10764 13829 10792
rect 12216 10752 12222 10764
rect 13817 10761 13829 10764
rect 13863 10761 13875 10795
rect 13817 10755 13875 10761
rect 14369 10795 14427 10801
rect 14369 10761 14381 10795
rect 14415 10792 14427 10795
rect 15562 10792 15568 10804
rect 14415 10764 15568 10792
rect 14415 10761 14427 10764
rect 14369 10755 14427 10761
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 15933 10795 15991 10801
rect 15933 10792 15945 10795
rect 15856 10764 15945 10792
rect 4816 10696 6960 10724
rect 7116 10696 7236 10724
rect 4816 10656 4844 10696
rect 4632 10628 4844 10656
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 6932 10665 6960 10696
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5316 10628 5641 10656
rect 5316 10616 5322 10628
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 5736 10520 5764 10551
rect 5902 10548 5908 10600
rect 5960 10548 5966 10600
rect 6914 10520 6920 10532
rect 5736 10492 6920 10520
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 6730 10412 6736 10464
rect 6788 10412 6794 10464
rect 7208 10452 7236 10696
rect 9398 10684 9404 10736
rect 9456 10684 9462 10736
rect 12342 10724 12348 10736
rect 12084 10696 12348 10724
rect 8754 10616 8760 10668
rect 8812 10616 8818 10668
rect 9582 10616 9588 10668
rect 9640 10656 9646 10668
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 9640 10628 10701 10656
rect 9640 10616 9646 10628
rect 10689 10625 10701 10628
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 12084 10665 12112 10696
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 12618 10684 12624 10736
rect 12676 10724 12682 10736
rect 14737 10727 14795 10733
rect 12676 10696 12834 10724
rect 12676 10684 12682 10696
rect 14737 10693 14749 10727
rect 14783 10724 14795 10727
rect 15746 10724 15752 10736
rect 14783 10696 15752 10724
rect 14783 10693 14795 10696
rect 14737 10687 14795 10693
rect 15746 10684 15752 10696
rect 15804 10684 15810 10736
rect 12069 10659 12127 10665
rect 12069 10656 12081 10659
rect 11296 10628 12081 10656
rect 11296 10616 11302 10628
rect 12069 10625 12081 10628
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 14274 10616 14280 10668
rect 14332 10656 14338 10668
rect 15856 10656 15884 10764
rect 15933 10761 15945 10764
rect 15979 10761 15991 10795
rect 15933 10755 15991 10761
rect 17402 10752 17408 10804
rect 17460 10792 17466 10804
rect 19245 10795 19303 10801
rect 19245 10792 19257 10795
rect 17460 10764 19257 10792
rect 17460 10752 17466 10764
rect 19245 10761 19257 10764
rect 19291 10761 19303 10795
rect 21450 10792 21456 10804
rect 19245 10755 19303 10761
rect 19536 10764 21456 10792
rect 17862 10684 17868 10736
rect 17920 10724 17926 10736
rect 17920 10696 18262 10724
rect 17920 10684 17926 10696
rect 14332 10628 15884 10656
rect 15948 10628 16712 10656
rect 14332 10616 14338 10628
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 7653 10591 7711 10597
rect 7432 10560 7512 10588
rect 7432 10548 7438 10560
rect 7374 10452 7380 10464
rect 7208 10424 7380 10452
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7484 10452 7512 10560
rect 7653 10557 7665 10591
rect 7699 10588 7711 10591
rect 7699 10560 9076 10588
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 9048 10520 9076 10560
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10376 10560 10793 10588
rect 10376 10548 10382 10560
rect 10781 10557 10793 10560
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 10965 10591 11023 10597
rect 10965 10557 10977 10591
rect 11011 10588 11023 10591
rect 11146 10588 11152 10600
rect 11011 10560 11152 10588
rect 11011 10557 11023 10560
rect 10965 10551 11023 10557
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 14829 10591 14887 10597
rect 14829 10588 14841 10591
rect 11900 10560 14841 10588
rect 9674 10520 9680 10532
rect 9048 10492 9680 10520
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 7834 10452 7840 10464
rect 7484 10424 7840 10452
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 8018 10412 8024 10464
rect 8076 10452 8082 10464
rect 11900 10452 11928 10560
rect 14829 10557 14841 10560
rect 14875 10557 14887 10591
rect 14829 10551 14887 10557
rect 14921 10591 14979 10597
rect 14921 10557 14933 10591
rect 14967 10588 14979 10591
rect 15948 10588 15976 10628
rect 14967 10560 15976 10588
rect 16025 10591 16083 10597
rect 14967 10557 14979 10560
rect 14921 10551 14979 10557
rect 16025 10557 16037 10591
rect 16071 10588 16083 10591
rect 16209 10591 16267 10597
rect 16071 10560 16160 10588
rect 16071 10557 16083 10560
rect 16025 10551 16083 10557
rect 15565 10523 15623 10529
rect 15565 10489 15577 10523
rect 15611 10520 15623 10523
rect 15654 10520 15660 10532
rect 15611 10492 15660 10520
rect 15611 10489 15623 10492
rect 15565 10483 15623 10489
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 8076 10424 11928 10452
rect 8076 10412 8082 10424
rect 11974 10412 11980 10464
rect 12032 10452 12038 10464
rect 12326 10455 12384 10461
rect 12326 10452 12338 10455
rect 12032 10424 12338 10452
rect 12032 10412 12038 10424
rect 12326 10421 12338 10424
rect 12372 10421 12384 10455
rect 12326 10415 12384 10421
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 16022 10452 16028 10464
rect 15252 10424 16028 10452
rect 15252 10412 15258 10424
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 16132 10452 16160 10560
rect 16209 10557 16221 10591
rect 16255 10588 16267 10591
rect 16298 10588 16304 10600
rect 16255 10560 16304 10588
rect 16255 10557 16267 10560
rect 16209 10551 16267 10557
rect 16298 10548 16304 10560
rect 16356 10548 16362 10600
rect 16684 10588 16712 10628
rect 17034 10616 17040 10668
rect 17092 10616 17098 10668
rect 17494 10616 17500 10668
rect 17552 10616 17558 10668
rect 17310 10588 17316 10600
rect 16684 10560 17316 10588
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 17773 10591 17831 10597
rect 17773 10588 17785 10591
rect 17604 10560 17785 10588
rect 17034 10480 17040 10532
rect 17092 10520 17098 10532
rect 17604 10520 17632 10560
rect 17773 10557 17785 10560
rect 17819 10588 17831 10591
rect 19536 10588 19564 10764
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 20714 10684 20720 10736
rect 20772 10684 20778 10736
rect 17819 10560 19564 10588
rect 17819 10557 17831 10560
rect 17773 10551 17831 10557
rect 19702 10548 19708 10600
rect 19760 10548 19766 10600
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 22646 10588 22652 10600
rect 20027 10560 22652 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 22646 10548 22652 10560
rect 22704 10548 22710 10600
rect 17092 10492 17632 10520
rect 17092 10480 17098 10492
rect 18782 10480 18788 10532
rect 18840 10520 18846 10532
rect 18840 10492 19564 10520
rect 18840 10480 18846 10492
rect 19426 10452 19432 10464
rect 16132 10424 19432 10452
rect 19426 10412 19432 10424
rect 19484 10412 19490 10464
rect 19536 10452 19564 10492
rect 21453 10455 21511 10461
rect 21453 10452 21465 10455
rect 19536 10424 21465 10452
rect 21453 10421 21465 10424
rect 21499 10421 21511 10455
rect 21453 10415 21511 10421
rect 24854 10412 24860 10464
rect 24912 10452 24918 10464
rect 32858 10452 32864 10464
rect 24912 10424 32864 10452
rect 24912 10412 24918 10424
rect 32858 10412 32864 10424
rect 32916 10412 32922 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 5997 10251 6055 10257
rect 5997 10217 6009 10251
rect 6043 10248 6055 10251
rect 9585 10251 9643 10257
rect 6043 10220 9168 10248
rect 6043 10217 6055 10220
rect 5997 10211 6055 10217
rect 1118 10140 1124 10192
rect 1176 10180 1182 10192
rect 1176 10152 2774 10180
rect 1176 10140 1182 10152
rect 934 10072 940 10124
rect 992 10112 998 10124
rect 1581 10115 1639 10121
rect 1581 10112 1593 10115
rect 992 10084 1593 10112
rect 992 10072 998 10084
rect 1581 10081 1593 10084
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10112 1915 10115
rect 2222 10112 2228 10124
rect 1903 10084 2228 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 2222 10072 2228 10084
rect 2280 10072 2286 10124
rect 2746 10112 2774 10152
rect 4801 10115 4859 10121
rect 4801 10112 4813 10115
rect 2746 10084 4813 10112
rect 4801 10081 4813 10084
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 7834 10112 7840 10124
rect 6871 10084 7840 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 2832 10016 3065 10044
rect 2832 10004 2838 10016
rect 3053 10013 3065 10016
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 6454 10044 6460 10056
rect 4571 10016 6460 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 2869 9911 2927 9917
rect 2869 9877 2881 9911
rect 2915 9908 2927 9911
rect 4540 9908 4568 10007
rect 6454 10004 6460 10016
rect 6512 10004 6518 10056
rect 8754 10044 8760 10056
rect 8234 10016 8760 10044
rect 8754 10004 8760 10016
rect 8812 10044 8818 10056
rect 9030 10044 9036 10056
rect 8812 10016 9036 10044
rect 8812 10004 8818 10016
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 9140 10044 9168 10220
rect 9585 10217 9597 10251
rect 9631 10248 9643 10251
rect 9631 10220 12756 10248
rect 9631 10217 9643 10220
rect 9585 10211 9643 10217
rect 12728 10180 12756 10220
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 13633 10251 13691 10257
rect 13633 10248 13645 10251
rect 12860 10220 13645 10248
rect 12860 10208 12866 10220
rect 13633 10217 13645 10220
rect 13679 10217 13691 10251
rect 15010 10248 15016 10260
rect 13633 10211 13691 10217
rect 14476 10220 15016 10248
rect 14182 10180 14188 10192
rect 12728 10152 14188 10180
rect 14182 10140 14188 10152
rect 14240 10140 14246 10192
rect 10502 10072 10508 10124
rect 10560 10072 10566 10124
rect 10597 10115 10655 10121
rect 10597 10081 10609 10115
rect 10643 10081 10655 10115
rect 10597 10075 10655 10081
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 9140 10016 10425 10044
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 7101 9979 7159 9985
rect 7101 9945 7113 9979
rect 7147 9976 7159 9979
rect 7190 9976 7196 9988
rect 7147 9948 7196 9976
rect 7147 9945 7159 9948
rect 7101 9939 7159 9945
rect 7190 9936 7196 9948
rect 7248 9936 7254 9988
rect 8386 9936 8392 9988
rect 8444 9976 8450 9988
rect 9490 9976 9496 9988
rect 8444 9948 9496 9976
rect 8444 9936 8450 9948
rect 9490 9936 9496 9948
rect 9548 9976 9554 9988
rect 10612 9976 10640 10075
rect 11238 10072 11244 10124
rect 11296 10072 11302 10124
rect 11514 10072 11520 10124
rect 11572 10072 11578 10124
rect 12250 10072 12256 10124
rect 12308 10112 12314 10124
rect 12894 10112 12900 10124
rect 12308 10084 12900 10112
rect 12308 10072 12314 10084
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 13004 10044 13032 10075
rect 13078 10072 13084 10124
rect 13136 10112 13142 10124
rect 14476 10112 14504 10220
rect 15010 10208 15016 10220
rect 15068 10248 15074 10260
rect 16301 10251 16359 10257
rect 16301 10248 16313 10251
rect 15068 10220 16313 10248
rect 15068 10208 15074 10220
rect 16301 10217 16313 10220
rect 16347 10248 16359 10251
rect 17586 10248 17592 10260
rect 16347 10220 17592 10248
rect 16347 10217 16359 10220
rect 16301 10211 16359 10217
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 18877 10251 18935 10257
rect 18877 10217 18889 10251
rect 18923 10248 18935 10251
rect 19242 10248 19248 10260
rect 18923 10220 19248 10248
rect 18923 10217 18935 10220
rect 18877 10211 18935 10217
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 23290 10248 23296 10260
rect 21652 10220 23296 10248
rect 15838 10140 15844 10192
rect 15896 10180 15902 10192
rect 16942 10180 16948 10192
rect 15896 10152 16948 10180
rect 15896 10140 15902 10152
rect 16942 10140 16948 10152
rect 17000 10140 17006 10192
rect 13136 10084 14504 10112
rect 13136 10072 13142 10084
rect 14550 10072 14556 10124
rect 14608 10072 14614 10124
rect 14826 10072 14832 10124
rect 14884 10072 14890 10124
rect 14918 10072 14924 10124
rect 14976 10112 14982 10124
rect 17034 10112 17040 10124
rect 14976 10084 17040 10112
rect 14976 10072 14982 10084
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 19429 10115 19487 10121
rect 19429 10112 19441 10115
rect 17144 10084 19441 10112
rect 13170 10044 13176 10056
rect 12676 10016 12940 10044
rect 13004 10016 13176 10044
rect 12676 10004 12682 10016
rect 9548 9948 10640 9976
rect 12912 9976 12940 10016
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 17144 10053 17172 10084
rect 19429 10081 19441 10084
rect 19475 10112 19487 10115
rect 19702 10112 19708 10124
rect 19475 10084 19708 10112
rect 19475 10081 19487 10084
rect 19429 10075 19487 10081
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16908 10016 17141 10044
rect 16908 10004 16914 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 13446 9976 13452 9988
rect 12912 9948 13452 9976
rect 9548 9936 9554 9948
rect 13446 9936 13452 9948
rect 13504 9936 13510 9988
rect 14734 9976 14740 9988
rect 13648 9948 14740 9976
rect 2915 9880 4568 9908
rect 2915 9877 2927 9880
rect 2869 9871 2927 9877
rect 6730 9868 6736 9920
rect 6788 9908 6794 9920
rect 8478 9908 8484 9920
rect 6788 9880 8484 9908
rect 6788 9868 6794 9880
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 8573 9911 8631 9917
rect 8573 9877 8585 9911
rect 8619 9908 8631 9911
rect 9674 9908 9680 9920
rect 8619 9880 9680 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 10042 9868 10048 9920
rect 10100 9868 10106 9920
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 13648 9908 13676 9948
rect 14734 9936 14740 9948
rect 14792 9936 14798 9988
rect 15286 9936 15292 9988
rect 15344 9936 15350 9988
rect 16224 9948 17356 9976
rect 12400 9880 13676 9908
rect 12400 9868 12406 9880
rect 13722 9868 13728 9920
rect 13780 9908 13786 9920
rect 16224 9908 16252 9948
rect 13780 9880 16252 9908
rect 17328 9908 17356 9948
rect 17402 9936 17408 9988
rect 17460 9936 17466 9988
rect 17862 9936 17868 9988
rect 17920 9936 17926 9988
rect 19705 9979 19763 9985
rect 19705 9976 19717 9979
rect 18800 9948 19717 9976
rect 18800 9908 18828 9948
rect 19705 9945 19717 9948
rect 19751 9945 19763 9979
rect 19705 9939 19763 9945
rect 17328 9880 18828 9908
rect 19720 9908 19748 9939
rect 20714 9936 20720 9988
rect 20772 9936 20778 9988
rect 21652 9985 21680 10220
rect 23290 10208 23296 10220
rect 23348 10208 23354 10260
rect 22094 10072 22100 10124
rect 22152 10112 22158 10124
rect 23842 10112 23848 10124
rect 22152 10084 23848 10112
rect 22152 10072 22158 10084
rect 23842 10072 23848 10084
rect 23900 10072 23906 10124
rect 21637 9979 21695 9985
rect 21637 9976 21649 9979
rect 21008 9948 21649 9976
rect 21008 9908 21036 9948
rect 21637 9945 21649 9948
rect 21683 9945 21695 9979
rect 21637 9939 21695 9945
rect 19720 9880 21036 9908
rect 13780 9868 13786 9880
rect 21174 9868 21180 9920
rect 21232 9868 21238 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 6914 9664 6920 9716
rect 6972 9664 6978 9716
rect 9858 9704 9864 9716
rect 9692 9676 9864 9704
rect 4893 9639 4951 9645
rect 4893 9636 4905 9639
rect 4356 9608 4905 9636
rect 1578 9528 1584 9580
rect 1636 9528 1642 9580
rect 3329 9571 3387 9577
rect 3329 9537 3341 9571
rect 3375 9568 3387 9571
rect 3418 9568 3424 9580
rect 3375 9540 3424 9568
rect 3375 9537 3387 9540
rect 3329 9531 3387 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 4356 9577 4384 9608
rect 4893 9605 4905 9608
rect 4939 9636 4951 9639
rect 6086 9636 6092 9648
rect 4939 9608 6092 9636
rect 4939 9605 4951 9608
rect 4893 9599 4951 9605
rect 6086 9596 6092 9608
rect 6144 9596 6150 9648
rect 6270 9596 6276 9648
rect 6328 9636 6334 9648
rect 6328 9608 7512 9636
rect 6328 9596 6334 9608
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9537 4399 9571
rect 4341 9531 4399 9537
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9568 5411 9571
rect 5626 9568 5632 9580
rect 5399 9540 5632 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9568 6055 9571
rect 7006 9568 7012 9580
rect 6043 9540 7012 9568
rect 6043 9537 6055 9540
rect 5997 9531 6055 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9500 1915 9503
rect 5902 9500 5908 9512
rect 1903 9472 5908 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 6730 9460 6736 9512
rect 6788 9500 6794 9512
rect 7300 9500 7328 9531
rect 7484 9509 7512 9608
rect 8386 9596 8392 9648
rect 8444 9596 8450 9648
rect 9030 9596 9036 9648
rect 9088 9596 9094 9648
rect 9692 9568 9720 9676
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 10318 9664 10324 9716
rect 10376 9664 10382 9716
rect 12158 9664 12164 9716
rect 12216 9704 12222 9716
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 12216 9676 13461 9704
rect 12216 9664 12222 9676
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 13449 9667 13507 9673
rect 15120 9676 16068 9704
rect 10778 9596 10784 9648
rect 10836 9596 10842 9648
rect 15120 9636 15148 9676
rect 14384 9608 15148 9636
rect 16040 9636 16068 9676
rect 17218 9636 17224 9648
rect 16040 9608 17224 9636
rect 9600 9540 9720 9568
rect 6788 9472 7328 9500
rect 7377 9503 7435 9509
rect 6788 9460 6794 9472
rect 7377 9469 7389 9503
rect 7423 9469 7435 9503
rect 7377 9463 7435 9469
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9469 7527 9503
rect 7469 9463 7527 9469
rect 3145 9435 3203 9441
rect 3145 9401 3157 9435
rect 3191 9432 3203 9435
rect 3786 9432 3792 9444
rect 3191 9404 3792 9432
rect 3191 9401 3203 9404
rect 3145 9395 3203 9401
rect 3786 9392 3792 9404
rect 3844 9392 3850 9444
rect 7392 9432 7420 9463
rect 7834 9460 7840 9512
rect 7892 9500 7898 9512
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 7892 9472 8125 9500
rect 7892 9460 7898 9472
rect 8113 9469 8125 9472
rect 8159 9469 8171 9503
rect 9600 9500 9628 9540
rect 9858 9528 9864 9580
rect 9916 9568 9922 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 9916 9540 10701 9568
rect 9916 9528 9922 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 11238 9528 11244 9580
rect 11296 9568 11302 9580
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11296 9540 11713 9568
rect 11296 9528 11302 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 13446 9568 13452 9580
rect 13110 9540 13452 9568
rect 11701 9531 11759 9537
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 8113 9463 8171 9469
rect 8220 9472 9628 9500
rect 10965 9503 11023 9509
rect 8220 9432 8248 9472
rect 10965 9469 10977 9503
rect 11011 9500 11023 9503
rect 11977 9503 12035 9509
rect 11977 9500 11989 9503
rect 11011 9472 11989 9500
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 11977 9469 11989 9472
rect 12023 9500 12035 9503
rect 13170 9500 13176 9512
rect 12023 9472 13176 9500
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 13630 9460 13636 9512
rect 13688 9500 13694 9512
rect 14384 9500 14412 9608
rect 17218 9596 17224 9608
rect 17276 9636 17282 9648
rect 17402 9636 17408 9648
rect 17276 9608 17408 9636
rect 17276 9596 17282 9608
rect 17402 9596 17408 9608
rect 17460 9596 17466 9648
rect 18414 9636 18420 9648
rect 18354 9608 18420 9636
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 19521 9639 19579 9645
rect 19521 9605 19533 9639
rect 19567 9636 19579 9639
rect 23566 9636 23572 9648
rect 19567 9608 23572 9636
rect 19567 9605 19579 9608
rect 19521 9599 19579 9605
rect 23566 9596 23572 9608
rect 23624 9596 23630 9648
rect 14458 9528 14464 9580
rect 14516 9528 14522 9580
rect 16114 9568 16120 9580
rect 15870 9540 16120 9568
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 19426 9528 19432 9580
rect 19484 9528 19490 9580
rect 27430 9528 27436 9580
rect 27488 9568 27494 9580
rect 27525 9571 27583 9577
rect 27525 9568 27537 9571
rect 27488 9540 27537 9568
rect 27488 9528 27494 9540
rect 27525 9537 27537 9540
rect 27571 9537 27583 9571
rect 27525 9531 27583 9537
rect 14737 9503 14795 9509
rect 14737 9500 14749 9503
rect 13688 9472 14749 9500
rect 13688 9460 13694 9472
rect 14737 9469 14749 9472
rect 14783 9469 14795 9503
rect 14737 9463 14795 9469
rect 14826 9460 14832 9512
rect 14884 9500 14890 9512
rect 16209 9503 16267 9509
rect 16209 9500 16221 9503
rect 14884 9472 16221 9500
rect 14884 9460 14890 9472
rect 16209 9469 16221 9472
rect 16255 9469 16267 9503
rect 16209 9463 16267 9469
rect 16850 9460 16856 9512
rect 16908 9460 16914 9512
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9500 17187 9503
rect 18322 9500 18328 9512
rect 17175 9472 18328 9500
rect 17175 9469 17187 9472
rect 17129 9463 17187 9469
rect 18322 9460 18328 9472
rect 18380 9500 18386 9512
rect 19242 9500 19248 9512
rect 18380 9472 19248 9500
rect 18380 9460 18386 9472
rect 19242 9460 19248 9472
rect 19300 9460 19306 9512
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 21174 9500 21180 9512
rect 19751 9472 21180 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 21174 9460 21180 9472
rect 21232 9460 21238 9512
rect 22554 9460 22560 9512
rect 22612 9500 22618 9512
rect 27985 9503 28043 9509
rect 27985 9500 27997 9503
rect 22612 9472 27997 9500
rect 22612 9460 22618 9472
rect 27985 9469 27997 9472
rect 28031 9469 28043 9503
rect 27985 9463 28043 9469
rect 11422 9432 11428 9444
rect 7392 9404 8248 9432
rect 9784 9404 11428 9432
rect 3053 9367 3111 9373
rect 3053 9333 3065 9367
rect 3099 9364 3111 9367
rect 3697 9367 3755 9373
rect 3697 9364 3709 9367
rect 3099 9336 3709 9364
rect 3099 9333 3111 9336
rect 3053 9327 3111 9333
rect 3697 9333 3709 9336
rect 3743 9364 3755 9367
rect 9784 9364 9812 9404
rect 11422 9392 11428 9404
rect 11480 9392 11486 9444
rect 19061 9435 19119 9441
rect 19061 9401 19073 9435
rect 19107 9432 19119 9435
rect 19610 9432 19616 9444
rect 19107 9404 19616 9432
rect 19107 9401 19119 9404
rect 19061 9395 19119 9401
rect 19610 9392 19616 9404
rect 19668 9392 19674 9444
rect 3743 9336 9812 9364
rect 9861 9367 9919 9373
rect 3743 9333 3755 9336
rect 3697 9327 3755 9333
rect 9861 9333 9873 9367
rect 9907 9364 9919 9367
rect 10134 9364 10140 9376
rect 9907 9336 10140 9364
rect 9907 9333 9919 9336
rect 9861 9327 9919 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10318 9324 10324 9376
rect 10376 9364 10382 9376
rect 14734 9364 14740 9376
rect 10376 9336 14740 9364
rect 10376 9324 10382 9336
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 18601 9367 18659 9373
rect 18601 9364 18613 9367
rect 16356 9336 18613 9364
rect 16356 9324 16362 9336
rect 18601 9333 18613 9336
rect 18647 9333 18659 9367
rect 18601 9327 18659 9333
rect 27801 9367 27859 9373
rect 27801 9333 27813 9367
rect 27847 9364 27859 9367
rect 31662 9364 31668 9376
rect 27847 9336 31668 9364
rect 27847 9333 27859 9336
rect 27801 9327 27859 9333
rect 31662 9324 31668 9336
rect 31720 9324 31726 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9160 4031 9163
rect 4062 9160 4068 9172
rect 4019 9132 4068 9160
rect 4019 9129 4031 9132
rect 3973 9123 4031 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 5166 9120 5172 9172
rect 5224 9120 5230 9172
rect 6822 9120 6828 9172
rect 6880 9120 6886 9172
rect 7024 9132 22094 9160
rect 4522 9052 4528 9104
rect 4580 9092 4586 9104
rect 6181 9095 6239 9101
rect 6181 9092 6193 9095
rect 4580 9064 6193 9092
rect 4580 9052 4586 9064
rect 6181 9061 6193 9064
rect 6227 9061 6239 9095
rect 6181 9055 6239 9061
rect 1854 8984 1860 9036
rect 1912 8984 1918 9036
rect 4982 8984 4988 9036
rect 5040 9024 5046 9036
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 5040 8996 5733 9024
rect 5040 8984 5046 8996
rect 5721 8993 5733 8996
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 992 8928 1593 8956
rect 992 8916 998 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 3326 8956 3332 8968
rect 3099 8928 3332 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 5368 8888 5396 8919
rect 6362 8916 6368 8968
rect 6420 8916 6426 8968
rect 7024 8965 7052 9132
rect 22066 9104 22094 9132
rect 8386 9052 8392 9104
rect 8444 9092 8450 9104
rect 9858 9092 9864 9104
rect 8444 9064 9864 9092
rect 8444 9052 8450 9064
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 10413 9095 10471 9101
rect 10413 9061 10425 9095
rect 10459 9092 10471 9095
rect 12805 9095 12863 9101
rect 10459 9064 12434 9092
rect 10459 9061 10471 9064
rect 10413 9055 10471 9061
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7745 9027 7803 9033
rect 7745 9024 7757 9027
rect 7156 8996 7757 9024
rect 7156 8984 7162 8996
rect 7745 8993 7757 8996
rect 7791 8993 7803 9027
rect 7745 8987 7803 8993
rect 9122 8984 9128 9036
rect 9180 8984 9186 9036
rect 9398 8984 9404 9036
rect 9456 8984 9462 9036
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 9732 8996 10977 9024
rect 9732 8984 9738 8996
rect 10965 8993 10977 8996
rect 11011 8993 11023 9027
rect 10965 8987 11023 8993
rect 12250 8984 12256 9036
rect 12308 8984 12314 9036
rect 12406 9024 12434 9064
rect 12805 9061 12817 9095
rect 12851 9092 12863 9095
rect 15470 9092 15476 9104
rect 12851 9064 15476 9092
rect 12851 9061 12863 9064
rect 12805 9055 12863 9061
rect 15470 9052 15476 9064
rect 15528 9052 15534 9104
rect 17402 9052 17408 9104
rect 17460 9092 17466 9104
rect 17773 9095 17831 9101
rect 17773 9092 17785 9095
rect 17460 9064 17785 9092
rect 17460 9052 17466 9064
rect 17773 9061 17785 9064
rect 17819 9061 17831 9095
rect 22066 9064 22100 9104
rect 17773 9055 17831 9061
rect 22094 9052 22100 9064
rect 22152 9052 22158 9104
rect 13814 9024 13820 9036
rect 12406 8996 13820 9024
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 14734 8984 14740 9036
rect 14792 8984 14798 9036
rect 14918 8984 14924 9036
rect 14976 8984 14982 9036
rect 16025 9027 16083 9033
rect 16025 8993 16037 9027
rect 16071 9024 16083 9027
rect 16850 9024 16856 9036
rect 16071 8996 16856 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 7466 8916 7472 8968
rect 7524 8916 7530 8968
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 10284 8928 10885 8956
rect 10284 8916 10290 8928
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 12066 8916 12072 8968
rect 12124 8916 12130 8968
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12492 8928 13001 8956
rect 12492 8916 12498 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8956 13783 8959
rect 14645 8959 14703 8965
rect 14645 8956 14657 8959
rect 13771 8928 14657 8956
rect 13771 8925 13783 8928
rect 13725 8919 13783 8925
rect 14645 8925 14657 8928
rect 14691 8925 14703 8959
rect 18414 8956 18420 8968
rect 17434 8928 18420 8956
rect 14645 8919 14703 8925
rect 18414 8916 18420 8928
rect 18472 8916 18478 8968
rect 8846 8888 8852 8900
rect 5368 8860 8852 8888
rect 8846 8848 8852 8860
rect 8904 8848 8910 8900
rect 10318 8888 10324 8900
rect 9784 8860 10324 8888
rect 2869 8823 2927 8829
rect 2869 8789 2881 8823
rect 2915 8820 2927 8823
rect 6454 8820 6460 8832
rect 2915 8792 6460 8820
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 6730 8780 6736 8832
rect 6788 8820 6794 8832
rect 9784 8820 9812 8860
rect 10318 8848 10324 8860
rect 10376 8848 10382 8900
rect 12084 8888 12112 8916
rect 11624 8860 12112 8888
rect 6788 8792 9812 8820
rect 6788 8780 6794 8792
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 11624 8829 11652 8860
rect 13078 8848 13084 8900
rect 13136 8888 13142 8900
rect 13136 8860 16068 8888
rect 13136 8848 13142 8860
rect 10781 8823 10839 8829
rect 10781 8820 10793 8823
rect 9916 8792 10793 8820
rect 9916 8780 9922 8792
rect 10781 8789 10793 8792
rect 10827 8789 10839 8823
rect 10781 8783 10839 8789
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8789 11667 8823
rect 11609 8783 11667 8789
rect 11974 8780 11980 8832
rect 12032 8780 12038 8832
rect 12066 8780 12072 8832
rect 12124 8780 12130 8832
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 13630 8820 13636 8832
rect 12676 8792 13636 8820
rect 12676 8780 12682 8792
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 14277 8823 14335 8829
rect 14277 8789 14289 8823
rect 14323 8820 14335 8823
rect 15930 8820 15936 8832
rect 14323 8792 15936 8820
rect 14323 8789 14335 8792
rect 14277 8783 14335 8789
rect 15930 8780 15936 8792
rect 15988 8780 15994 8832
rect 16040 8820 16068 8860
rect 16298 8848 16304 8900
rect 16356 8848 16362 8900
rect 19426 8888 19432 8900
rect 17604 8860 19432 8888
rect 17604 8820 17632 8860
rect 19426 8848 19432 8860
rect 19484 8848 19490 8900
rect 16040 8792 17632 8820
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 3602 8616 3608 8628
rect 1780 8588 3608 8616
rect 1780 8489 1808 8588
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 4430 8576 4436 8628
rect 4488 8616 4494 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 4488 8588 5825 8616
rect 4488 8576 4494 8588
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 11790 8616 11796 8628
rect 5813 8579 5871 8585
rect 6656 8588 11796 8616
rect 6656 8557 6684 8588
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12802 8616 12808 8628
rect 11931 8588 12808 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 13078 8576 13084 8628
rect 13136 8576 13142 8628
rect 14737 8619 14795 8625
rect 14737 8616 14749 8619
rect 13372 8588 14749 8616
rect 6641 8551 6699 8557
rect 6641 8517 6653 8551
rect 6687 8517 6699 8551
rect 6641 8511 6699 8517
rect 6825 8551 6883 8557
rect 6825 8517 6837 8551
rect 6871 8548 6883 8551
rect 7558 8548 7564 8560
rect 6871 8520 7564 8548
rect 6871 8517 6883 8520
rect 6825 8511 6883 8517
rect 7558 8508 7564 8520
rect 7616 8508 7622 8560
rect 11330 8548 11336 8560
rect 9416 8520 11336 8548
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8480 2467 8483
rect 2866 8480 2872 8492
rect 2455 8452 2872 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3510 8480 3516 8492
rect 3099 8452 3516 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 5994 8440 6000 8492
rect 6052 8440 6058 8492
rect 7742 8440 7748 8492
rect 7800 8440 7806 8492
rect 8938 8440 8944 8492
rect 8996 8440 9002 8492
rect 9416 8489 9444 8520
rect 11330 8508 11336 8520
rect 11388 8508 11394 8560
rect 13372 8548 13400 8588
rect 14737 8585 14749 8588
rect 14783 8585 14795 8619
rect 14737 8579 14795 8585
rect 11440 8520 13400 8548
rect 13449 8551 13507 8557
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8480 9735 8483
rect 9950 8480 9956 8492
rect 9723 8452 9956 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 11440 8480 11468 8520
rect 13449 8517 13461 8551
rect 13495 8548 13507 8551
rect 13495 8520 15700 8548
rect 13495 8517 13507 8520
rect 13449 8511 13507 8517
rect 11164 8452 11468 8480
rect 12253 8483 12311 8489
rect 2038 8412 2044 8424
rect 1596 8384 2044 8412
rect 1596 8353 1624 8384
rect 2038 8372 2044 8384
rect 2096 8372 2102 8424
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8381 7527 8415
rect 7469 8375 7527 8381
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8313 1639 8347
rect 1581 8307 1639 8313
rect 1670 8304 1676 8356
rect 1728 8344 1734 8356
rect 2225 8347 2283 8353
rect 2225 8344 2237 8347
rect 1728 8316 2237 8344
rect 1728 8304 1734 8316
rect 2225 8313 2237 8316
rect 2271 8313 2283 8347
rect 2225 8307 2283 8313
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8344 2927 8347
rect 4246 8344 4252 8356
rect 2915 8316 4252 8344
rect 2915 8313 2927 8316
rect 2869 8307 2927 8313
rect 4246 8304 4252 8316
rect 4304 8304 4310 8356
rect 7484 8344 7512 8375
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 11164 8412 11192 8452
rect 12253 8449 12265 8483
rect 12299 8480 12311 8483
rect 13354 8480 13360 8492
rect 12299 8452 13360 8480
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8480 14703 8483
rect 15378 8480 15384 8492
rect 14691 8452 15384 8480
rect 14691 8449 14703 8452
rect 14645 8443 14703 8449
rect 15378 8440 15384 8452
rect 15436 8440 15442 8492
rect 15672 8489 15700 8520
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 16942 8440 16948 8492
rect 17000 8480 17006 8492
rect 17037 8483 17095 8489
rect 17037 8480 17049 8483
rect 17000 8452 17049 8480
rect 17000 8440 17006 8452
rect 17037 8449 17049 8452
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 9272 8384 11192 8412
rect 9272 8372 9278 8384
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 12345 8415 12403 8421
rect 12345 8412 12357 8415
rect 11296 8384 12357 8412
rect 11296 8372 11302 8384
rect 12345 8381 12357 8384
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 12434 8372 12440 8424
rect 12492 8372 12498 8424
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 8757 8347 8815 8353
rect 8757 8344 8769 8347
rect 7484 8316 8769 8344
rect 8757 8313 8769 8316
rect 8803 8313 8815 8347
rect 8757 8307 8815 8313
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 13556 8344 13584 8375
rect 13722 8372 13728 8424
rect 13780 8372 13786 8424
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8412 14979 8415
rect 18322 8412 18328 8424
rect 14967 8384 18328 8412
rect 14967 8381 14979 8384
rect 14921 8375 14979 8381
rect 18322 8372 18328 8384
rect 18380 8372 18386 8424
rect 11204 8316 13584 8344
rect 11204 8304 11210 8316
rect 14274 8304 14280 8356
rect 14332 8304 14338 8356
rect 10226 8236 10232 8288
rect 10284 8276 10290 8288
rect 10873 8279 10931 8285
rect 10873 8276 10885 8279
rect 10284 8248 10885 8276
rect 10284 8236 10290 8248
rect 10873 8245 10885 8248
rect 10919 8245 10931 8279
rect 10873 8239 10931 8245
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 13998 8276 14004 8288
rect 11112 8248 14004 8276
rect 11112 8236 11118 8248
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 2130 8072 2136 8084
rect 1627 8044 2136 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 2130 8032 2136 8044
rect 2188 8032 2194 8084
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 8662 8072 8668 8084
rect 2915 8044 8668 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 9582 8032 9588 8084
rect 9640 8032 9646 8084
rect 11054 8072 11060 8084
rect 9692 8044 11060 8072
rect 7929 8007 7987 8013
rect 7929 7973 7941 8007
rect 7975 8004 7987 8007
rect 8573 8007 8631 8013
rect 8573 8004 8585 8007
rect 7975 7976 8585 8004
rect 7975 7973 7987 7976
rect 7929 7967 7987 7973
rect 8573 7973 8585 7976
rect 8619 8004 8631 8007
rect 9692 8004 9720 8044
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 12069 8075 12127 8081
rect 12069 8041 12081 8075
rect 12115 8072 12127 8075
rect 12710 8072 12716 8084
rect 12115 8044 12716 8072
rect 12115 8041 12127 8044
rect 12069 8035 12127 8041
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 13354 8032 13360 8084
rect 13412 8032 13418 8084
rect 23934 8032 23940 8084
rect 23992 8072 23998 8084
rect 28350 8072 28356 8084
rect 23992 8044 28356 8072
rect 23992 8032 23998 8044
rect 28350 8032 28356 8044
rect 28408 8032 28414 8084
rect 12434 8004 12440 8016
rect 8619 7976 9720 8004
rect 10520 7976 12440 8004
rect 8619 7973 8631 7976
rect 8573 7967 8631 7973
rect 1302 7896 1308 7948
rect 1360 7936 1366 7948
rect 1360 7908 3096 7936
rect 1360 7896 1366 7908
rect 1762 7828 1768 7880
rect 1820 7828 1826 7880
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7868 2467 7871
rect 2774 7868 2780 7880
rect 2455 7840 2780 7868
rect 2455 7837 2467 7840
rect 2409 7831 2467 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 3068 7877 3096 7908
rect 8478 7896 8484 7948
rect 8536 7936 8542 7948
rect 10520 7945 10548 7976
rect 12434 7964 12440 7976
rect 12492 7964 12498 8016
rect 12544 7976 15056 8004
rect 10505 7939 10563 7945
rect 8536 7908 10364 7936
rect 8536 7896 8542 7908
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 10226 7828 10232 7880
rect 10284 7828 10290 7880
rect 10336 7868 10364 7908
rect 10505 7905 10517 7939
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 10612 7908 10824 7936
rect 10612 7868 10640 7908
rect 10336 7840 10640 7868
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7837 10747 7871
rect 10796 7868 10824 7908
rect 10962 7896 10968 7948
rect 11020 7896 11026 7948
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 12544 7936 12572 7976
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 11572 7908 12572 7936
rect 12636 7908 14841 7936
rect 11572 7896 11578 7908
rect 12636 7868 12664 7908
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 15028 7877 15056 7976
rect 15194 7964 15200 8016
rect 15252 7964 15258 8016
rect 22186 7896 22192 7948
rect 22244 7896 22250 7948
rect 10796 7840 12664 7868
rect 15013 7871 15071 7877
rect 10689 7831 10747 7837
rect 15013 7837 15025 7871
rect 15059 7868 15071 7871
rect 15059 7840 22094 7868
rect 15059 7837 15071 7840
rect 15013 7831 15071 7837
rect 8294 7800 8300 7812
rect 2240 7772 8300 7800
rect 2240 7741 2268 7772
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 10704 7800 10732 7831
rect 16666 7800 16672 7812
rect 9876 7772 10640 7800
rect 10704 7772 16672 7800
rect 9876 7741 9904 7772
rect 2225 7735 2283 7741
rect 2225 7701 2237 7735
rect 2271 7701 2283 7735
rect 2225 7695 2283 7701
rect 9861 7735 9919 7741
rect 9861 7701 9873 7735
rect 9907 7701 9919 7735
rect 9861 7695 9919 7701
rect 10318 7692 10324 7744
rect 10376 7692 10382 7744
rect 10612 7732 10640 7772
rect 16666 7760 16672 7772
rect 16724 7760 16730 7812
rect 13446 7732 13452 7744
rect 10612 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 22066 7732 22094 7840
rect 22462 7760 22468 7812
rect 22520 7760 22526 7812
rect 23842 7800 23848 7812
rect 23690 7772 23848 7800
rect 23842 7760 23848 7772
rect 23900 7760 23906 7812
rect 22554 7732 22560 7744
rect 22066 7704 22560 7732
rect 22554 7692 22560 7704
rect 22612 7692 22618 7744
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7528 2283 7531
rect 8386 7528 8392 7540
rect 2271 7500 8392 7528
rect 2271 7497 2283 7500
rect 2225 7491 2283 7497
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 9585 7531 9643 7537
rect 9585 7497 9597 7531
rect 9631 7528 9643 7531
rect 9858 7528 9864 7540
rect 9631 7500 9864 7528
rect 9631 7497 9643 7500
rect 9585 7491 9643 7497
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 10042 7528 10048 7540
rect 9999 7500 10048 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 3694 7420 3700 7472
rect 3752 7460 3758 7472
rect 3752 7432 12112 7460
rect 3752 7420 3758 7432
rect 1394 7352 1400 7404
rect 1452 7392 1458 7404
rect 1765 7395 1823 7401
rect 1765 7392 1777 7395
rect 1452 7364 1777 7392
rect 1452 7352 1458 7364
rect 1765 7361 1777 7364
rect 1811 7361 1823 7395
rect 1765 7355 1823 7361
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 2774 7392 2780 7404
rect 2455 7364 2780 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 9364 7364 10057 7392
rect 9364 7352 9370 7364
rect 10045 7361 10057 7364
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7392 11023 7395
rect 11974 7392 11980 7404
rect 11011 7364 11980 7392
rect 11011 7361 11023 7364
rect 10965 7355 11023 7361
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12084 7401 12112 7432
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 10134 7284 10140 7336
rect 10192 7284 10198 7336
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 7650 7256 7656 7268
rect 1627 7228 7656 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 7650 7216 7656 7228
rect 7708 7216 7714 7268
rect 11885 7259 11943 7265
rect 11885 7225 11897 7259
rect 11931 7256 11943 7259
rect 15562 7256 15568 7268
rect 11931 7228 15568 7256
rect 11931 7225 11943 7228
rect 11885 7219 11943 7225
rect 15562 7216 15568 7228
rect 15620 7216 15626 7268
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7188 13691 7191
rect 16482 7188 16488 7200
rect 13679 7160 16488 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 16482 7148 16488 7160
rect 16540 7148 16546 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 23293 6987 23351 6993
rect 23293 6953 23305 6987
rect 23339 6984 23351 6987
rect 23934 6984 23940 6996
rect 23339 6956 23940 6984
rect 23339 6953 23351 6956
rect 23293 6947 23351 6953
rect 23934 6944 23940 6956
rect 23992 6944 23998 6996
rect 1762 6740 1768 6792
rect 1820 6740 1826 6792
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6749 2467 6783
rect 2409 6743 2467 6749
rect 1210 6672 1216 6724
rect 1268 6712 1274 6724
rect 2424 6712 2452 6743
rect 2866 6740 2872 6792
rect 2924 6780 2930 6792
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 2924 6752 3065 6780
rect 2924 6740 2930 6752
rect 3053 6749 3065 6752
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 20898 6740 20904 6792
rect 20956 6780 20962 6792
rect 23017 6783 23075 6789
rect 23017 6780 23029 6783
rect 20956 6752 23029 6780
rect 20956 6740 20962 6752
rect 23017 6749 23029 6752
rect 23063 6780 23075 6783
rect 27430 6780 27436 6792
rect 23063 6752 27436 6780
rect 23063 6749 23075 6752
rect 23017 6743 23075 6749
rect 27430 6740 27436 6752
rect 27488 6740 27494 6792
rect 6638 6712 6644 6724
rect 1268 6684 2452 6712
rect 2746 6684 6644 6712
rect 1268 6672 1274 6684
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 1670 6644 1676 6656
rect 1627 6616 1676 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 1670 6604 1676 6616
rect 1728 6604 1734 6656
rect 2225 6647 2283 6653
rect 2225 6613 2237 6647
rect 2271 6644 2283 6647
rect 2746 6644 2774 6684
rect 6638 6672 6644 6684
rect 6696 6672 6702 6724
rect 2271 6616 2774 6644
rect 2869 6647 2927 6653
rect 2271 6613 2283 6616
rect 2225 6607 2283 6613
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 7282 6644 7288 6656
rect 2915 6616 7288 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 22094 6604 22100 6656
rect 22152 6644 22158 6656
rect 23477 6647 23535 6653
rect 23477 6644 23489 6647
rect 22152 6616 23489 6644
rect 22152 6604 22158 6616
rect 23477 6613 23489 6616
rect 23523 6613 23535 6647
rect 23477 6607 23535 6613
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 22440 6307 22498 6313
rect 22440 6273 22452 6307
rect 22486 6304 22498 6307
rect 22554 6304 22560 6316
rect 22486 6276 22560 6304
rect 22486 6273 22498 6276
rect 22440 6267 22498 6273
rect 22554 6264 22560 6276
rect 22612 6264 22618 6316
rect 934 6196 940 6248
rect 992 6236 998 6248
rect 1581 6239 1639 6245
rect 1581 6236 1593 6239
rect 992 6208 1593 6236
rect 992 6196 998 6208
rect 1581 6205 1593 6208
rect 1627 6205 1639 6239
rect 1581 6199 1639 6205
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 11698 6236 11704 6248
rect 1903 6208 11704 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 22511 6103 22569 6109
rect 22511 6069 22523 6103
rect 22557 6100 22569 6103
rect 24762 6100 24768 6112
rect 22557 6072 24768 6100
rect 22557 6069 22569 6072
rect 22511 6063 22569 6069
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 18877 5899 18935 5905
rect 18877 5865 18889 5899
rect 18923 5896 18935 5899
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 18923 5868 21005 5896
rect 18923 5865 18935 5868
rect 18877 5859 18935 5865
rect 20993 5865 21005 5868
rect 21039 5896 21051 5899
rect 22462 5896 22468 5908
rect 21039 5868 22468 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 12618 5788 12624 5840
rect 12676 5828 12682 5840
rect 12676 5800 17264 5828
rect 12676 5788 12682 5800
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 15764 5769 15792 5800
rect 15565 5763 15623 5769
rect 15565 5760 15577 5763
rect 15528 5732 15577 5760
rect 15528 5720 15534 5732
rect 15565 5729 15577 5732
rect 15611 5729 15623 5763
rect 15565 5723 15623 5729
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5729 15807 5763
rect 15749 5723 15807 5729
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 17129 5763 17187 5769
rect 17129 5760 17141 5763
rect 16908 5732 17141 5760
rect 16908 5720 16914 5732
rect 17129 5729 17141 5732
rect 17175 5729 17187 5763
rect 17236 5760 17264 5800
rect 22094 5760 22100 5772
rect 17236 5732 22100 5760
rect 17129 5723 17187 5729
rect 22094 5720 22100 5732
rect 22152 5720 22158 5772
rect 24762 5720 24768 5772
rect 24820 5720 24826 5772
rect 26881 5763 26939 5769
rect 26881 5729 26893 5763
rect 26927 5760 26939 5763
rect 28902 5760 28908 5772
rect 26927 5732 28908 5760
rect 26927 5729 26939 5732
rect 26881 5723 26939 5729
rect 28902 5720 28908 5732
rect 28960 5720 28966 5772
rect 934 5652 940 5704
rect 992 5692 998 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 992 5664 1593 5692
rect 992 5652 998 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 10594 5692 10600 5704
rect 1903 5664 10600 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 20898 5652 20904 5704
rect 20956 5652 20962 5704
rect 24581 5695 24639 5701
rect 24581 5661 24593 5695
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 17402 5584 17408 5636
rect 17460 5584 17466 5636
rect 18414 5584 18420 5636
rect 18472 5584 18478 5636
rect 24596 5624 24624 5655
rect 25498 5624 25504 5636
rect 24596 5596 25504 5624
rect 25498 5584 25504 5596
rect 25556 5584 25562 5636
rect 26421 5627 26479 5633
rect 26421 5593 26433 5627
rect 26467 5593 26479 5627
rect 26421 5587 26479 5593
rect 16209 5559 16267 5565
rect 16209 5525 16221 5559
rect 16255 5556 16267 5559
rect 17034 5556 17040 5568
rect 16255 5528 17040 5556
rect 16255 5525 16267 5528
rect 16209 5519 16267 5525
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 21358 5516 21364 5568
rect 21416 5516 21422 5568
rect 26436 5556 26464 5587
rect 27062 5584 27068 5636
rect 27120 5584 27126 5636
rect 28718 5584 28724 5636
rect 28776 5584 28782 5636
rect 27614 5556 27620 5568
rect 26436 5528 27620 5556
rect 27614 5516 27620 5528
rect 27672 5556 27678 5568
rect 28350 5556 28356 5568
rect 27672 5528 28356 5556
rect 27672 5516 27678 5528
rect 28350 5516 28356 5528
rect 28408 5516 28414 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 22879 5355 22937 5361
rect 22879 5321 22891 5355
rect 22925 5352 22937 5355
rect 27062 5352 27068 5364
rect 22925 5324 27068 5352
rect 22925 5321 22937 5324
rect 22879 5315 22937 5321
rect 27062 5312 27068 5324
rect 27120 5312 27126 5364
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 992 5188 1593 5216
rect 992 5176 998 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 7374 5216 7380 5228
rect 1903 5188 7380 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 15562 5176 15568 5228
rect 15620 5176 15626 5228
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 17497 5219 17555 5225
rect 17497 5216 17509 5219
rect 16540 5188 17509 5216
rect 16540 5176 16546 5188
rect 17497 5185 17509 5188
rect 17543 5185 17555 5219
rect 21358 5216 21364 5228
rect 17497 5179 17555 5185
rect 17604 5188 21364 5216
rect 15470 5108 15476 5160
rect 15528 5148 15534 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15528 5120 15761 5148
rect 15528 5108 15534 5120
rect 15749 5117 15761 5120
rect 15795 5148 15807 5151
rect 17604 5148 17632 5188
rect 21358 5176 21364 5188
rect 21416 5176 21422 5228
rect 22094 5176 22100 5228
rect 22152 5225 22158 5228
rect 22152 5219 22190 5225
rect 22178 5185 22190 5219
rect 22776 5219 22834 5225
rect 22776 5216 22788 5219
rect 22152 5179 22190 5185
rect 22296 5188 22788 5216
rect 22152 5176 22158 5179
rect 15795 5120 17632 5148
rect 15795 5117 15807 5120
rect 15749 5111 15807 5117
rect 17678 5108 17684 5160
rect 17736 5108 17742 5160
rect 21376 5148 21404 5176
rect 22296 5148 22324 5188
rect 22776 5185 22788 5188
rect 22822 5185 22834 5219
rect 22776 5179 22834 5185
rect 21376 5120 22324 5148
rect 28629 5151 28687 5157
rect 28629 5117 28641 5151
rect 28675 5117 28687 5151
rect 28629 5111 28687 5117
rect 28644 5080 28672 5111
rect 28810 5108 28816 5160
rect 28868 5108 28874 5160
rect 30285 5151 30343 5157
rect 30285 5117 30297 5151
rect 30331 5148 30343 5151
rect 30374 5148 30380 5160
rect 30331 5120 30380 5148
rect 30331 5117 30343 5120
rect 30285 5111 30343 5117
rect 30374 5108 30380 5120
rect 30432 5148 30438 5160
rect 31386 5148 31392 5160
rect 30432 5120 31392 5148
rect 30432 5108 30438 5120
rect 31386 5108 31392 5120
rect 31444 5108 31450 5160
rect 33502 5080 33508 5092
rect 28644 5052 33508 5080
rect 33502 5040 33508 5052
rect 33560 5040 33566 5092
rect 16209 5015 16267 5021
rect 16209 4981 16221 5015
rect 16255 5012 16267 5015
rect 17862 5012 17868 5024
rect 16255 4984 17868 5012
rect 16255 4981 16267 4984
rect 16209 4975 16267 4981
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 18141 5015 18199 5021
rect 18141 4981 18153 5015
rect 18187 5012 18199 5015
rect 20530 5012 20536 5024
rect 18187 4984 20536 5012
rect 18187 4981 18199 4984
rect 18141 4975 18199 4981
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 22235 5015 22293 5021
rect 22235 4981 22247 5015
rect 22281 5012 22293 5015
rect 25958 5012 25964 5024
rect 22281 4984 25964 5012
rect 22281 4981 22293 4984
rect 22235 4975 22293 4981
rect 25958 4972 25964 4984
rect 26016 4972 26022 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 17402 4768 17408 4820
rect 17460 4808 17466 4820
rect 19521 4811 19579 4817
rect 19521 4808 19533 4811
rect 17460 4780 19533 4808
rect 17460 4768 17466 4780
rect 19521 4777 19533 4780
rect 19567 4777 19579 4811
rect 19521 4771 19579 4777
rect 24719 4811 24777 4817
rect 24719 4777 24731 4811
rect 24765 4808 24777 4811
rect 28810 4808 28816 4820
rect 24765 4780 28816 4808
rect 24765 4777 24777 4780
rect 24719 4771 24777 4777
rect 28810 4768 28816 4780
rect 28868 4768 28874 4820
rect 934 4632 940 4684
rect 992 4672 998 4684
rect 1581 4675 1639 4681
rect 1581 4672 1593 4675
rect 992 4644 1593 4672
rect 992 4632 998 4644
rect 1581 4641 1593 4644
rect 1627 4641 1639 4675
rect 1581 4635 1639 4641
rect 25777 4675 25835 4681
rect 25777 4641 25789 4675
rect 25823 4672 25835 4675
rect 27798 4672 27804 4684
rect 25823 4644 27804 4672
rect 25823 4641 25835 4644
rect 25777 4635 25835 4641
rect 27798 4632 27804 4644
rect 27856 4632 27862 4684
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4604 1915 4607
rect 11606 4604 11612 4616
rect 1903 4576 11612 4604
rect 1903 4573 1915 4576
rect 1857 4567 1915 4573
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 20898 4604 20904 4616
rect 19475 4576 20904 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 24616 4607 24674 4613
rect 24616 4604 24628 4607
rect 22066 4576 24628 4604
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 19889 4471 19947 4477
rect 19889 4468 19901 4471
rect 17736 4440 19901 4468
rect 17736 4428 17742 4440
rect 19889 4437 19901 4440
rect 19935 4468 19947 4471
rect 22066 4468 22094 4576
rect 24616 4573 24628 4576
rect 24662 4573 24674 4607
rect 24616 4567 24674 4573
rect 25958 4496 25964 4548
rect 26016 4496 26022 4548
rect 27338 4496 27344 4548
rect 27396 4536 27402 4548
rect 27522 4536 27528 4548
rect 27396 4508 27528 4536
rect 27396 4496 27402 4508
rect 27522 4496 27528 4508
rect 27580 4536 27586 4548
rect 27617 4539 27675 4545
rect 27617 4536 27629 4539
rect 27580 4508 27629 4536
rect 27580 4496 27586 4508
rect 27617 4505 27629 4508
rect 27663 4505 27675 4539
rect 27617 4499 27675 4505
rect 19935 4440 22094 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 1302 4088 1308 4140
rect 1360 4128 1366 4140
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 1360 4100 3065 4128
rect 1360 4088 1366 4100
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 934 4020 940 4072
rect 992 4060 998 4072
rect 1581 4063 1639 4069
rect 1581 4060 1593 4063
rect 992 4032 1593 4060
rect 992 4020 998 4032
rect 1581 4029 1593 4032
rect 1627 4029 1639 4063
rect 1581 4023 1639 4029
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4060 1915 4063
rect 9214 4060 9220 4072
rect 1903 4032 9220 4060
rect 1903 4029 1915 4032
rect 1857 4023 1915 4029
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 2869 3995 2927 4001
rect 2869 3961 2881 3995
rect 2915 3992 2927 3995
rect 10318 3992 10324 4004
rect 2915 3964 10324 3992
rect 2915 3961 2927 3964
rect 2869 3955 2927 3961
rect 10318 3952 10324 3964
rect 10376 3952 10382 4004
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 6730 3924 6736 3936
rect 2832 3896 6736 3924
rect 2832 3884 2838 3896
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 15010 3884 15016 3936
rect 15068 3884 15074 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 2225 3723 2283 3729
rect 2225 3689 2237 3723
rect 2271 3720 2283 3723
rect 2774 3720 2780 3732
rect 2271 3692 2780 3720
rect 2271 3689 2283 3692
rect 2225 3683 2283 3689
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3720 2927 3723
rect 11146 3720 11152 3732
rect 2915 3692 11152 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 30374 3680 30380 3732
rect 30432 3720 30438 3732
rect 41414 3720 41420 3732
rect 30432 3692 41420 3720
rect 30432 3680 30438 3692
rect 41414 3680 41420 3692
rect 41472 3680 41478 3732
rect 1581 3655 1639 3661
rect 1581 3621 1593 3655
rect 1627 3652 1639 3655
rect 12066 3652 12072 3664
rect 1627 3624 12072 3652
rect 1627 3621 1639 3624
rect 1581 3615 1639 3621
rect 12066 3612 12072 3624
rect 12124 3612 12130 3664
rect 28718 3612 28724 3664
rect 28776 3652 28782 3664
rect 44082 3652 44088 3664
rect 28776 3624 44088 3652
rect 28776 3612 28782 3624
rect 44082 3612 44088 3624
rect 44140 3612 44146 3664
rect 27522 3544 27528 3596
rect 27580 3584 27586 3596
rect 46750 3584 46756 3596
rect 27580 3556 46756 3584
rect 27580 3544 27586 3556
rect 46750 3544 46756 3556
rect 46808 3544 46814 3596
rect 1762 3476 1768 3528
rect 1820 3476 1826 3528
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 1210 3408 1216 3460
rect 1268 3448 1274 3460
rect 2424 3448 2452 3479
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2924 3488 3065 3516
rect 2924 3476 2930 3488
rect 3053 3485 3065 3488
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 11514 3476 11520 3528
rect 11572 3476 11578 3528
rect 28350 3476 28356 3528
rect 28408 3516 28414 3528
rect 49418 3516 49424 3528
rect 28408 3488 49424 3516
rect 28408 3476 28414 3488
rect 49418 3476 49424 3488
rect 49476 3476 49482 3528
rect 1268 3420 2452 3448
rect 1268 3408 1274 3420
rect 17126 3408 17132 3460
rect 17184 3448 17190 3460
rect 38746 3448 38752 3460
rect 17184 3420 38752 3448
rect 17184 3408 17190 3420
rect 38746 3408 38752 3420
rect 38804 3408 38810 3460
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 11238 3380 11244 3392
rect 3016 3352 11244 3380
rect 3016 3340 3022 3352
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 11606 3340 11612 3392
rect 11664 3340 11670 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 2958 3176 2964 3188
rect 2915 3148 2964 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 14001 3179 14059 3185
rect 14001 3176 14013 3179
rect 9824 3148 14013 3176
rect 9824 3136 9830 3148
rect 14001 3145 14013 3148
rect 14047 3145 14059 3179
rect 14001 3139 14059 3145
rect 7190 3108 7196 3120
rect 1872 3080 7196 3108
rect 1872 3049 1900 3080
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 9030 3068 9036 3120
rect 9088 3108 9094 3120
rect 9088 3080 9614 3108
rect 9088 3068 9094 3080
rect 12618 3068 12624 3120
rect 12676 3068 12682 3120
rect 13909 3111 13967 3117
rect 13909 3077 13921 3111
rect 13955 3108 13967 3111
rect 15470 3108 15476 3120
rect 13955 3080 15476 3108
rect 13955 3077 13967 3080
rect 13909 3071 13967 3077
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 15565 3111 15623 3117
rect 15565 3077 15577 3111
rect 15611 3108 15623 3111
rect 17678 3108 17684 3120
rect 15611 3080 17684 3108
rect 15611 3077 15623 3080
rect 15565 3071 15623 3077
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 2832 3012 3065 3040
rect 2832 3000 2838 3012
rect 3053 3009 3065 3012
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 7892 3012 8861 3040
rect 7892 3000 7898 3012
rect 8849 3009 8861 3012
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18325 3043 18383 3049
rect 18325 3040 18337 3043
rect 17920 3012 18337 3040
rect 17920 3000 17926 3012
rect 18325 3009 18337 3012
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 20530 3000 20536 3052
rect 20588 3000 20594 3052
rect 934 2932 940 2984
rect 992 2972 998 2984
rect 1581 2975 1639 2981
rect 1581 2972 1593 2975
rect 992 2944 1593 2972
rect 992 2932 998 2944
rect 1581 2941 1593 2944
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 8018 2932 8024 2984
rect 8076 2972 8082 2984
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 8076 2944 9137 2972
rect 8076 2932 8082 2944
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 10597 2975 10655 2981
rect 10597 2941 10609 2975
rect 10643 2972 10655 2975
rect 17402 2972 17408 2984
rect 10643 2944 17408 2972
rect 10643 2941 10655 2944
rect 10597 2935 10655 2941
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 12526 2864 12532 2916
rect 12584 2904 12590 2916
rect 15749 2907 15807 2913
rect 15749 2904 15761 2907
rect 12584 2876 15761 2904
rect 12584 2864 12590 2876
rect 15749 2873 15761 2876
rect 15795 2873 15807 2907
rect 15749 2867 15807 2873
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 12713 2839 12771 2845
rect 12713 2836 12725 2839
rect 8352 2808 12725 2836
rect 8352 2796 8358 2808
rect 12713 2805 12725 2808
rect 12759 2805 12771 2839
rect 12713 2799 12771 2805
rect 16853 2839 16911 2845
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 17494 2836 17500 2848
rect 16899 2808 17500 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 18141 2839 18199 2845
rect 18141 2805 18153 2839
rect 18187 2836 18199 2839
rect 20070 2836 20076 2848
rect 18187 2808 20076 2836
rect 18187 2805 18199 2808
rect 18141 2799 18199 2805
rect 20070 2796 20076 2808
rect 20128 2796 20134 2848
rect 20349 2839 20407 2845
rect 20349 2805 20361 2839
rect 20395 2836 20407 2839
rect 22002 2836 22008 2848
rect 20395 2808 22008 2836
rect 20395 2805 20407 2808
rect 20349 2799 20407 2805
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 9674 2632 9680 2644
rect 1872 2604 9680 2632
rect 1872 2505 1900 2604
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 25498 2592 25504 2644
rect 25556 2592 25562 2644
rect 27798 2592 27804 2644
rect 27856 2632 27862 2644
rect 28169 2635 28227 2641
rect 28169 2632 28181 2635
rect 27856 2604 28181 2632
rect 27856 2592 27862 2604
rect 28169 2601 28181 2604
rect 28215 2601 28227 2635
rect 28169 2595 28227 2601
rect 28902 2592 28908 2644
rect 28960 2632 28966 2644
rect 30837 2635 30895 2641
rect 30837 2632 30849 2635
rect 28960 2604 30849 2632
rect 28960 2592 28966 2604
rect 30837 2601 30849 2604
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 33502 2592 33508 2644
rect 33560 2592 33566 2644
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4120 2468 4629 2496
rect 4120 2456 4126 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6788 2468 7297 2496
rect 6788 2456 6794 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9456 2468 9965 2496
rect 9456 2456 9462 2468
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12124 2468 12633 2496
rect 12124 2456 12130 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 14734 2456 14740 2508
rect 14792 2496 14798 2508
rect 15289 2499 15347 2505
rect 15289 2496 15301 2499
rect 14792 2468 15301 2496
rect 14792 2456 14798 2468
rect 15289 2465 15301 2468
rect 15335 2465 15347 2499
rect 15289 2459 15347 2465
rect 17402 2456 17408 2508
rect 17460 2496 17466 2508
rect 17957 2499 18015 2505
rect 17957 2496 17969 2499
rect 17460 2468 17969 2496
rect 17460 2456 17466 2468
rect 17957 2465 17969 2468
rect 18003 2465 18015 2499
rect 17957 2459 18015 2465
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20220 2468 20545 2496
rect 20220 2456 20226 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22738 2456 22744 2508
rect 22796 2496 22802 2508
rect 23109 2499 23167 2505
rect 23109 2496 23121 2499
rect 22796 2468 23121 2496
rect 22796 2456 22802 2468
rect 23109 2465 23121 2468
rect 23155 2465 23167 2499
rect 23109 2459 23167 2465
rect 27430 2456 27436 2508
rect 27488 2496 27494 2508
rect 36357 2499 36415 2505
rect 36357 2496 36369 2499
rect 27488 2468 36369 2496
rect 27488 2456 27494 2468
rect 36357 2465 36369 2468
rect 36403 2465 36415 2499
rect 36357 2459 36415 2465
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 992 2400 1593 2428
rect 992 2388 998 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1762 2388 1768 2440
rect 1820 2428 1826 2440
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 1820 2400 3065 2428
rect 1820 2388 1826 2400
rect 3053 2397 3065 2400
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2397 4399 2431
rect 4341 2391 4399 2397
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 8294 2428 8300 2440
rect 7055 2400 8300 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 4356 2360 4384 2391
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 9766 2428 9772 2440
rect 9631 2400 9772 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 12526 2428 12532 2440
rect 12391 2400 12532 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12526 2388 12532 2400
rect 12584 2388 12590 2440
rect 15010 2388 15016 2440
rect 15068 2388 15074 2440
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 22002 2388 22008 2440
rect 22060 2428 22066 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22060 2400 22661 2428
rect 22060 2388 22066 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 25406 2388 25412 2440
rect 25464 2428 25470 2440
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25464 2400 25697 2428
rect 25464 2388 25470 2400
rect 25685 2397 25697 2400
rect 25731 2397 25743 2431
rect 25685 2391 25743 2397
rect 28350 2388 28356 2440
rect 28408 2388 28414 2440
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 33689 2431 33747 2437
rect 33689 2428 33701 2431
rect 33468 2400 33701 2428
rect 33468 2388 33474 2400
rect 33689 2397 33701 2400
rect 33735 2397 33747 2431
rect 33689 2391 33747 2397
rect 36078 2388 36084 2440
rect 36136 2388 36142 2440
rect 11606 2360 11612 2372
rect 4356 2332 11612 2360
rect 11606 2320 11612 2332
rect 11664 2320 11670 2372
rect 2869 2295 2927 2301
rect 2869 2261 2881 2295
rect 2915 2292 2927 2295
rect 8018 2292 8024 2304
rect 2915 2264 8024 2292
rect 2915 2261 2927 2264
rect 2869 2255 2927 2261
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
<< via1 >>
rect 20812 25508 20864 25560
rect 24124 25508 24176 25560
rect 13452 25440 13504 25492
rect 31760 25440 31812 25492
rect 10876 25372 10928 25424
rect 34520 25372 34572 25424
rect 12256 25304 12308 25356
rect 32128 25304 32180 25356
rect 11060 25236 11112 25288
rect 33416 25236 33468 25288
rect 12164 25168 12216 25220
rect 34152 25168 34204 25220
rect 9956 25100 10008 25152
rect 32036 25100 32088 25152
rect 15844 25032 15896 25084
rect 39304 25032 39356 25084
rect 11428 24964 11480 25016
rect 35900 24964 35952 25016
rect 13912 24896 13964 24948
rect 38660 24896 38712 24948
rect 3332 24828 3384 24880
rect 8576 24828 8628 24880
rect 17224 24760 17276 24812
rect 18604 24760 18656 24812
rect 22560 24828 22612 24880
rect 22284 24760 22336 24812
rect 25964 24760 26016 24812
rect 26056 24760 26108 24812
rect 28632 24760 28684 24812
rect 9588 24692 9640 24744
rect 23480 24692 23532 24744
rect 25228 24692 25280 24744
rect 29092 24692 29144 24744
rect 9128 24624 9180 24676
rect 18788 24624 18840 24676
rect 19064 24624 19116 24676
rect 25872 24624 25924 24676
rect 25964 24624 26016 24676
rect 32312 24624 32364 24676
rect 12348 24556 12400 24608
rect 25780 24556 25832 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 9128 24395 9180 24404
rect 9128 24361 9137 24395
rect 9137 24361 9171 24395
rect 9171 24361 9180 24395
rect 9128 24352 9180 24361
rect 7472 24284 7524 24336
rect 9312 24284 9364 24336
rect 3516 24216 3568 24268
rect 7380 24216 7432 24268
rect 11796 24284 11848 24336
rect 13820 24284 13872 24336
rect 2412 24148 2464 24200
rect 4804 24191 4856 24200
rect 4804 24157 4813 24191
rect 4813 24157 4847 24191
rect 4847 24157 4856 24191
rect 4804 24148 4856 24157
rect 6644 24148 6696 24200
rect 6828 24148 6880 24200
rect 9588 24148 9640 24200
rect 9956 24191 10008 24200
rect 9956 24157 9965 24191
rect 9965 24157 9999 24191
rect 9999 24157 10008 24191
rect 9956 24148 10008 24157
rect 11796 24148 11848 24200
rect 11980 24148 12032 24200
rect 12532 24191 12584 24200
rect 12532 24157 12541 24191
rect 12541 24157 12575 24191
rect 12575 24157 12584 24191
rect 12532 24148 12584 24157
rect 14280 24216 14332 24268
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 17132 24216 17184 24268
rect 10048 24080 10100 24132
rect 16212 24080 16264 24132
rect 17224 24080 17276 24132
rect 18512 24080 18564 24132
rect 4712 24012 4764 24064
rect 10140 24012 10192 24064
rect 17500 24012 17552 24064
rect 21548 24352 21600 24404
rect 18788 24148 18840 24200
rect 19800 24148 19852 24200
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 21548 24148 21600 24200
rect 21916 24148 21968 24200
rect 22560 24352 22612 24404
rect 25228 24259 25280 24268
rect 25228 24225 25237 24259
rect 25237 24225 25271 24259
rect 25271 24225 25280 24259
rect 25228 24216 25280 24225
rect 25780 24395 25832 24404
rect 25780 24361 25789 24395
rect 25789 24361 25823 24395
rect 25823 24361 25832 24395
rect 25780 24352 25832 24361
rect 25872 24352 25924 24404
rect 27252 24352 27304 24404
rect 30380 24352 30432 24404
rect 32312 24395 32364 24404
rect 32312 24361 32321 24395
rect 32321 24361 32355 24395
rect 32355 24361 32364 24395
rect 32312 24352 32364 24361
rect 33416 24395 33468 24404
rect 33416 24361 33425 24395
rect 33425 24361 33459 24395
rect 33459 24361 33468 24395
rect 33416 24352 33468 24361
rect 34152 24395 34204 24404
rect 34152 24361 34161 24395
rect 34161 24361 34195 24395
rect 34195 24361 34204 24395
rect 34152 24352 34204 24361
rect 34520 24352 34572 24404
rect 35900 24352 35952 24404
rect 39304 24395 39356 24404
rect 39304 24361 39313 24395
rect 39313 24361 39347 24395
rect 39347 24361 39356 24395
rect 39304 24352 39356 24361
rect 28080 24284 28132 24336
rect 28356 24216 28408 24268
rect 25412 24148 25464 24200
rect 26700 24148 26752 24200
rect 28632 24148 28684 24200
rect 29552 24216 29604 24268
rect 31944 24216 31996 24268
rect 30564 24148 30616 24200
rect 20812 24012 20864 24064
rect 28724 24080 28776 24132
rect 33324 24191 33376 24200
rect 33324 24157 33333 24191
rect 33333 24157 33367 24191
rect 33367 24157 33376 24191
rect 33324 24148 33376 24157
rect 33784 24148 33836 24200
rect 34520 24148 34572 24200
rect 35072 24148 35124 24200
rect 35900 24148 35952 24200
rect 37280 24148 37332 24200
rect 38476 24191 38528 24200
rect 38476 24157 38485 24191
rect 38485 24157 38519 24191
rect 38519 24157 38528 24191
rect 38476 24148 38528 24157
rect 38660 24191 38712 24200
rect 38660 24157 38669 24191
rect 38669 24157 38703 24191
rect 38703 24157 38712 24191
rect 38660 24148 38712 24157
rect 39212 24191 39264 24200
rect 39212 24157 39221 24191
rect 39221 24157 39255 24191
rect 39255 24157 39264 24191
rect 39212 24148 39264 24157
rect 40040 24259 40092 24268
rect 40040 24225 40049 24259
rect 40049 24225 40083 24259
rect 40083 24225 40092 24259
rect 40040 24216 40092 24225
rect 40592 24148 40644 24200
rect 41604 24148 41656 24200
rect 44732 24148 44784 24200
rect 45560 24148 45612 24200
rect 46020 24148 46072 24200
rect 47308 24148 47360 24200
rect 47952 24148 48004 24200
rect 34704 24080 34756 24132
rect 23940 24012 23992 24064
rect 24676 24012 24728 24064
rect 25044 24055 25096 24064
rect 25044 24021 25053 24055
rect 25053 24021 25087 24055
rect 25087 24021 25096 24055
rect 25044 24012 25096 24021
rect 25688 24012 25740 24064
rect 26240 24055 26292 24064
rect 26240 24021 26249 24055
rect 26249 24021 26283 24055
rect 26283 24021 26292 24055
rect 26240 24012 26292 24021
rect 27160 24055 27212 24064
rect 27160 24021 27169 24055
rect 27169 24021 27203 24055
rect 27203 24021 27212 24055
rect 27160 24012 27212 24021
rect 27436 24012 27488 24064
rect 27712 24012 27764 24064
rect 29000 24055 29052 24064
rect 29000 24021 29009 24055
rect 29009 24021 29043 24055
rect 29043 24021 29052 24055
rect 29000 24012 29052 24021
rect 29184 24012 29236 24064
rect 34520 24012 34572 24064
rect 40040 24080 40092 24132
rect 38660 24012 38712 24064
rect 45376 24055 45428 24064
rect 45376 24021 45385 24055
rect 45385 24021 45419 24055
rect 45419 24021 45428 24055
rect 45376 24012 45428 24021
rect 46112 24055 46164 24064
rect 46112 24021 46121 24055
rect 46121 24021 46155 24055
rect 46155 24021 46164 24055
rect 46112 24012 46164 24021
rect 46388 24012 46440 24064
rect 48780 24012 48832 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 1584 23808 1636 23860
rect 12256 23851 12308 23860
rect 12256 23817 12265 23851
rect 12265 23817 12299 23851
rect 12299 23817 12308 23851
rect 12256 23808 12308 23817
rect 12348 23851 12400 23860
rect 12348 23817 12357 23851
rect 12357 23817 12391 23851
rect 12391 23817 12400 23851
rect 12348 23808 12400 23817
rect 14464 23808 14516 23860
rect 21916 23808 21968 23860
rect 3792 23740 3844 23792
rect 4068 23740 4120 23792
rect 9680 23740 9732 23792
rect 12440 23740 12492 23792
rect 15752 23740 15804 23792
rect 19340 23740 19392 23792
rect 21456 23740 21508 23792
rect 25044 23808 25096 23860
rect 27252 23808 27304 23860
rect 27344 23808 27396 23860
rect 24492 23740 24544 23792
rect 26608 23740 26660 23792
rect 28908 23740 28960 23792
rect 29184 23740 29236 23792
rect 1124 23604 1176 23656
rect 4620 23715 4672 23724
rect 4620 23681 4629 23715
rect 4629 23681 4663 23715
rect 4663 23681 4672 23715
rect 4620 23672 4672 23681
rect 4896 23672 4948 23724
rect 7472 23715 7524 23724
rect 7472 23681 7481 23715
rect 7481 23681 7515 23715
rect 7515 23681 7524 23715
rect 7472 23672 7524 23681
rect 8116 23715 8168 23724
rect 8116 23681 8125 23715
rect 8125 23681 8159 23715
rect 8159 23681 8168 23715
rect 8116 23672 8168 23681
rect 9956 23715 10008 23724
rect 9956 23681 9965 23715
rect 9965 23681 9999 23715
rect 9999 23681 10008 23715
rect 9956 23672 10008 23681
rect 10048 23672 10100 23724
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 13452 23672 13504 23724
rect 2320 23579 2372 23588
rect 2320 23545 2329 23579
rect 2329 23545 2363 23579
rect 2363 23545 2372 23579
rect 2320 23536 2372 23545
rect 13544 23604 13596 23656
rect 15200 23672 15252 23724
rect 21732 23672 21784 23724
rect 24676 23672 24728 23724
rect 15292 23536 15344 23588
rect 18328 23604 18380 23656
rect 17776 23536 17828 23588
rect 1860 23468 1912 23520
rect 12348 23468 12400 23520
rect 19064 23647 19116 23656
rect 19064 23613 19073 23647
rect 19073 23613 19107 23647
rect 19107 23613 19116 23647
rect 19064 23604 19116 23613
rect 19616 23604 19668 23656
rect 20352 23604 20404 23656
rect 21824 23536 21876 23588
rect 24860 23647 24912 23656
rect 24860 23613 24869 23647
rect 24869 23613 24903 23647
rect 24903 23613 24912 23647
rect 24860 23604 24912 23613
rect 25872 23604 25924 23656
rect 19708 23468 19760 23520
rect 20076 23468 20128 23520
rect 23756 23511 23808 23520
rect 23756 23477 23765 23511
rect 23765 23477 23799 23511
rect 23799 23477 23808 23511
rect 23756 23468 23808 23477
rect 24860 23468 24912 23520
rect 26884 23604 26936 23656
rect 27068 23672 27120 23724
rect 29000 23672 29052 23724
rect 29736 23808 29788 23860
rect 29644 23740 29696 23792
rect 32588 23740 32640 23792
rect 30012 23715 30064 23724
rect 30012 23681 30021 23715
rect 30021 23681 30055 23715
rect 30055 23681 30064 23715
rect 30012 23672 30064 23681
rect 28632 23604 28684 23656
rect 31852 23672 31904 23724
rect 30288 23647 30340 23656
rect 30288 23613 30297 23647
rect 30297 23613 30331 23647
rect 30331 23613 30340 23647
rect 30288 23604 30340 23613
rect 31208 23604 31260 23656
rect 35164 23851 35216 23860
rect 35164 23817 35173 23851
rect 35173 23817 35207 23851
rect 35207 23817 35216 23851
rect 35164 23808 35216 23817
rect 34612 23740 34664 23792
rect 46112 23808 46164 23860
rect 34060 23672 34112 23724
rect 34428 23672 34480 23724
rect 35992 23783 36044 23792
rect 35992 23749 36001 23783
rect 36001 23749 36035 23783
rect 36035 23749 36044 23783
rect 35992 23740 36044 23749
rect 43628 23783 43680 23792
rect 43628 23749 43637 23783
rect 43637 23749 43671 23783
rect 43671 23749 43680 23783
rect 43628 23740 43680 23749
rect 35072 23715 35124 23724
rect 35072 23681 35081 23715
rect 35081 23681 35115 23715
rect 35115 23681 35124 23715
rect 35072 23672 35124 23681
rect 35808 23715 35860 23724
rect 35808 23681 35817 23715
rect 35817 23681 35851 23715
rect 35851 23681 35860 23715
rect 35808 23672 35860 23681
rect 36636 23715 36688 23724
rect 36636 23681 36645 23715
rect 36645 23681 36679 23715
rect 36679 23681 36688 23715
rect 36636 23672 36688 23681
rect 37648 23672 37700 23724
rect 41144 23672 41196 23724
rect 44180 23672 44232 23724
rect 46664 23672 46716 23724
rect 48320 23715 48372 23724
rect 48320 23681 48329 23715
rect 48329 23681 48363 23715
rect 48363 23681 48372 23715
rect 48320 23672 48372 23681
rect 49056 23715 49108 23724
rect 49056 23681 49065 23715
rect 49065 23681 49099 23715
rect 49099 23681 49108 23715
rect 49056 23672 49108 23681
rect 26240 23536 26292 23588
rect 26608 23511 26660 23520
rect 26608 23477 26617 23511
rect 26617 23477 26651 23511
rect 26651 23477 26660 23511
rect 26608 23468 26660 23477
rect 31024 23536 31076 23588
rect 37188 23604 37240 23656
rect 28724 23468 28776 23520
rect 30564 23468 30616 23520
rect 31760 23468 31812 23520
rect 35256 23468 35308 23520
rect 37740 23511 37792 23520
rect 37740 23477 37749 23511
rect 37749 23477 37783 23511
rect 37783 23477 37792 23511
rect 37740 23468 37792 23477
rect 41328 23511 41380 23520
rect 41328 23477 41337 23511
rect 41337 23477 41371 23511
rect 41371 23477 41380 23511
rect 41328 23468 41380 23477
rect 46940 23511 46992 23520
rect 46940 23477 46949 23511
rect 46949 23477 46983 23511
rect 46983 23477 46992 23511
rect 46940 23468 46992 23477
rect 48504 23511 48556 23520
rect 48504 23477 48513 23511
rect 48513 23477 48547 23511
rect 48547 23477 48556 23511
rect 48504 23468 48556 23477
rect 48688 23468 48740 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 1676 23264 1728 23316
rect 16212 23264 16264 23316
rect 18972 23264 19024 23316
rect 19524 23264 19576 23316
rect 2872 23196 2924 23248
rect 4160 23196 4212 23248
rect 9036 23196 9088 23248
rect 19064 23196 19116 23248
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 12440 23128 12492 23180
rect 12716 23128 12768 23180
rect 15200 23128 15252 23180
rect 17408 23128 17460 23180
rect 1768 23103 1820 23112
rect 1768 23069 1777 23103
rect 1777 23069 1811 23103
rect 1811 23069 1820 23103
rect 1768 23060 1820 23069
rect 2780 23035 2832 23044
rect 2780 23001 2789 23035
rect 2789 23001 2823 23035
rect 2823 23001 2832 23035
rect 2780 22992 2832 23001
rect 5448 23103 5500 23112
rect 5448 23069 5457 23103
rect 5457 23069 5491 23103
rect 5491 23069 5500 23103
rect 5448 23060 5500 23069
rect 7288 23103 7340 23112
rect 7288 23069 7297 23103
rect 7297 23069 7331 23103
rect 7331 23069 7340 23103
rect 7288 23060 7340 23069
rect 8484 23060 8536 23112
rect 10968 23060 11020 23112
rect 3884 22924 3936 22976
rect 4804 22924 4856 22976
rect 4988 22924 5040 22976
rect 8208 22924 8260 22976
rect 9496 23035 9548 23044
rect 9496 23001 9505 23035
rect 9505 23001 9539 23035
rect 9539 23001 9548 23035
rect 9496 22992 9548 23001
rect 10784 22992 10836 23044
rect 16948 23060 17000 23112
rect 17132 23103 17184 23112
rect 17132 23069 17141 23103
rect 17141 23069 17175 23103
rect 17175 23069 17184 23103
rect 17132 23060 17184 23069
rect 18512 23060 18564 23112
rect 24768 23264 24820 23316
rect 25872 23264 25924 23316
rect 27436 23264 27488 23316
rect 27620 23264 27672 23316
rect 29736 23264 29788 23316
rect 22284 23196 22336 23248
rect 23756 23196 23808 23248
rect 19708 23128 19760 23180
rect 20352 23128 20404 23180
rect 21456 23060 21508 23112
rect 10968 22967 11020 22976
rect 10968 22933 10977 22967
rect 10977 22933 11011 22967
rect 11011 22933 11020 22967
rect 10968 22924 11020 22933
rect 13820 22992 13872 23044
rect 12624 22924 12676 22976
rect 13176 22967 13228 22976
rect 13176 22933 13185 22967
rect 13185 22933 13219 22967
rect 13219 22933 13228 22967
rect 13176 22924 13228 22933
rect 15292 22992 15344 23044
rect 17500 22992 17552 23044
rect 20352 23035 20404 23044
rect 20352 23001 20361 23035
rect 20361 23001 20395 23035
rect 20395 23001 20404 23035
rect 20352 22992 20404 23001
rect 25136 23171 25188 23180
rect 25136 23137 25145 23171
rect 25145 23137 25179 23171
rect 25179 23137 25188 23171
rect 25136 23128 25188 23137
rect 25688 23128 25740 23180
rect 25872 23128 25924 23180
rect 22284 23103 22336 23112
rect 22284 23069 22293 23103
rect 22293 23069 22327 23103
rect 22327 23069 22336 23103
rect 22284 23060 22336 23069
rect 23848 23060 23900 23112
rect 25964 23060 26016 23112
rect 24492 22992 24544 23044
rect 27068 23128 27120 23180
rect 29092 23239 29144 23248
rect 29092 23205 29101 23239
rect 29101 23205 29135 23239
rect 29135 23205 29144 23239
rect 29092 23196 29144 23205
rect 29184 23196 29236 23248
rect 30012 23264 30064 23316
rect 31116 23196 31168 23248
rect 32128 23307 32180 23316
rect 32128 23273 32137 23307
rect 32137 23273 32171 23307
rect 32171 23273 32180 23307
rect 32128 23264 32180 23273
rect 28264 23128 28316 23180
rect 28356 23128 28408 23180
rect 29000 23060 29052 23112
rect 29184 23060 29236 23112
rect 40040 23196 40092 23248
rect 21824 22967 21876 22976
rect 21824 22933 21833 22967
rect 21833 22933 21867 22967
rect 21867 22933 21876 22967
rect 21824 22924 21876 22933
rect 23388 22924 23440 22976
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 24952 22967 25004 22976
rect 24952 22933 24961 22967
rect 24961 22933 24995 22967
rect 24995 22933 25004 22967
rect 24952 22924 25004 22933
rect 25780 22967 25832 22976
rect 25780 22933 25789 22967
rect 25789 22933 25823 22967
rect 25823 22933 25832 22967
rect 25780 22924 25832 22933
rect 27712 22924 27764 22976
rect 29092 22992 29144 23044
rect 28632 22924 28684 22976
rect 29552 22924 29604 22976
rect 48596 23103 48648 23112
rect 48596 23069 48605 23103
rect 48605 23069 48639 23103
rect 48639 23069 48648 23103
rect 48596 23060 48648 23069
rect 49056 23103 49108 23112
rect 49056 23069 49065 23103
rect 49065 23069 49099 23103
rect 49099 23069 49108 23103
rect 49056 23060 49108 23069
rect 32680 23035 32732 23044
rect 32680 23001 32689 23035
rect 32689 23001 32723 23035
rect 32723 23001 32732 23035
rect 32680 22992 32732 23001
rect 34152 23035 34204 23044
rect 34152 23001 34161 23035
rect 34161 23001 34195 23035
rect 34195 23001 34204 23035
rect 34152 22992 34204 23001
rect 31484 22967 31536 22976
rect 31484 22933 31493 22967
rect 31493 22933 31527 22967
rect 31527 22933 31536 22967
rect 31484 22924 31536 22933
rect 32772 22967 32824 22976
rect 32772 22933 32781 22967
rect 32781 22933 32815 22967
rect 32815 22933 32824 22967
rect 32772 22924 32824 22933
rect 33508 22967 33560 22976
rect 33508 22933 33517 22967
rect 33517 22933 33551 22967
rect 33551 22933 33560 22967
rect 33508 22924 33560 22933
rect 34244 22967 34296 22976
rect 34244 22933 34253 22967
rect 34253 22933 34287 22967
rect 34287 22933 34296 22967
rect 34244 22924 34296 22933
rect 42800 22924 42852 22976
rect 48412 22967 48464 22976
rect 48412 22933 48421 22967
rect 48421 22933 48455 22967
rect 48455 22933 48464 22967
rect 48412 22924 48464 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 1768 22652 1820 22704
rect 14464 22720 14516 22772
rect 1676 22627 1728 22636
rect 1676 22593 1685 22627
rect 1685 22593 1719 22627
rect 1719 22593 1728 22627
rect 1676 22584 1728 22593
rect 6920 22652 6972 22704
rect 10692 22695 10744 22704
rect 10692 22661 10701 22695
rect 10701 22661 10735 22695
rect 10735 22661 10744 22695
rect 10692 22652 10744 22661
rect 11888 22652 11940 22704
rect 12624 22652 12676 22704
rect 16120 22695 16172 22704
rect 16120 22661 16129 22695
rect 16129 22661 16163 22695
rect 16163 22661 16172 22695
rect 16120 22652 16172 22661
rect 2872 22516 2924 22568
rect 3700 22516 3752 22568
rect 4252 22516 4304 22568
rect 3516 22448 3568 22500
rect 7012 22584 7064 22636
rect 7840 22584 7892 22636
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 7380 22559 7432 22568
rect 7380 22525 7389 22559
rect 7389 22525 7423 22559
rect 7423 22525 7432 22559
rect 7380 22516 7432 22525
rect 5356 22448 5408 22500
rect 9956 22627 10008 22636
rect 9956 22593 9965 22627
rect 9965 22593 9999 22627
rect 9999 22593 10008 22627
rect 9956 22584 10008 22593
rect 11980 22584 12032 22636
rect 13820 22584 13872 22636
rect 16580 22584 16632 22636
rect 19708 22720 19760 22772
rect 20352 22720 20404 22772
rect 25136 22720 25188 22772
rect 26148 22720 26200 22772
rect 27620 22763 27672 22772
rect 27620 22729 27629 22763
rect 27629 22729 27663 22763
rect 27663 22729 27672 22763
rect 27620 22720 27672 22729
rect 18512 22652 18564 22704
rect 19156 22584 19208 22636
rect 20076 22652 20128 22704
rect 21456 22584 21508 22636
rect 23664 22652 23716 22704
rect 24676 22652 24728 22704
rect 24492 22584 24544 22636
rect 25228 22584 25280 22636
rect 25504 22584 25556 22636
rect 8668 22559 8720 22568
rect 8668 22525 8677 22559
rect 8677 22525 8711 22559
rect 8711 22525 8720 22559
rect 8668 22516 8720 22525
rect 12440 22559 12492 22568
rect 12440 22525 12449 22559
rect 12449 22525 12483 22559
rect 12483 22525 12492 22559
rect 12440 22516 12492 22525
rect 10508 22448 10560 22500
rect 10784 22448 10836 22500
rect 3424 22423 3476 22432
rect 3424 22389 3433 22423
rect 3433 22389 3467 22423
rect 3467 22389 3476 22423
rect 3424 22380 3476 22389
rect 3608 22380 3660 22432
rect 4528 22380 4580 22432
rect 6644 22380 6696 22432
rect 6828 22380 6880 22432
rect 12256 22380 12308 22432
rect 13176 22380 13228 22432
rect 13452 22380 13504 22432
rect 17224 22516 17276 22568
rect 18604 22559 18656 22568
rect 18604 22525 18613 22559
rect 18613 22525 18647 22559
rect 18647 22525 18656 22559
rect 18604 22516 18656 22525
rect 22284 22516 22336 22568
rect 18512 22380 18564 22432
rect 19064 22423 19116 22432
rect 19064 22389 19073 22423
rect 19073 22389 19107 22423
rect 19107 22389 19116 22423
rect 19064 22380 19116 22389
rect 19340 22380 19392 22432
rect 21824 22380 21876 22432
rect 23388 22559 23440 22568
rect 23388 22525 23397 22559
rect 23397 22525 23431 22559
rect 23431 22525 23440 22559
rect 23388 22516 23440 22525
rect 23480 22516 23532 22568
rect 24584 22516 24636 22568
rect 23388 22380 23440 22432
rect 23940 22380 23992 22432
rect 27436 22652 27488 22704
rect 31484 22720 31536 22772
rect 32496 22763 32548 22772
rect 32496 22729 32505 22763
rect 32505 22729 32539 22763
rect 32539 22729 32548 22763
rect 32496 22720 32548 22729
rect 27344 22584 27396 22636
rect 26056 22516 26108 22568
rect 26148 22516 26200 22568
rect 30012 22652 30064 22704
rect 31024 22695 31076 22704
rect 31024 22661 31033 22695
rect 31033 22661 31067 22695
rect 31067 22661 31076 22695
rect 31024 22652 31076 22661
rect 31116 22652 31168 22704
rect 28356 22627 28408 22636
rect 28356 22593 28365 22627
rect 28365 22593 28399 22627
rect 28399 22593 28408 22627
rect 28356 22584 28408 22593
rect 30932 22627 30984 22636
rect 30932 22593 30941 22627
rect 30941 22593 30975 22627
rect 30975 22593 30984 22627
rect 30932 22584 30984 22593
rect 32404 22627 32456 22636
rect 32404 22593 32413 22627
rect 32413 22593 32447 22627
rect 32447 22593 32456 22627
rect 32404 22584 32456 22593
rect 33324 22584 33376 22636
rect 33508 22584 33560 22636
rect 40040 22652 40092 22704
rect 28724 22516 28776 22568
rect 48412 22516 48464 22568
rect 27804 22448 27856 22500
rect 29920 22448 29972 22500
rect 25320 22423 25372 22432
rect 25320 22389 25329 22423
rect 25329 22389 25363 22423
rect 25363 22389 25372 22423
rect 25320 22380 25372 22389
rect 25412 22380 25464 22432
rect 26608 22380 26660 22432
rect 29000 22380 29052 22432
rect 30380 22448 30432 22500
rect 31668 22448 31720 22500
rect 31576 22380 31628 22432
rect 33232 22423 33284 22432
rect 33232 22389 33241 22423
rect 33241 22389 33275 22423
rect 33275 22389 33284 22423
rect 33232 22380 33284 22389
rect 34336 22423 34388 22432
rect 34336 22389 34345 22423
rect 34345 22389 34379 22423
rect 34379 22389 34388 22423
rect 34336 22380 34388 22389
rect 39672 22423 39724 22432
rect 39672 22389 39681 22423
rect 39681 22389 39715 22423
rect 39715 22389 39724 22423
rect 39672 22380 39724 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 3608 22176 3660 22228
rect 3792 22176 3844 22228
rect 6552 22176 6604 22228
rect 6828 22176 6880 22228
rect 7012 22176 7064 22228
rect 10324 22176 10376 22228
rect 14464 22219 14516 22228
rect 14464 22185 14473 22219
rect 14473 22185 14507 22219
rect 14507 22185 14516 22219
rect 14464 22176 14516 22185
rect 6736 22108 6788 22160
rect 1308 22040 1360 22092
rect 4436 22083 4488 22092
rect 4436 22049 4445 22083
rect 4445 22049 4479 22083
rect 4479 22049 4488 22083
rect 4436 22040 4488 22049
rect 10968 22108 11020 22160
rect 15108 22108 15160 22160
rect 10600 22083 10652 22092
rect 10600 22049 10609 22083
rect 10609 22049 10643 22083
rect 10643 22049 10652 22083
rect 10600 22040 10652 22049
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 2320 21972 2372 22024
rect 7012 22015 7064 22024
rect 7012 21981 7021 22015
rect 7021 21981 7055 22015
rect 7055 21981 7064 22015
rect 7012 21972 7064 21981
rect 11152 21972 11204 22024
rect 11244 21972 11296 22024
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 19524 22176 19576 22228
rect 19984 22176 20036 22228
rect 32772 22176 32824 22228
rect 18880 22108 18932 22160
rect 19340 22108 19392 22160
rect 22836 22151 22888 22160
rect 22836 22117 22845 22151
rect 22845 22117 22879 22151
rect 22879 22117 22888 22151
rect 22836 22108 22888 22117
rect 17132 22083 17184 22092
rect 17132 22049 17141 22083
rect 17141 22049 17175 22083
rect 17175 22049 17184 22083
rect 17132 22040 17184 22049
rect 18696 22040 18748 22092
rect 18512 21972 18564 22024
rect 20168 22040 20220 22092
rect 20260 22040 20312 22092
rect 25412 22108 25464 22160
rect 27068 22108 27120 22160
rect 25136 22083 25188 22092
rect 25136 22049 25145 22083
rect 25145 22049 25179 22083
rect 25179 22049 25188 22083
rect 25136 22040 25188 22049
rect 27252 22040 27304 22092
rect 27436 22040 27488 22092
rect 19064 21972 19116 22024
rect 19294 21972 19346 22024
rect 19616 21972 19668 22024
rect 23388 21972 23440 22024
rect 24860 21972 24912 22024
rect 25780 22015 25832 22024
rect 25780 21981 25789 22015
rect 25789 21981 25823 22015
rect 25823 21981 25832 22015
rect 25780 21972 25832 21981
rect 29184 22040 29236 22092
rect 29644 22040 29696 22092
rect 31484 22108 31536 22160
rect 31576 22108 31628 22160
rect 39672 22108 39724 22160
rect 27804 21972 27856 22024
rect 34520 22040 34572 22092
rect 32588 22015 32640 22024
rect 32588 21981 32597 22015
rect 32597 21981 32631 22015
rect 32631 21981 32640 22015
rect 32588 21972 32640 21981
rect 32864 22015 32916 22024
rect 32864 21981 32873 22015
rect 32873 21981 32907 22015
rect 32907 21981 32916 22015
rect 32864 21972 32916 21981
rect 49056 22015 49108 22024
rect 49056 21981 49065 22015
rect 49065 21981 49099 22015
rect 49099 21981 49108 22015
rect 49056 21972 49108 21981
rect 6460 21904 6512 21956
rect 11888 21904 11940 21956
rect 14372 21947 14424 21956
rect 14372 21913 14381 21947
rect 14381 21913 14415 21947
rect 14415 21913 14424 21947
rect 14372 21904 14424 21913
rect 16672 21904 16724 21956
rect 17500 21904 17552 21956
rect 18788 21904 18840 21956
rect 20536 21904 20588 21956
rect 23480 21904 23532 21956
rect 23664 21947 23716 21956
rect 23664 21913 23673 21947
rect 23673 21913 23707 21947
rect 23707 21913 23716 21947
rect 23664 21904 23716 21913
rect 24676 21904 24728 21956
rect 25688 21904 25740 21956
rect 25964 21904 26016 21956
rect 26792 21904 26844 21956
rect 6000 21836 6052 21888
rect 6276 21879 6328 21888
rect 6276 21845 6285 21879
rect 6285 21845 6319 21879
rect 6319 21845 6328 21879
rect 6276 21836 6328 21845
rect 8944 21836 8996 21888
rect 9404 21836 9456 21888
rect 14924 21836 14976 21888
rect 15016 21879 15068 21888
rect 15016 21845 15025 21879
rect 15025 21845 15059 21879
rect 15059 21845 15068 21879
rect 15016 21836 15068 21845
rect 17224 21836 17276 21888
rect 18972 21836 19024 21888
rect 19340 21836 19392 21888
rect 20076 21836 20128 21888
rect 23296 21879 23348 21888
rect 23296 21845 23305 21879
rect 23305 21845 23339 21879
rect 23339 21845 23348 21879
rect 23296 21836 23348 21845
rect 23572 21836 23624 21888
rect 29184 21904 29236 21956
rect 29000 21836 29052 21888
rect 31300 21836 31352 21888
rect 31484 21879 31536 21888
rect 31484 21845 31493 21879
rect 31493 21845 31527 21879
rect 31527 21845 31536 21879
rect 31484 21836 31536 21845
rect 49240 21879 49292 21888
rect 49240 21845 49249 21879
rect 49249 21845 49283 21879
rect 49283 21845 49292 21879
rect 49240 21836 49292 21845
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 1768 21632 1820 21684
rect 6276 21632 6328 21684
rect 2136 21564 2188 21616
rect 6092 21564 6144 21616
rect 6736 21564 6788 21616
rect 7380 21607 7432 21616
rect 7380 21573 7389 21607
rect 7389 21573 7423 21607
rect 7423 21573 7432 21607
rect 7380 21564 7432 21573
rect 9588 21564 9640 21616
rect 11888 21675 11940 21684
rect 11888 21641 11897 21675
rect 11897 21641 11931 21675
rect 11931 21641 11940 21675
rect 11888 21632 11940 21641
rect 12808 21632 12860 21684
rect 18788 21632 18840 21684
rect 2320 21496 2372 21548
rect 3608 21539 3660 21548
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 2044 21471 2096 21480
rect 2044 21437 2053 21471
rect 2053 21437 2087 21471
rect 2087 21437 2096 21471
rect 2044 21428 2096 21437
rect 4160 21471 4212 21480
rect 4160 21437 4169 21471
rect 4169 21437 4203 21471
rect 4203 21437 4212 21471
rect 4160 21428 4212 21437
rect 5540 21428 5592 21480
rect 6828 21539 6880 21548
rect 6828 21505 6837 21539
rect 6837 21505 6871 21539
rect 6871 21505 6880 21539
rect 6828 21496 6880 21505
rect 9312 21496 9364 21548
rect 12072 21496 12124 21548
rect 1952 21360 2004 21412
rect 7104 21471 7156 21480
rect 7104 21437 7113 21471
rect 7113 21437 7147 21471
rect 7147 21437 7156 21471
rect 7104 21428 7156 21437
rect 9956 21428 10008 21480
rect 10048 21428 10100 21480
rect 10784 21428 10836 21480
rect 14924 21564 14976 21616
rect 19708 21632 19760 21684
rect 20536 21632 20588 21684
rect 25136 21632 25188 21684
rect 26700 21632 26752 21684
rect 26792 21632 26844 21684
rect 27252 21632 27304 21684
rect 20260 21564 20312 21616
rect 21088 21564 21140 21616
rect 23940 21564 23992 21616
rect 25228 21564 25280 21616
rect 12532 21496 12584 21548
rect 15016 21496 15068 21548
rect 1492 21292 1544 21344
rect 3332 21292 3384 21344
rect 4436 21292 4488 21344
rect 9496 21360 9548 21412
rect 13452 21428 13504 21480
rect 13820 21428 13872 21480
rect 14280 21428 14332 21480
rect 15200 21428 15252 21480
rect 7104 21292 7156 21344
rect 8484 21292 8536 21344
rect 9312 21335 9364 21344
rect 9312 21301 9321 21335
rect 9321 21301 9355 21335
rect 9355 21301 9364 21335
rect 9312 21292 9364 21301
rect 9864 21335 9916 21344
rect 9864 21301 9873 21335
rect 9873 21301 9907 21335
rect 9907 21301 9916 21335
rect 9864 21292 9916 21301
rect 9956 21292 10008 21344
rect 10784 21292 10836 21344
rect 12808 21292 12860 21344
rect 13820 21292 13872 21344
rect 14096 21292 14148 21344
rect 14740 21292 14792 21344
rect 15476 21292 15528 21344
rect 16580 21496 16632 21548
rect 22468 21539 22520 21548
rect 22468 21505 22477 21539
rect 22477 21505 22511 21539
rect 22511 21505 22520 21539
rect 22468 21496 22520 21505
rect 17040 21428 17092 21480
rect 18696 21471 18748 21480
rect 18696 21437 18705 21471
rect 18705 21437 18739 21471
rect 18739 21437 18748 21471
rect 18696 21428 18748 21437
rect 17224 21360 17276 21412
rect 18328 21360 18380 21412
rect 19064 21428 19116 21480
rect 23204 21496 23256 21548
rect 23388 21539 23440 21548
rect 23388 21505 23397 21539
rect 23397 21505 23431 21539
rect 23431 21505 23440 21539
rect 23388 21496 23440 21505
rect 29000 21564 29052 21616
rect 29736 21564 29788 21616
rect 24676 21428 24728 21480
rect 25964 21428 26016 21480
rect 27896 21496 27948 21548
rect 20536 21360 20588 21412
rect 20904 21360 20956 21412
rect 25596 21403 25648 21412
rect 25596 21369 25605 21403
rect 25605 21369 25639 21403
rect 25639 21369 25648 21403
rect 25596 21360 25648 21369
rect 27712 21428 27764 21480
rect 27804 21471 27856 21480
rect 27804 21437 27813 21471
rect 27813 21437 27847 21471
rect 27847 21437 27856 21471
rect 27804 21428 27856 21437
rect 28356 21428 28408 21480
rect 29092 21428 29144 21480
rect 32036 21632 32088 21684
rect 34152 21632 34204 21684
rect 35256 21564 35308 21616
rect 31024 21539 31076 21548
rect 31024 21505 31033 21539
rect 31033 21505 31067 21539
rect 31067 21505 31076 21539
rect 31024 21496 31076 21505
rect 31760 21496 31812 21548
rect 32220 21496 32272 21548
rect 33416 21496 33468 21548
rect 47860 21496 47912 21548
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 17500 21292 17552 21344
rect 21456 21292 21508 21344
rect 22468 21292 22520 21344
rect 25320 21292 25372 21344
rect 27252 21335 27304 21344
rect 27252 21301 27261 21335
rect 27261 21301 27295 21335
rect 27295 21301 27304 21335
rect 27252 21292 27304 21301
rect 30196 21335 30248 21344
rect 30196 21301 30205 21335
rect 30205 21301 30239 21335
rect 30239 21301 30248 21335
rect 30196 21292 30248 21301
rect 30656 21335 30708 21344
rect 30656 21301 30665 21335
rect 30665 21301 30699 21335
rect 30699 21301 30708 21335
rect 30656 21292 30708 21301
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 6000 21088 6052 21140
rect 12256 21088 12308 21140
rect 12808 21088 12860 21140
rect 17868 21088 17920 21140
rect 19524 21088 19576 21140
rect 20444 21088 20496 21140
rect 20720 21088 20772 21140
rect 21916 21088 21968 21140
rect 4988 21020 5040 21072
rect 6828 21020 6880 21072
rect 12348 21020 12400 21072
rect 5172 20952 5224 21004
rect 4344 20884 4396 20936
rect 4804 20884 4856 20936
rect 2872 20816 2924 20868
rect 4988 20816 5040 20868
rect 4160 20791 4212 20800
rect 4160 20757 4169 20791
rect 4169 20757 4203 20791
rect 4203 20757 4212 20791
rect 4160 20748 4212 20757
rect 6276 20816 6328 20868
rect 7564 20884 7616 20936
rect 8392 20952 8444 21004
rect 12624 20995 12676 21004
rect 12624 20961 12633 20995
rect 12633 20961 12667 20995
rect 12667 20961 12676 20995
rect 12624 20952 12676 20961
rect 14832 20995 14884 21004
rect 14832 20961 14841 20995
rect 14841 20961 14875 20995
rect 14875 20961 14884 20995
rect 14832 20952 14884 20961
rect 8760 20884 8812 20936
rect 9404 20884 9456 20936
rect 12716 20884 12768 20936
rect 16672 20952 16724 21004
rect 20812 21020 20864 21072
rect 30656 21088 30708 21140
rect 31852 21088 31904 21140
rect 17040 20884 17092 20936
rect 17408 20884 17460 20936
rect 7472 20816 7524 20868
rect 11336 20859 11388 20868
rect 11336 20825 11345 20859
rect 11345 20825 11379 20859
rect 11379 20825 11388 20859
rect 11336 20816 11388 20825
rect 7196 20748 7248 20800
rect 7380 20748 7432 20800
rect 11152 20748 11204 20800
rect 15476 20816 15528 20868
rect 14004 20748 14056 20800
rect 14740 20791 14792 20800
rect 14740 20757 14749 20791
rect 14749 20757 14783 20791
rect 14783 20757 14792 20791
rect 14740 20748 14792 20757
rect 15200 20791 15252 20800
rect 15200 20757 15209 20791
rect 15209 20757 15243 20791
rect 15243 20757 15252 20791
rect 15200 20748 15252 20757
rect 16856 20816 16908 20868
rect 16396 20791 16448 20800
rect 16396 20757 16405 20791
rect 16405 20757 16439 20791
rect 16439 20757 16448 20791
rect 16396 20748 16448 20757
rect 17132 20816 17184 20868
rect 18604 20995 18656 21004
rect 18604 20961 18613 20995
rect 18613 20961 18647 20995
rect 18647 20961 18656 20995
rect 18604 20952 18656 20961
rect 19064 20952 19116 21004
rect 19708 20952 19760 21004
rect 20352 20952 20404 21004
rect 21180 20952 21232 21004
rect 23204 20952 23256 21004
rect 23664 20952 23716 21004
rect 23848 20995 23900 21004
rect 23848 20961 23857 20995
rect 23857 20961 23891 20995
rect 23891 20961 23900 20995
rect 23848 20952 23900 20961
rect 25964 21020 26016 21072
rect 27528 21020 27580 21072
rect 25780 20952 25832 21004
rect 26056 20995 26108 21004
rect 26056 20961 26065 20995
rect 26065 20961 26099 20995
rect 26099 20961 26108 20995
rect 26056 20952 26108 20961
rect 28356 20952 28408 21004
rect 21088 20884 21140 20936
rect 21548 20884 21600 20936
rect 19984 20816 20036 20868
rect 17408 20791 17460 20800
rect 17408 20757 17417 20791
rect 17417 20757 17451 20791
rect 17451 20757 17460 20791
rect 17408 20748 17460 20757
rect 18420 20748 18472 20800
rect 19248 20748 19300 20800
rect 19340 20748 19392 20800
rect 20628 20748 20680 20800
rect 20720 20748 20772 20800
rect 23480 20884 23532 20936
rect 24952 20884 25004 20936
rect 27712 20884 27764 20936
rect 28448 20884 28500 20936
rect 28540 20927 28592 20936
rect 28540 20893 28549 20927
rect 28549 20893 28583 20927
rect 28583 20893 28592 20927
rect 28540 20884 28592 20893
rect 29368 20884 29420 20936
rect 29828 20884 29880 20936
rect 31300 20927 31352 20936
rect 31300 20893 31309 20927
rect 31309 20893 31343 20927
rect 31343 20893 31352 20927
rect 31300 20884 31352 20893
rect 26240 20816 26292 20868
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 27068 20816 27120 20868
rect 27712 20748 27764 20800
rect 32312 20816 32364 20868
rect 27896 20748 27948 20800
rect 28540 20748 28592 20800
rect 31024 20748 31076 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 6092 20544 6144 20596
rect 10416 20544 10468 20596
rect 11888 20587 11940 20596
rect 11888 20553 11897 20587
rect 11897 20553 11931 20587
rect 11931 20553 11940 20587
rect 11888 20544 11940 20553
rect 17224 20544 17276 20596
rect 17316 20587 17368 20596
rect 17316 20553 17325 20587
rect 17325 20553 17359 20587
rect 17359 20553 17368 20587
rect 17316 20544 17368 20553
rect 1860 20408 1912 20460
rect 6920 20476 6972 20528
rect 10232 20476 10284 20528
rect 13360 20476 13412 20528
rect 14280 20476 14332 20528
rect 18972 20476 19024 20528
rect 6552 20451 6604 20460
rect 6552 20417 6561 20451
rect 6561 20417 6595 20451
rect 6595 20417 6604 20451
rect 6552 20408 6604 20417
rect 8392 20451 8444 20460
rect 8392 20417 8401 20451
rect 8401 20417 8435 20451
rect 8435 20417 8444 20451
rect 8392 20408 8444 20417
rect 9680 20408 9732 20460
rect 10508 20408 10560 20460
rect 11060 20408 11112 20460
rect 11612 20408 11664 20460
rect 12256 20408 12308 20460
rect 15292 20408 15344 20460
rect 16396 20408 16448 20460
rect 17408 20408 17460 20460
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 5724 20383 5776 20392
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 5816 20383 5868 20392
rect 5816 20349 5825 20383
rect 5825 20349 5859 20383
rect 5859 20349 5868 20383
rect 5816 20340 5868 20349
rect 5908 20340 5960 20392
rect 7104 20340 7156 20392
rect 7472 20340 7524 20392
rect 11704 20340 11756 20392
rect 13452 20340 13504 20392
rect 13728 20383 13780 20392
rect 13728 20349 13737 20383
rect 13737 20349 13771 20383
rect 13771 20349 13780 20383
rect 13728 20340 13780 20349
rect 14096 20340 14148 20392
rect 18420 20408 18472 20460
rect 18512 20451 18564 20460
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 19708 20451 19760 20460
rect 19708 20417 19717 20451
rect 19717 20417 19751 20451
rect 19751 20417 19760 20451
rect 19708 20408 19760 20417
rect 21088 20408 21140 20460
rect 7196 20272 7248 20324
rect 5632 20204 5684 20256
rect 12532 20315 12584 20324
rect 12532 20281 12541 20315
rect 12541 20281 12575 20315
rect 12575 20281 12584 20315
rect 12532 20272 12584 20281
rect 15292 20272 15344 20324
rect 15936 20272 15988 20324
rect 18880 20340 18932 20392
rect 19984 20383 20036 20392
rect 19984 20349 19993 20383
rect 19993 20349 20027 20383
rect 20027 20349 20036 20383
rect 19984 20340 20036 20349
rect 21456 20587 21508 20596
rect 21456 20553 21465 20587
rect 21465 20553 21499 20587
rect 21499 20553 21508 20587
rect 21456 20544 21508 20553
rect 22836 20544 22888 20596
rect 27252 20544 27304 20596
rect 28908 20544 28960 20596
rect 23388 20476 23440 20528
rect 24860 20476 24912 20528
rect 26424 20476 26476 20528
rect 34704 20544 34756 20596
rect 29644 20476 29696 20528
rect 23572 20340 23624 20392
rect 10048 20204 10100 20256
rect 10416 20204 10468 20256
rect 14648 20204 14700 20256
rect 15108 20204 15160 20256
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 15568 20204 15620 20256
rect 17316 20204 17368 20256
rect 19064 20204 19116 20256
rect 21640 20272 21692 20324
rect 20536 20204 20588 20256
rect 20720 20204 20772 20256
rect 22192 20247 22244 20256
rect 22192 20213 22201 20247
rect 22201 20213 22235 20247
rect 22235 20213 22244 20247
rect 22192 20204 22244 20213
rect 24676 20340 24728 20392
rect 25228 20340 25280 20392
rect 27068 20408 27120 20460
rect 27160 20408 27212 20460
rect 27528 20451 27580 20460
rect 27528 20417 27537 20451
rect 27537 20417 27571 20451
rect 27571 20417 27580 20451
rect 27528 20408 27580 20417
rect 28356 20451 28408 20460
rect 28356 20417 28365 20451
rect 28365 20417 28399 20451
rect 28399 20417 28408 20451
rect 28356 20408 28408 20417
rect 30104 20408 30156 20460
rect 25688 20272 25740 20324
rect 30196 20340 30248 20392
rect 25872 20204 25924 20256
rect 27160 20247 27212 20256
rect 27160 20213 27169 20247
rect 27169 20213 27203 20247
rect 27203 20213 27212 20247
rect 27160 20204 27212 20213
rect 27344 20204 27396 20256
rect 30288 20204 30340 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 2504 20000 2556 20052
rect 5908 20000 5960 20052
rect 6736 20000 6788 20052
rect 10048 20000 10100 20052
rect 11704 20043 11756 20052
rect 11704 20009 11713 20043
rect 11713 20009 11747 20043
rect 11747 20009 11756 20043
rect 11704 20000 11756 20009
rect 12532 20000 12584 20052
rect 15384 20000 15436 20052
rect 8392 19932 8444 19984
rect 9220 19932 9272 19984
rect 12440 19932 12492 19984
rect 13728 19932 13780 19984
rect 18880 20000 18932 20052
rect 23572 20000 23624 20052
rect 27160 20000 27212 20052
rect 27804 20000 27856 20052
rect 19524 19932 19576 19984
rect 21548 19932 21600 19984
rect 1400 19864 1452 19916
rect 7012 19864 7064 19916
rect 7472 19864 7524 19916
rect 1768 19839 1820 19848
rect 1768 19805 1777 19839
rect 1777 19805 1811 19839
rect 1811 19805 1820 19839
rect 1768 19796 1820 19805
rect 8484 19864 8536 19916
rect 9680 19864 9732 19916
rect 15476 19864 15528 19916
rect 17132 19864 17184 19916
rect 18236 19864 18288 19916
rect 18420 19864 18472 19916
rect 19708 19864 19760 19916
rect 20536 19907 20588 19916
rect 20536 19873 20545 19907
rect 20545 19873 20579 19907
rect 20579 19873 20588 19907
rect 20536 19864 20588 19873
rect 22560 19932 22612 19984
rect 22928 19932 22980 19984
rect 27528 19932 27580 19984
rect 31392 19932 31444 19984
rect 23848 19907 23900 19916
rect 23848 19873 23857 19907
rect 23857 19873 23891 19907
rect 23891 19873 23900 19907
rect 23848 19864 23900 19873
rect 25320 19907 25372 19916
rect 25320 19873 25329 19907
rect 25329 19873 25363 19907
rect 25363 19873 25372 19907
rect 25320 19864 25372 19873
rect 26240 19864 26292 19916
rect 6276 19728 6328 19780
rect 7472 19728 7524 19780
rect 6552 19660 6604 19712
rect 6736 19660 6788 19712
rect 9772 19796 9824 19848
rect 13268 19796 13320 19848
rect 9312 19771 9364 19780
rect 9312 19737 9321 19771
rect 9321 19737 9355 19771
rect 9355 19737 9364 19771
rect 9312 19728 9364 19737
rect 8852 19660 8904 19712
rect 9404 19703 9456 19712
rect 9404 19669 9413 19703
rect 9413 19669 9447 19703
rect 9447 19669 9456 19703
rect 9404 19660 9456 19669
rect 11796 19728 11848 19780
rect 12164 19728 12216 19780
rect 13544 19728 13596 19780
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 18788 19796 18840 19848
rect 19892 19796 19944 19848
rect 21640 19796 21692 19848
rect 23388 19796 23440 19848
rect 25780 19796 25832 19848
rect 25872 19839 25924 19848
rect 25872 19805 25881 19839
rect 25881 19805 25915 19839
rect 25915 19805 25924 19839
rect 25872 19796 25924 19805
rect 27252 19796 27304 19848
rect 27436 19796 27488 19848
rect 31576 19907 31628 19916
rect 31576 19873 31585 19907
rect 31585 19873 31619 19907
rect 31619 19873 31628 19907
rect 31576 19864 31628 19873
rect 29920 19796 29972 19848
rect 15292 19728 15344 19780
rect 11244 19660 11296 19712
rect 11520 19660 11572 19712
rect 12992 19703 13044 19712
rect 12992 19669 13001 19703
rect 13001 19669 13035 19703
rect 13035 19669 13044 19703
rect 12992 19660 13044 19669
rect 18236 19728 18288 19780
rect 20812 19728 20864 19780
rect 18420 19660 18472 19712
rect 19524 19660 19576 19712
rect 19892 19660 19944 19712
rect 21364 19660 21416 19712
rect 24032 19728 24084 19780
rect 25504 19728 25556 19780
rect 26148 19771 26200 19780
rect 26148 19737 26157 19771
rect 26157 19737 26191 19771
rect 26191 19737 26200 19771
rect 26148 19728 26200 19737
rect 23664 19703 23716 19712
rect 23664 19669 23673 19703
rect 23673 19669 23707 19703
rect 23707 19669 23716 19703
rect 23664 19660 23716 19669
rect 27620 19660 27672 19712
rect 41328 19728 41380 19780
rect 31392 19703 31444 19712
rect 31392 19669 31401 19703
rect 31401 19669 31435 19703
rect 31435 19669 31444 19703
rect 31392 19660 31444 19669
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 5632 19456 5684 19508
rect 6828 19456 6880 19508
rect 8760 19499 8812 19508
rect 8760 19465 8769 19499
rect 8769 19465 8803 19499
rect 8803 19465 8812 19499
rect 8760 19456 8812 19465
rect 9956 19456 10008 19508
rect 14556 19456 14608 19508
rect 4528 19431 4580 19440
rect 4528 19397 4537 19431
rect 4537 19397 4571 19431
rect 4571 19397 4580 19431
rect 4528 19388 4580 19397
rect 6920 19388 6972 19440
rect 8576 19388 8628 19440
rect 6736 19320 6788 19372
rect 7012 19363 7064 19372
rect 7012 19329 7028 19363
rect 7028 19329 7062 19363
rect 7062 19329 7064 19363
rect 7012 19320 7064 19329
rect 8392 19320 8444 19372
rect 8668 19320 8720 19372
rect 11980 19388 12032 19440
rect 13360 19388 13412 19440
rect 13728 19388 13780 19440
rect 20628 19456 20680 19508
rect 20812 19456 20864 19508
rect 22376 19456 22428 19508
rect 22560 19456 22612 19508
rect 23572 19456 23624 19508
rect 15384 19388 15436 19440
rect 15844 19388 15896 19440
rect 17132 19388 17184 19440
rect 15660 19363 15712 19372
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 16764 19320 16816 19372
rect 2044 19295 2096 19304
rect 2044 19261 2053 19295
rect 2053 19261 2087 19295
rect 2087 19261 2096 19295
rect 2044 19252 2096 19261
rect 3424 19252 3476 19304
rect 4252 19116 4304 19168
rect 7656 19252 7708 19304
rect 13636 19252 13688 19304
rect 13728 19252 13780 19304
rect 15844 19295 15896 19304
rect 15844 19261 15853 19295
rect 15853 19261 15887 19295
rect 15887 19261 15896 19295
rect 15844 19252 15896 19261
rect 16304 19252 16356 19304
rect 18696 19388 18748 19440
rect 18880 19320 18932 19372
rect 19340 19320 19392 19372
rect 21640 19388 21692 19440
rect 21732 19388 21784 19440
rect 22652 19388 22704 19440
rect 24032 19499 24084 19508
rect 24032 19465 24041 19499
rect 24041 19465 24075 19499
rect 24075 19465 24084 19499
rect 24032 19456 24084 19465
rect 35072 19456 35124 19508
rect 29644 19388 29696 19440
rect 18052 19252 18104 19304
rect 18604 19295 18656 19304
rect 18604 19261 18613 19295
rect 18613 19261 18647 19295
rect 18647 19261 18656 19295
rect 18604 19252 18656 19261
rect 8484 19184 8536 19236
rect 11428 19184 11480 19236
rect 12992 19184 13044 19236
rect 7288 19116 7340 19168
rect 11244 19116 11296 19168
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 15292 19116 15344 19125
rect 15936 19116 15988 19168
rect 16672 19116 16724 19168
rect 16856 19159 16908 19168
rect 16856 19125 16865 19159
rect 16865 19125 16899 19159
rect 16899 19125 16908 19159
rect 16856 19116 16908 19125
rect 18328 19184 18380 19236
rect 18972 19252 19024 19304
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 18144 19159 18196 19168
rect 18144 19125 18153 19159
rect 18153 19125 18187 19159
rect 18187 19125 18196 19159
rect 18144 19116 18196 19125
rect 19616 19184 19668 19236
rect 20352 19252 20404 19304
rect 23572 19252 23624 19304
rect 24124 19363 24176 19372
rect 24124 19329 24133 19363
rect 24133 19329 24167 19363
rect 24167 19329 24176 19363
rect 24124 19320 24176 19329
rect 25044 19363 25096 19372
rect 25044 19329 25053 19363
rect 25053 19329 25087 19363
rect 25087 19329 25096 19363
rect 25044 19320 25096 19329
rect 27620 19320 27672 19372
rect 24952 19252 25004 19304
rect 25872 19295 25924 19304
rect 25872 19261 25881 19295
rect 25881 19261 25915 19295
rect 25915 19261 25924 19295
rect 25872 19252 25924 19261
rect 26332 19252 26384 19304
rect 28356 19295 28408 19304
rect 28356 19261 28365 19295
rect 28365 19261 28399 19295
rect 28399 19261 28408 19295
rect 28356 19252 28408 19261
rect 26148 19184 26200 19236
rect 26424 19184 26476 19236
rect 19984 19116 20036 19168
rect 20168 19116 20220 19168
rect 25412 19116 25464 19168
rect 25780 19116 25832 19168
rect 28448 19116 28500 19168
rect 30932 19184 30984 19236
rect 30104 19159 30156 19168
rect 30104 19125 30113 19159
rect 30113 19125 30147 19159
rect 30147 19125 30156 19159
rect 30104 19116 30156 19125
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 11520 18912 11572 18964
rect 12072 18955 12124 18964
rect 12072 18921 12081 18955
rect 12081 18921 12115 18955
rect 12115 18921 12124 18955
rect 12072 18912 12124 18921
rect 3332 18776 3384 18828
rect 4712 18708 4764 18760
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 6276 18776 6328 18828
rect 6552 18819 6604 18828
rect 6552 18785 6561 18819
rect 6561 18785 6595 18819
rect 6595 18785 6604 18819
rect 6552 18776 6604 18785
rect 2504 18683 2556 18692
rect 2504 18649 2513 18683
rect 2513 18649 2547 18683
rect 2547 18649 2556 18683
rect 2504 18640 2556 18649
rect 5172 18640 5224 18692
rect 12532 18844 12584 18896
rect 14096 18844 14148 18896
rect 8300 18776 8352 18828
rect 8760 18776 8812 18828
rect 11244 18776 11296 18828
rect 11520 18776 11572 18828
rect 11888 18776 11940 18828
rect 12256 18776 12308 18828
rect 12440 18776 12492 18828
rect 12900 18776 12952 18828
rect 13544 18776 13596 18828
rect 10508 18708 10560 18760
rect 8576 18640 8628 18692
rect 13176 18708 13228 18760
rect 13912 18708 13964 18760
rect 11428 18640 11480 18692
rect 18144 18912 18196 18964
rect 19984 18912 20036 18964
rect 23664 18912 23716 18964
rect 26148 18912 26200 18964
rect 28816 18955 28868 18964
rect 28816 18921 28825 18955
rect 28825 18921 28859 18955
rect 28859 18921 28868 18955
rect 28816 18912 28868 18921
rect 14648 18887 14700 18896
rect 14648 18853 14657 18887
rect 14657 18853 14691 18887
rect 14691 18853 14700 18887
rect 14648 18844 14700 18853
rect 17224 18844 17276 18896
rect 16120 18776 16172 18828
rect 16672 18708 16724 18760
rect 17776 18708 17828 18760
rect 20812 18844 20864 18896
rect 18328 18776 18380 18828
rect 19708 18776 19760 18828
rect 21180 18819 21232 18828
rect 21180 18785 21189 18819
rect 21189 18785 21223 18819
rect 21223 18785 21232 18819
rect 21180 18776 21232 18785
rect 21456 18819 21508 18828
rect 21456 18785 21465 18819
rect 21465 18785 21499 18819
rect 21499 18785 21508 18819
rect 21456 18776 21508 18785
rect 22100 18776 22152 18828
rect 27068 18844 27120 18896
rect 25780 18776 25832 18828
rect 27528 18776 27580 18828
rect 18696 18708 18748 18760
rect 23572 18751 23624 18760
rect 23572 18717 23581 18751
rect 23581 18717 23615 18751
rect 23615 18717 23624 18751
rect 23572 18708 23624 18717
rect 27160 18708 27212 18760
rect 30012 18776 30064 18828
rect 29000 18751 29052 18760
rect 29000 18717 29009 18751
rect 29009 18717 29043 18751
rect 29043 18717 29052 18751
rect 29000 18708 29052 18717
rect 29092 18708 29144 18760
rect 34428 18844 34480 18896
rect 45376 18844 45428 18896
rect 3332 18572 3384 18624
rect 7288 18572 7340 18624
rect 9680 18572 9732 18624
rect 10876 18615 10928 18624
rect 10876 18581 10885 18615
rect 10885 18581 10919 18615
rect 10919 18581 10928 18615
rect 10876 18572 10928 18581
rect 11888 18572 11940 18624
rect 12072 18572 12124 18624
rect 14464 18572 14516 18624
rect 15016 18640 15068 18692
rect 15476 18640 15528 18692
rect 17684 18640 17736 18692
rect 18052 18640 18104 18692
rect 18880 18640 18932 18692
rect 19708 18683 19760 18692
rect 19708 18649 19717 18683
rect 19717 18649 19751 18683
rect 19751 18649 19760 18683
rect 19708 18640 19760 18649
rect 20628 18640 20680 18692
rect 23848 18640 23900 18692
rect 24492 18640 24544 18692
rect 25688 18683 25740 18692
rect 25688 18649 25697 18683
rect 25697 18649 25731 18683
rect 25731 18649 25740 18683
rect 25688 18640 25740 18649
rect 27252 18640 27304 18692
rect 30288 18640 30340 18692
rect 30380 18640 30432 18692
rect 48504 18640 48556 18692
rect 15568 18572 15620 18624
rect 16672 18572 16724 18624
rect 18328 18615 18380 18624
rect 18328 18581 18337 18615
rect 18337 18581 18371 18615
rect 18371 18581 18380 18615
rect 18328 18572 18380 18581
rect 21824 18572 21876 18624
rect 22928 18572 22980 18624
rect 24860 18572 24912 18624
rect 25320 18572 25372 18624
rect 26608 18572 26660 18624
rect 26700 18572 26752 18624
rect 27712 18572 27764 18624
rect 29460 18572 29512 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 5080 18368 5132 18420
rect 10968 18368 11020 18420
rect 12072 18368 12124 18420
rect 12440 18368 12492 18420
rect 2228 18300 2280 18352
rect 1952 18232 2004 18284
rect 3424 18275 3476 18284
rect 3424 18241 3433 18275
rect 3433 18241 3467 18275
rect 3467 18241 3476 18275
rect 3424 18232 3476 18241
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 9128 18300 9180 18352
rect 13728 18343 13780 18352
rect 13728 18309 13737 18343
rect 13737 18309 13771 18343
rect 13771 18309 13780 18343
rect 13728 18300 13780 18309
rect 14556 18343 14608 18352
rect 14556 18309 14565 18343
rect 14565 18309 14599 18343
rect 14599 18309 14608 18343
rect 14556 18300 14608 18309
rect 15108 18411 15160 18420
rect 15108 18377 15117 18411
rect 15117 18377 15151 18411
rect 15151 18377 15160 18411
rect 15108 18368 15160 18377
rect 20168 18368 20220 18420
rect 20352 18368 20404 18420
rect 25136 18368 25188 18420
rect 37740 18368 37792 18420
rect 17500 18300 17552 18352
rect 5632 18275 5684 18284
rect 5632 18241 5641 18275
rect 5641 18241 5675 18275
rect 5675 18241 5684 18275
rect 5632 18232 5684 18241
rect 6368 18232 6420 18284
rect 8024 18232 8076 18284
rect 4160 18164 4212 18216
rect 7012 18207 7064 18216
rect 7012 18173 7021 18207
rect 7021 18173 7055 18207
rect 7055 18173 7064 18207
rect 7012 18164 7064 18173
rect 8392 18164 8444 18216
rect 9496 18232 9548 18284
rect 11428 18232 11480 18284
rect 12808 18232 12860 18284
rect 13544 18232 13596 18284
rect 18420 18300 18472 18352
rect 18604 18300 18656 18352
rect 19248 18300 19300 18352
rect 9588 18096 9640 18148
rect 13360 18164 13412 18216
rect 16672 18164 16724 18216
rect 1584 18028 1636 18080
rect 5080 18028 5132 18080
rect 6368 18028 6420 18080
rect 7472 18028 7524 18080
rect 9496 18028 9548 18080
rect 12072 18071 12124 18080
rect 12072 18037 12081 18071
rect 12081 18037 12115 18071
rect 12115 18037 12124 18071
rect 12072 18028 12124 18037
rect 12440 18096 12492 18148
rect 12532 18096 12584 18148
rect 14464 18096 14516 18148
rect 17776 18096 17828 18148
rect 18420 18207 18472 18216
rect 18420 18173 18429 18207
rect 18429 18173 18463 18207
rect 18463 18173 18472 18207
rect 18420 18164 18472 18173
rect 19800 18232 19852 18284
rect 22468 18343 22520 18352
rect 22468 18309 22477 18343
rect 22477 18309 22511 18343
rect 22511 18309 22520 18343
rect 22468 18300 22520 18309
rect 22836 18300 22888 18352
rect 23848 18300 23900 18352
rect 25044 18300 25096 18352
rect 26056 18343 26108 18352
rect 26056 18309 26065 18343
rect 26065 18309 26099 18343
rect 26099 18309 26108 18343
rect 26056 18300 26108 18309
rect 20168 18207 20220 18216
rect 20168 18173 20177 18207
rect 20177 18173 20211 18207
rect 20211 18173 20220 18207
rect 20168 18164 20220 18173
rect 20812 18164 20864 18216
rect 21640 18164 21692 18216
rect 22928 18232 22980 18284
rect 24676 18232 24728 18284
rect 26700 18232 26752 18284
rect 27712 18232 27764 18284
rect 27804 18232 27856 18284
rect 28356 18300 28408 18352
rect 30932 18300 30984 18352
rect 29460 18232 29512 18284
rect 29644 18232 29696 18284
rect 22652 18207 22704 18216
rect 22652 18173 22661 18207
rect 22661 18173 22695 18207
rect 22695 18173 22704 18207
rect 22652 18164 22704 18173
rect 22744 18096 22796 18148
rect 12900 18028 12952 18080
rect 13176 18028 13228 18080
rect 21272 18028 21324 18080
rect 21456 18071 21508 18080
rect 21456 18037 21465 18071
rect 21465 18037 21499 18071
rect 21499 18037 21508 18071
rect 21456 18028 21508 18037
rect 22100 18071 22152 18080
rect 22100 18037 22109 18071
rect 22109 18037 22143 18071
rect 22143 18037 22152 18071
rect 22100 18028 22152 18037
rect 25320 18164 25372 18216
rect 30104 18164 30156 18216
rect 30840 18207 30892 18216
rect 30840 18173 30849 18207
rect 30849 18173 30883 18207
rect 30883 18173 30892 18207
rect 30840 18164 30892 18173
rect 24768 18028 24820 18080
rect 27528 18028 27580 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 1676 17824 1728 17876
rect 1952 17824 2004 17876
rect 4344 17867 4396 17876
rect 4344 17833 4353 17867
rect 4353 17833 4387 17867
rect 4387 17833 4396 17867
rect 4344 17824 4396 17833
rect 5172 17824 5224 17876
rect 6920 17824 6972 17876
rect 12348 17824 12400 17876
rect 13820 17824 13872 17876
rect 18328 17824 18380 17876
rect 18420 17824 18472 17876
rect 24492 17824 24544 17876
rect 26424 17824 26476 17876
rect 26608 17867 26660 17876
rect 26608 17833 26617 17867
rect 26617 17833 26651 17867
rect 26651 17833 26660 17867
rect 26608 17824 26660 17833
rect 27528 17824 27580 17876
rect 27620 17824 27672 17876
rect 1216 17688 1268 17740
rect 5816 17688 5868 17740
rect 7932 17688 7984 17740
rect 1768 17663 1820 17672
rect 1768 17629 1777 17663
rect 1777 17629 1811 17663
rect 1811 17629 1820 17663
rect 1768 17620 1820 17629
rect 4160 17620 4212 17672
rect 4804 17620 4856 17672
rect 6276 17620 6328 17672
rect 6920 17620 6972 17672
rect 9772 17756 9824 17808
rect 13636 17756 13688 17808
rect 9312 17688 9364 17740
rect 9956 17688 10008 17740
rect 13268 17688 13320 17740
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 16672 17688 16724 17740
rect 17132 17688 17184 17740
rect 18420 17688 18472 17740
rect 5080 17552 5132 17604
rect 7012 17552 7064 17604
rect 7748 17552 7800 17604
rect 8852 17552 8904 17604
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 15568 17620 15620 17672
rect 15752 17620 15804 17672
rect 17684 17620 17736 17672
rect 19248 17620 19300 17672
rect 19616 17663 19668 17672
rect 19616 17629 19625 17663
rect 19625 17629 19659 17663
rect 19659 17629 19668 17663
rect 19616 17620 19668 17629
rect 21088 17620 21140 17672
rect 10232 17552 10284 17604
rect 7932 17484 7984 17536
rect 9680 17484 9732 17536
rect 12716 17552 12768 17604
rect 15384 17552 15436 17604
rect 15936 17552 15988 17604
rect 24768 17688 24820 17740
rect 25872 17688 25924 17740
rect 27712 17688 27764 17740
rect 21916 17620 21968 17672
rect 24400 17620 24452 17672
rect 29460 17688 29512 17740
rect 30012 17688 30064 17740
rect 28816 17620 28868 17672
rect 13728 17484 13780 17536
rect 16212 17484 16264 17536
rect 18420 17484 18472 17536
rect 18880 17484 18932 17536
rect 20168 17527 20220 17536
rect 20168 17493 20177 17527
rect 20177 17493 20211 17527
rect 20211 17493 20220 17527
rect 20168 17484 20220 17493
rect 20996 17484 21048 17536
rect 21180 17527 21232 17536
rect 21180 17493 21189 17527
rect 21189 17493 21223 17527
rect 21223 17493 21232 17527
rect 21180 17484 21232 17493
rect 22468 17484 22520 17536
rect 23848 17484 23900 17536
rect 25228 17552 25280 17604
rect 26424 17552 26476 17604
rect 26700 17552 26752 17604
rect 24216 17484 24268 17536
rect 27160 17484 27212 17536
rect 30840 17552 30892 17604
rect 42800 17552 42852 17604
rect 30196 17527 30248 17536
rect 30196 17493 30205 17527
rect 30205 17493 30239 17527
rect 30239 17493 30248 17527
rect 30196 17484 30248 17493
rect 46388 17484 46440 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 7104 17280 7156 17332
rect 7196 17323 7248 17332
rect 7196 17289 7205 17323
rect 7205 17289 7239 17323
rect 7239 17289 7248 17323
rect 7196 17280 7248 17289
rect 7288 17323 7340 17332
rect 7288 17289 7297 17323
rect 7297 17289 7331 17323
rect 7331 17289 7340 17323
rect 7288 17280 7340 17289
rect 7840 17280 7892 17332
rect 9496 17280 9548 17332
rect 2320 17212 2372 17264
rect 5172 17212 5224 17264
rect 6000 17212 6052 17264
rect 8484 17255 8536 17264
rect 8484 17221 8493 17255
rect 8493 17221 8527 17255
rect 8527 17221 8536 17255
rect 8484 17212 8536 17221
rect 10048 17212 10100 17264
rect 11336 17280 11388 17332
rect 11888 17280 11940 17332
rect 20168 17280 20220 17332
rect 3332 17144 3384 17196
rect 3424 17187 3476 17196
rect 3424 17153 3433 17187
rect 3433 17153 3467 17187
rect 3467 17153 3476 17187
rect 3424 17144 3476 17153
rect 8300 17144 8352 17196
rect 1308 17076 1360 17128
rect 3792 17076 3844 17128
rect 5356 17076 5408 17128
rect 5908 17119 5960 17128
rect 5908 17085 5917 17119
rect 5917 17085 5951 17119
rect 5951 17085 5960 17119
rect 5908 17076 5960 17085
rect 7196 17076 7248 17128
rect 7656 17076 7708 17128
rect 9404 17144 9456 17196
rect 9956 17144 10008 17196
rect 10324 17144 10376 17196
rect 13912 17212 13964 17264
rect 17684 17212 17736 17264
rect 21456 17280 21508 17332
rect 21548 17280 21600 17332
rect 8576 17119 8628 17128
rect 8576 17085 8585 17119
rect 8585 17085 8619 17119
rect 8619 17085 8628 17119
rect 8576 17076 8628 17085
rect 8760 17076 8812 17128
rect 9496 17076 9548 17128
rect 9588 17076 9640 17128
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 10968 17119 11020 17128
rect 10968 17085 10977 17119
rect 10977 17085 11011 17119
rect 11011 17085 11020 17119
rect 10968 17076 11020 17085
rect 16856 17144 16908 17196
rect 6460 17008 6512 17060
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 5632 16940 5684 16992
rect 6000 16940 6052 16992
rect 8576 16940 8628 16992
rect 9312 16940 9364 16992
rect 10692 16940 10744 16992
rect 13636 17076 13688 17128
rect 12624 17008 12676 17060
rect 16028 17076 16080 17128
rect 17500 17119 17552 17128
rect 17500 17085 17509 17119
rect 17509 17085 17543 17119
rect 17543 17085 17552 17119
rect 17500 17076 17552 17085
rect 14924 17008 14976 17060
rect 16948 17008 17000 17060
rect 17040 17008 17092 17060
rect 18420 17119 18472 17128
rect 18420 17085 18429 17119
rect 18429 17085 18463 17119
rect 18463 17085 18472 17119
rect 18420 17076 18472 17085
rect 18880 17076 18932 17128
rect 22744 17280 22796 17332
rect 25136 17212 25188 17264
rect 26424 17212 26476 17264
rect 27160 17212 27212 17264
rect 14188 16940 14240 16992
rect 14832 16940 14884 16992
rect 15936 16940 15988 16992
rect 17132 16940 17184 16992
rect 19524 16940 19576 16992
rect 20260 17076 20312 17128
rect 21272 17119 21324 17128
rect 21272 17085 21281 17119
rect 21281 17085 21315 17119
rect 21315 17085 21324 17119
rect 22284 17187 22336 17196
rect 22284 17153 22293 17187
rect 22293 17153 22327 17187
rect 22327 17153 22336 17187
rect 22284 17144 22336 17153
rect 22836 17144 22888 17196
rect 23572 17144 23624 17196
rect 24492 17187 24544 17196
rect 24492 17153 24501 17187
rect 24501 17153 24535 17187
rect 24535 17153 24544 17187
rect 24492 17144 24544 17153
rect 24768 17187 24820 17196
rect 24768 17153 24777 17187
rect 24777 17153 24811 17187
rect 24811 17153 24820 17187
rect 24768 17144 24820 17153
rect 21272 17076 21324 17085
rect 22744 17008 22796 17060
rect 22836 17008 22888 17060
rect 23848 17119 23900 17128
rect 23848 17085 23857 17119
rect 23857 17085 23891 17119
rect 23891 17085 23900 17119
rect 23848 17076 23900 17085
rect 26700 17076 26752 17128
rect 30196 17280 30248 17332
rect 29460 17212 29512 17264
rect 30104 17212 30156 17264
rect 27804 17144 27856 17196
rect 30012 17076 30064 17128
rect 28172 16940 28224 16992
rect 28264 16940 28316 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 2228 16600 2280 16652
rect 8116 16736 8168 16788
rect 10232 16668 10284 16720
rect 10324 16668 10376 16720
rect 10876 16668 10928 16720
rect 5264 16600 5316 16652
rect 7196 16643 7248 16652
rect 7196 16609 7205 16643
rect 7205 16609 7239 16643
rect 7239 16609 7248 16643
rect 7196 16600 7248 16609
rect 1308 16464 1360 16516
rect 3976 16464 4028 16516
rect 5172 16464 5224 16516
rect 6552 16532 6604 16584
rect 10968 16600 11020 16652
rect 11520 16600 11572 16652
rect 12348 16736 12400 16788
rect 15936 16736 15988 16788
rect 16856 16779 16908 16788
rect 16856 16745 16865 16779
rect 16865 16745 16899 16779
rect 16899 16745 16908 16779
rect 16856 16736 16908 16745
rect 16948 16736 17000 16788
rect 12440 16643 12492 16652
rect 12440 16609 12449 16643
rect 12449 16609 12483 16643
rect 12483 16609 12492 16643
rect 12440 16600 12492 16609
rect 8208 16575 8260 16584
rect 8208 16541 8217 16575
rect 8217 16541 8251 16575
rect 8251 16541 8260 16575
rect 8208 16532 8260 16541
rect 9772 16532 9824 16584
rect 10140 16532 10192 16584
rect 10600 16575 10652 16584
rect 10600 16541 10609 16575
rect 10609 16541 10643 16575
rect 10643 16541 10652 16575
rect 10600 16532 10652 16541
rect 12072 16532 12124 16584
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 18420 16668 18472 16720
rect 18788 16779 18840 16788
rect 18788 16745 18797 16779
rect 18797 16745 18831 16779
rect 18831 16745 18840 16779
rect 18788 16736 18840 16745
rect 18880 16736 18932 16788
rect 19432 16736 19484 16788
rect 20260 16736 20312 16788
rect 21180 16736 21232 16788
rect 25780 16736 25832 16788
rect 20812 16668 20864 16720
rect 21548 16668 21600 16720
rect 22928 16668 22980 16720
rect 23388 16668 23440 16720
rect 25228 16668 25280 16720
rect 15384 16600 15436 16652
rect 15844 16600 15896 16652
rect 21272 16600 21324 16652
rect 22744 16600 22796 16652
rect 25136 16643 25188 16652
rect 25136 16609 25145 16643
rect 25145 16609 25179 16643
rect 25179 16609 25188 16643
rect 25136 16600 25188 16609
rect 25688 16600 25740 16652
rect 27068 16643 27120 16652
rect 27068 16609 27077 16643
rect 27077 16609 27111 16643
rect 27111 16609 27120 16643
rect 27068 16600 27120 16609
rect 27252 16643 27304 16652
rect 27252 16609 27261 16643
rect 27261 16609 27295 16643
rect 27295 16609 27304 16643
rect 27252 16600 27304 16609
rect 28264 16600 28316 16652
rect 31576 16600 31628 16652
rect 16764 16532 16816 16584
rect 17868 16532 17920 16584
rect 18420 16532 18472 16584
rect 19432 16575 19484 16584
rect 19432 16541 19441 16575
rect 19441 16541 19475 16575
rect 19475 16541 19484 16575
rect 19432 16532 19484 16541
rect 23480 16532 23532 16584
rect 24124 16532 24176 16584
rect 6000 16464 6052 16516
rect 6460 16396 6512 16448
rect 7380 16464 7432 16516
rect 8116 16464 8168 16516
rect 8484 16464 8536 16516
rect 10232 16464 10284 16516
rect 11152 16464 11204 16516
rect 7012 16439 7064 16448
rect 7012 16405 7021 16439
rect 7021 16405 7055 16439
rect 7055 16405 7064 16439
rect 7012 16396 7064 16405
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 9404 16396 9456 16448
rect 10140 16396 10192 16448
rect 10508 16439 10560 16448
rect 10508 16405 10517 16439
rect 10517 16405 10551 16439
rect 10551 16405 10560 16439
rect 10508 16396 10560 16405
rect 13544 16464 13596 16516
rect 11888 16396 11940 16448
rect 13268 16396 13320 16448
rect 19340 16464 19392 16516
rect 20996 16464 21048 16516
rect 21456 16507 21508 16516
rect 21456 16473 21465 16507
rect 21465 16473 21499 16507
rect 21499 16473 21508 16507
rect 21456 16464 21508 16473
rect 15384 16439 15436 16448
rect 15384 16405 15393 16439
rect 15393 16405 15427 16439
rect 15427 16405 15436 16439
rect 15384 16396 15436 16405
rect 15476 16439 15528 16448
rect 15476 16405 15485 16439
rect 15485 16405 15519 16439
rect 15519 16405 15528 16439
rect 15476 16396 15528 16405
rect 15660 16396 15712 16448
rect 19156 16396 19208 16448
rect 20720 16396 20772 16448
rect 23388 16464 23440 16516
rect 23756 16396 23808 16448
rect 24216 16396 24268 16448
rect 25228 16464 25280 16516
rect 27620 16532 27672 16584
rect 28172 16575 28224 16584
rect 28172 16541 28181 16575
rect 28181 16541 28215 16575
rect 28215 16541 28224 16575
rect 28172 16532 28224 16541
rect 25504 16464 25556 16516
rect 27896 16464 27948 16516
rect 28448 16464 28500 16516
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 6092 16192 6144 16244
rect 7564 16192 7616 16244
rect 7748 16192 7800 16244
rect 7932 16192 7984 16244
rect 12716 16192 12768 16244
rect 13360 16192 13412 16244
rect 14832 16235 14884 16244
rect 14832 16201 14841 16235
rect 14841 16201 14875 16235
rect 14875 16201 14884 16235
rect 14832 16192 14884 16201
rect 15384 16192 15436 16244
rect 20812 16192 20864 16244
rect 21088 16235 21140 16244
rect 21088 16201 21097 16235
rect 21097 16201 21131 16235
rect 21131 16201 21140 16235
rect 21088 16192 21140 16201
rect 22192 16235 22244 16244
rect 22192 16201 22201 16235
rect 22201 16201 22235 16235
rect 22235 16201 22244 16235
rect 22192 16192 22244 16201
rect 22652 16192 22704 16244
rect 22928 16192 22980 16244
rect 23756 16235 23808 16244
rect 23756 16201 23765 16235
rect 23765 16201 23799 16235
rect 23799 16201 23808 16235
rect 23756 16192 23808 16201
rect 24952 16192 25004 16244
rect 4344 16167 4396 16176
rect 4344 16133 4353 16167
rect 4353 16133 4387 16167
rect 4387 16133 4396 16167
rect 4344 16124 4396 16133
rect 1308 15988 1360 16040
rect 5724 16099 5776 16108
rect 5724 16065 5733 16099
rect 5733 16065 5767 16099
rect 5767 16065 5776 16099
rect 5724 16056 5776 16065
rect 6460 16056 6512 16108
rect 4804 15988 4856 16040
rect 6552 15988 6604 16040
rect 6552 15852 6604 15904
rect 8668 16124 8720 16176
rect 8852 16124 8904 16176
rect 10048 16124 10100 16176
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 7748 16031 7800 16040
rect 7748 15997 7757 16031
rect 7757 15997 7791 16031
rect 7791 15997 7800 16031
rect 7748 15988 7800 15997
rect 7932 16056 7984 16108
rect 8392 16056 8444 16108
rect 8024 15988 8076 16040
rect 12624 16124 12676 16176
rect 11152 16099 11204 16108
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 11152 16056 11204 16065
rect 11980 16056 12032 16108
rect 10232 16031 10284 16040
rect 10232 15997 10241 16031
rect 10241 15997 10275 16031
rect 10275 15997 10284 16031
rect 10232 15988 10284 15997
rect 10416 15988 10468 16040
rect 13544 15988 13596 16040
rect 7932 15920 7984 15972
rect 10508 15920 10560 15972
rect 10600 15852 10652 15904
rect 11520 15852 11572 15904
rect 12164 15852 12216 15904
rect 21456 16124 21508 16176
rect 27160 16124 27212 16176
rect 14464 15988 14516 16040
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 18512 16056 18564 16108
rect 18972 16056 19024 16108
rect 20168 16099 20220 16108
rect 20168 16065 20177 16099
rect 20177 16065 20211 16099
rect 20211 16065 20220 16099
rect 20168 16056 20220 16065
rect 17408 15988 17460 16040
rect 18328 15988 18380 16040
rect 23848 16031 23900 16040
rect 23848 15997 23857 16031
rect 23857 15997 23891 16031
rect 23891 15997 23900 16031
rect 23848 15988 23900 15997
rect 24860 16099 24912 16108
rect 24860 16065 24869 16099
rect 24869 16065 24903 16099
rect 24903 16065 24912 16099
rect 24860 16056 24912 16065
rect 27252 15988 27304 16040
rect 13912 15852 13964 15904
rect 16120 15895 16172 15904
rect 16120 15861 16129 15895
rect 16129 15861 16163 15895
rect 16163 15861 16172 15895
rect 16120 15852 16172 15861
rect 16672 15852 16724 15904
rect 17868 15920 17920 15972
rect 20628 15852 20680 15904
rect 21364 15852 21416 15904
rect 22560 15920 22612 15972
rect 24676 15852 24728 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 7012 15648 7064 15700
rect 7932 15648 7984 15700
rect 9496 15648 9548 15700
rect 10692 15648 10744 15700
rect 10784 15648 10836 15700
rect 8668 15580 8720 15632
rect 10232 15623 10284 15632
rect 10232 15589 10241 15623
rect 10241 15589 10275 15623
rect 10275 15589 10284 15623
rect 10232 15580 10284 15589
rect 10876 15623 10928 15632
rect 10876 15589 10885 15623
rect 10885 15589 10919 15623
rect 10919 15589 10928 15623
rect 10876 15580 10928 15589
rect 12072 15691 12124 15700
rect 12072 15657 12081 15691
rect 12081 15657 12115 15691
rect 12115 15657 12124 15691
rect 12072 15648 12124 15657
rect 12256 15648 12308 15700
rect 16120 15648 16172 15700
rect 19524 15648 19576 15700
rect 19984 15648 20036 15700
rect 15476 15580 15528 15632
rect 16028 15580 16080 15632
rect 22192 15580 22244 15632
rect 1308 15512 1360 15564
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 4712 15512 4764 15564
rect 5540 15512 5592 15564
rect 6736 15512 6788 15564
rect 7012 15555 7064 15564
rect 7012 15521 7021 15555
rect 7021 15521 7055 15555
rect 7055 15521 7064 15555
rect 7012 15512 7064 15521
rect 7380 15512 7432 15564
rect 8024 15512 8076 15564
rect 8852 15512 8904 15564
rect 2504 15444 2556 15496
rect 6368 15444 6420 15496
rect 5816 15376 5868 15428
rect 6092 15376 6144 15428
rect 4068 15308 4120 15360
rect 5172 15351 5224 15360
rect 5172 15317 5181 15351
rect 5181 15317 5215 15351
rect 5215 15317 5224 15351
rect 5172 15308 5224 15317
rect 6644 15376 6696 15428
rect 7196 15444 7248 15496
rect 9036 15444 9088 15496
rect 11428 15555 11480 15564
rect 11428 15521 11437 15555
rect 11437 15521 11471 15555
rect 11471 15521 11480 15555
rect 11428 15512 11480 15521
rect 12716 15555 12768 15564
rect 12716 15521 12725 15555
rect 12725 15521 12759 15555
rect 12759 15521 12768 15555
rect 12716 15512 12768 15521
rect 14924 15512 14976 15564
rect 16488 15512 16540 15564
rect 18420 15512 18472 15564
rect 19432 15512 19484 15564
rect 20628 15512 20680 15564
rect 22100 15512 22152 15564
rect 23756 15512 23808 15564
rect 25688 15512 25740 15564
rect 6368 15351 6420 15360
rect 6368 15317 6377 15351
rect 6377 15317 6411 15351
rect 6411 15317 6420 15351
rect 6368 15308 6420 15317
rect 8576 15376 8628 15428
rect 9220 15419 9272 15428
rect 9220 15385 9229 15419
rect 9229 15385 9263 15419
rect 9263 15385 9272 15419
rect 9220 15376 9272 15385
rect 10232 15444 10284 15496
rect 10968 15444 11020 15496
rect 11152 15444 11204 15496
rect 12072 15444 12124 15496
rect 16948 15444 17000 15496
rect 17040 15444 17092 15496
rect 19340 15444 19392 15496
rect 20996 15444 21048 15496
rect 22008 15444 22060 15496
rect 22836 15444 22888 15496
rect 10784 15376 10836 15428
rect 11336 15419 11388 15428
rect 11336 15385 11345 15419
rect 11345 15385 11379 15419
rect 11379 15385 11388 15419
rect 11336 15376 11388 15385
rect 15200 15419 15252 15428
rect 15200 15385 15209 15419
rect 15209 15385 15243 15419
rect 15243 15385 15252 15419
rect 15200 15376 15252 15385
rect 17684 15376 17736 15428
rect 19984 15419 20036 15428
rect 19984 15385 19993 15419
rect 19993 15385 20027 15419
rect 20027 15385 20036 15419
rect 19984 15376 20036 15385
rect 24584 15444 24636 15496
rect 25044 15444 25096 15496
rect 25412 15444 25464 15496
rect 26148 15444 26200 15496
rect 8208 15351 8260 15360
rect 8208 15317 8217 15351
rect 8217 15317 8251 15351
rect 8251 15317 8260 15351
rect 8208 15308 8260 15317
rect 12256 15308 12308 15360
rect 12440 15351 12492 15360
rect 12440 15317 12449 15351
rect 12449 15317 12483 15351
rect 12483 15317 12492 15351
rect 12440 15308 12492 15317
rect 14740 15308 14792 15360
rect 16304 15351 16356 15360
rect 16304 15317 16313 15351
rect 16313 15317 16347 15351
rect 16347 15317 16356 15351
rect 16304 15308 16356 15317
rect 17224 15308 17276 15360
rect 17500 15308 17552 15360
rect 19708 15308 19760 15360
rect 23940 15419 23992 15428
rect 23940 15385 23949 15419
rect 23949 15385 23983 15419
rect 23983 15385 23992 15419
rect 23940 15376 23992 15385
rect 24860 15376 24912 15428
rect 25780 15376 25832 15428
rect 21456 15351 21508 15360
rect 21456 15317 21465 15351
rect 21465 15317 21499 15351
rect 21499 15317 21508 15351
rect 21456 15308 21508 15317
rect 21548 15308 21600 15360
rect 22100 15308 22152 15360
rect 23572 15308 23624 15360
rect 24124 15308 24176 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 4804 15104 4856 15156
rect 4712 15036 4764 15088
rect 6000 15036 6052 15088
rect 8576 15104 8628 15156
rect 8852 15104 8904 15156
rect 9404 15104 9456 15156
rect 11888 15104 11940 15156
rect 12808 15104 12860 15156
rect 13820 15104 13872 15156
rect 7840 15036 7892 15088
rect 1860 14968 1912 15020
rect 4160 15011 4212 15020
rect 4160 14977 4169 15011
rect 4169 14977 4203 15011
rect 4203 14977 4212 15011
rect 4160 14968 4212 14977
rect 6276 14968 6328 15020
rect 6644 15011 6696 15020
rect 6644 14977 6653 15011
rect 6653 14977 6687 15011
rect 6687 14977 6696 15011
rect 6644 14968 6696 14977
rect 6736 14968 6788 15020
rect 1308 14900 1360 14952
rect 2320 14900 2372 14952
rect 3608 14900 3660 14952
rect 1492 14832 1544 14884
rect 7748 14900 7800 14952
rect 7932 14943 7984 14952
rect 7932 14909 7941 14943
rect 7941 14909 7975 14943
rect 7975 14909 7984 14943
rect 7932 14900 7984 14909
rect 5816 14832 5868 14884
rect 7104 14832 7156 14884
rect 7564 14832 7616 14884
rect 9312 15036 9364 15088
rect 10784 15079 10836 15088
rect 10784 15045 10793 15079
rect 10793 15045 10827 15079
rect 10827 15045 10836 15079
rect 10784 15036 10836 15045
rect 11520 15036 11572 15088
rect 15108 15036 15160 15088
rect 16948 15104 17000 15156
rect 20628 15104 20680 15156
rect 21916 15104 21968 15156
rect 21548 15036 21600 15088
rect 11428 14968 11480 15020
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14968 12032 14977
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 9496 14900 9548 14952
rect 9772 14943 9824 14952
rect 9772 14909 9781 14943
rect 9781 14909 9815 14943
rect 9815 14909 9824 14943
rect 9772 14900 9824 14909
rect 10416 14875 10468 14884
rect 10416 14841 10425 14875
rect 10425 14841 10459 14875
rect 10459 14841 10468 14875
rect 10416 14832 10468 14841
rect 7288 14764 7340 14816
rect 7932 14764 7984 14816
rect 12348 14900 12400 14952
rect 13452 14943 13504 14952
rect 13452 14909 13461 14943
rect 13461 14909 13495 14943
rect 13495 14909 13504 14943
rect 13452 14900 13504 14909
rect 13544 14943 13596 14952
rect 13544 14909 13553 14943
rect 13553 14909 13587 14943
rect 13587 14909 13596 14943
rect 13544 14900 13596 14909
rect 14556 14943 14608 14952
rect 14556 14909 14565 14943
rect 14565 14909 14599 14943
rect 14599 14909 14608 14943
rect 14556 14900 14608 14909
rect 14924 14900 14976 14952
rect 15292 14900 15344 14952
rect 15476 14900 15528 14952
rect 15844 14900 15896 14952
rect 18880 14943 18932 14952
rect 18880 14909 18889 14943
rect 18889 14909 18923 14943
rect 18923 14909 18932 14943
rect 18880 14900 18932 14909
rect 19064 14900 19116 14952
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 22284 15104 22336 15156
rect 23940 15104 23992 15156
rect 24952 15104 25004 15156
rect 23572 15036 23624 15088
rect 24400 15036 24452 15088
rect 27160 15036 27212 15088
rect 23940 14968 23992 15020
rect 23756 14943 23808 14952
rect 23756 14909 23765 14943
rect 23765 14909 23799 14943
rect 23799 14909 23808 14943
rect 23756 14900 23808 14909
rect 21456 14832 21508 14884
rect 11612 14764 11664 14816
rect 16120 14764 16172 14816
rect 22468 14764 22520 14816
rect 26608 14807 26660 14816
rect 26608 14773 26617 14807
rect 26617 14773 26651 14807
rect 26651 14773 26660 14807
rect 26608 14764 26660 14773
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 4068 14560 4120 14612
rect 12256 14560 12308 14612
rect 14740 14560 14792 14612
rect 15292 14560 15344 14612
rect 6644 14492 6696 14544
rect 1308 14424 1360 14476
rect 5540 14467 5592 14476
rect 5540 14433 5549 14467
rect 5549 14433 5583 14467
rect 5583 14433 5592 14467
rect 5540 14424 5592 14433
rect 5632 14424 5684 14476
rect 6000 14424 6052 14476
rect 6552 14424 6604 14476
rect 2872 14356 2924 14408
rect 4068 14356 4120 14408
rect 4620 14356 4672 14408
rect 4804 14356 4856 14408
rect 7380 14356 7432 14408
rect 7564 14356 7616 14408
rect 9496 14424 9548 14476
rect 9864 14492 9916 14544
rect 10508 14492 10560 14544
rect 11060 14492 11112 14544
rect 13544 14492 13596 14544
rect 18788 14492 18840 14544
rect 19064 14492 19116 14544
rect 22928 14560 22980 14612
rect 10140 14424 10192 14476
rect 10324 14424 10376 14476
rect 12716 14424 12768 14476
rect 13452 14424 13504 14476
rect 15476 14424 15528 14476
rect 16120 14424 16172 14476
rect 8484 14356 8536 14408
rect 9036 14356 9088 14408
rect 9404 14356 9456 14408
rect 9772 14356 9824 14408
rect 10876 14356 10928 14408
rect 11796 14356 11848 14408
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 4160 14288 4212 14340
rect 4896 14288 4948 14340
rect 6276 14288 6328 14340
rect 4344 14263 4396 14272
rect 4344 14229 4353 14263
rect 4353 14229 4387 14263
rect 4387 14229 4396 14263
rect 4344 14220 4396 14229
rect 4528 14220 4580 14272
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 9864 14220 9916 14272
rect 10140 14220 10192 14272
rect 10692 14220 10744 14272
rect 12256 14220 12308 14272
rect 12716 14288 12768 14340
rect 20812 14356 20864 14408
rect 17040 14288 17092 14340
rect 17224 14288 17276 14340
rect 17592 14288 17644 14340
rect 19156 14288 19208 14340
rect 22284 14467 22336 14476
rect 22284 14433 22293 14467
rect 22293 14433 22327 14467
rect 22327 14433 22336 14467
rect 22284 14424 22336 14433
rect 22652 14424 22704 14476
rect 26608 14424 26660 14476
rect 21456 14288 21508 14340
rect 23572 14288 23624 14340
rect 13912 14220 13964 14272
rect 15108 14220 15160 14272
rect 15200 14220 15252 14272
rect 19432 14220 19484 14272
rect 21640 14220 21692 14272
rect 22100 14220 22152 14272
rect 24860 14356 24912 14408
rect 25228 14356 25280 14408
rect 25780 14356 25832 14408
rect 27528 14356 27580 14408
rect 35808 14356 35860 14408
rect 23940 14220 23992 14272
rect 25688 14288 25740 14340
rect 26148 14331 26200 14340
rect 26148 14297 26157 14331
rect 26157 14297 26191 14331
rect 26191 14297 26200 14331
rect 26148 14288 26200 14297
rect 24860 14220 24912 14272
rect 25136 14220 25188 14272
rect 25780 14263 25832 14272
rect 25780 14229 25789 14263
rect 25789 14229 25823 14263
rect 25823 14229 25832 14263
rect 25780 14220 25832 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 4620 14016 4672 14068
rect 6368 14016 6420 14068
rect 4528 13948 4580 14000
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 8668 14016 8720 14068
rect 10048 13948 10100 14000
rect 3700 13923 3752 13932
rect 3700 13889 3709 13923
rect 3709 13889 3743 13923
rect 3743 13889 3752 13923
rect 3700 13880 3752 13889
rect 5172 13880 5224 13932
rect 11060 14016 11112 14068
rect 11152 13948 11204 14000
rect 5724 13855 5776 13864
rect 5724 13821 5733 13855
rect 5733 13821 5767 13855
rect 5767 13821 5776 13855
rect 5724 13812 5776 13821
rect 7104 13812 7156 13864
rect 7564 13855 7616 13864
rect 7564 13821 7573 13855
rect 7573 13821 7607 13855
rect 7607 13821 7616 13855
rect 7564 13812 7616 13821
rect 8484 13812 8536 13864
rect 5908 13744 5960 13796
rect 7288 13744 7340 13796
rect 8208 13744 8260 13796
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 9588 13812 9640 13864
rect 11244 13880 11296 13932
rect 11612 13880 11664 13932
rect 11704 13880 11756 13932
rect 14832 14059 14884 14068
rect 14832 14025 14841 14059
rect 14841 14025 14875 14059
rect 14875 14025 14884 14059
rect 14832 14016 14884 14025
rect 18328 14016 18380 14068
rect 18420 14016 18472 14068
rect 19248 14016 19300 14068
rect 21088 14016 21140 14068
rect 23572 14016 23624 14068
rect 25780 14016 25832 14068
rect 15292 13948 15344 14000
rect 16396 13948 16448 14000
rect 17408 13991 17460 14000
rect 17408 13957 17417 13991
rect 17417 13957 17451 13991
rect 17451 13957 17460 13991
rect 17408 13948 17460 13957
rect 17684 13948 17736 14000
rect 18696 13948 18748 14000
rect 22100 13948 22152 14000
rect 22192 13948 22244 14000
rect 12808 13880 12860 13932
rect 15384 13880 15436 13932
rect 16212 13880 16264 13932
rect 18788 13880 18840 13932
rect 18972 13880 19024 13932
rect 20076 13880 20128 13932
rect 12164 13744 12216 13796
rect 14464 13812 14516 13864
rect 15200 13812 15252 13864
rect 16028 13855 16080 13864
rect 16028 13821 16037 13855
rect 16037 13821 16071 13855
rect 16071 13821 16080 13855
rect 16028 13812 16080 13821
rect 7564 13676 7616 13728
rect 8300 13676 8352 13728
rect 10600 13676 10652 13728
rect 11152 13676 11204 13728
rect 12440 13676 12492 13728
rect 15384 13676 15436 13728
rect 16304 13812 16356 13864
rect 17040 13812 17092 13864
rect 21364 13880 21416 13932
rect 22928 13948 22980 14000
rect 24860 13948 24912 14000
rect 19800 13744 19852 13796
rect 22744 13855 22796 13864
rect 22744 13821 22753 13855
rect 22753 13821 22787 13855
rect 22787 13821 22796 13855
rect 22744 13812 22796 13821
rect 21824 13744 21876 13796
rect 23848 13744 23900 13796
rect 24032 13744 24084 13796
rect 49240 13812 49292 13864
rect 18972 13676 19024 13728
rect 19524 13676 19576 13728
rect 21180 13676 21232 13728
rect 22100 13676 22152 13728
rect 25136 13676 25188 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 8208 13404 8260 13456
rect 13452 13472 13504 13524
rect 15016 13472 15068 13524
rect 17408 13472 17460 13524
rect 21364 13472 21416 13524
rect 4804 13336 4856 13388
rect 8300 13336 8352 13388
rect 14096 13404 14148 13456
rect 15660 13404 15712 13456
rect 22468 13404 22520 13456
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 14648 13336 14700 13388
rect 15844 13336 15896 13388
rect 17040 13336 17092 13388
rect 17500 13336 17552 13388
rect 22192 13336 22244 13388
rect 23388 13336 23440 13388
rect 23480 13379 23532 13388
rect 23480 13345 23489 13379
rect 23489 13345 23523 13379
rect 23523 13345 23532 13379
rect 23480 13336 23532 13345
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 19340 13268 19392 13320
rect 23020 13268 23072 13320
rect 4528 13200 4580 13252
rect 6276 13200 6328 13252
rect 6644 13200 6696 13252
rect 7104 13200 7156 13252
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 7380 13132 7432 13184
rect 8576 13132 8628 13184
rect 10692 13175 10744 13184
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 10692 13132 10744 13141
rect 12348 13200 12400 13252
rect 12532 13200 12584 13252
rect 12716 13200 12768 13252
rect 13636 13132 13688 13184
rect 15016 13200 15068 13252
rect 15200 13132 15252 13184
rect 15384 13132 15436 13184
rect 16488 13175 16540 13184
rect 16488 13141 16497 13175
rect 16497 13141 16531 13175
rect 16531 13141 16540 13175
rect 16488 13132 16540 13141
rect 17684 13200 17736 13252
rect 18972 13200 19024 13252
rect 21640 13200 21692 13252
rect 24124 13200 24176 13252
rect 24584 13243 24636 13252
rect 24584 13209 24593 13243
rect 24593 13209 24627 13243
rect 24627 13209 24636 13243
rect 24584 13200 24636 13209
rect 26884 13200 26936 13252
rect 18420 13132 18472 13184
rect 18788 13132 18840 13184
rect 28540 13132 28592 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 3516 12971 3568 12980
rect 3516 12937 3525 12971
rect 3525 12937 3559 12971
rect 3559 12937 3568 12971
rect 3516 12928 3568 12937
rect 5724 12928 5776 12980
rect 7380 12971 7432 12980
rect 7380 12937 7389 12971
rect 7389 12937 7423 12971
rect 7423 12937 7432 12971
rect 7380 12928 7432 12937
rect 7564 12928 7616 12980
rect 8300 12928 8352 12980
rect 9312 12928 9364 12980
rect 10968 12928 11020 12980
rect 2780 12903 2832 12912
rect 2780 12869 2789 12903
rect 2789 12869 2823 12903
rect 2823 12869 2832 12903
rect 2780 12860 2832 12869
rect 3792 12860 3844 12912
rect 4436 12903 4488 12912
rect 4436 12869 4445 12903
rect 4445 12869 4479 12903
rect 4479 12869 4488 12903
rect 4436 12860 4488 12869
rect 4528 12860 4580 12912
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 4528 12767 4580 12776
rect 4528 12733 4537 12767
rect 4537 12733 4571 12767
rect 4571 12733 4580 12767
rect 4528 12724 4580 12733
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 5540 12724 5592 12776
rect 6736 12792 6788 12844
rect 8484 12903 8536 12912
rect 8484 12869 8493 12903
rect 8493 12869 8527 12903
rect 8527 12869 8536 12903
rect 8484 12860 8536 12869
rect 8760 12860 8812 12912
rect 10232 12903 10284 12912
rect 10232 12869 10241 12903
rect 10241 12869 10275 12903
rect 10275 12869 10284 12903
rect 10232 12860 10284 12869
rect 12072 12860 12124 12912
rect 5816 12656 5868 12708
rect 6276 12724 6328 12776
rect 9864 12792 9916 12844
rect 12808 12792 12860 12844
rect 14740 12792 14792 12844
rect 16028 12928 16080 12980
rect 15016 12903 15068 12912
rect 15016 12869 15025 12903
rect 15025 12869 15059 12903
rect 15059 12869 15068 12903
rect 15016 12860 15068 12869
rect 18880 12860 18932 12912
rect 19156 12903 19208 12912
rect 19156 12869 19165 12903
rect 19165 12869 19199 12903
rect 19199 12869 19208 12903
rect 19156 12860 19208 12869
rect 21088 12903 21140 12912
rect 21088 12869 21097 12903
rect 21097 12869 21131 12903
rect 21131 12869 21140 12903
rect 21088 12860 21140 12869
rect 17868 12792 17920 12844
rect 20720 12792 20772 12844
rect 22008 12928 22060 12980
rect 23480 12928 23532 12980
rect 22100 12792 22152 12844
rect 22192 12792 22244 12844
rect 23020 12835 23072 12844
rect 23020 12801 23029 12835
rect 23029 12801 23063 12835
rect 23063 12801 23072 12835
rect 23020 12792 23072 12801
rect 24400 12792 24452 12844
rect 5264 12631 5316 12640
rect 5264 12597 5273 12631
rect 5273 12597 5307 12631
rect 5307 12597 5316 12631
rect 5264 12588 5316 12597
rect 8484 12588 8536 12640
rect 9128 12588 9180 12640
rect 9680 12588 9732 12640
rect 14464 12767 14516 12776
rect 14464 12733 14473 12767
rect 14473 12733 14507 12767
rect 14507 12733 14516 12767
rect 14464 12724 14516 12733
rect 15844 12767 15896 12776
rect 15844 12733 15853 12767
rect 15853 12733 15887 12767
rect 15887 12733 15896 12767
rect 15844 12724 15896 12733
rect 15936 12724 15988 12776
rect 16304 12724 16356 12776
rect 18788 12724 18840 12776
rect 12624 12588 12676 12640
rect 15384 12656 15436 12708
rect 17500 12656 17552 12708
rect 20076 12724 20128 12776
rect 21456 12724 21508 12776
rect 23940 12724 23992 12776
rect 22560 12656 22612 12708
rect 13360 12588 13412 12640
rect 13820 12631 13872 12640
rect 13820 12597 13829 12631
rect 13829 12597 13863 12631
rect 13863 12597 13872 12631
rect 13820 12588 13872 12597
rect 15476 12588 15528 12640
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 23940 12588 23992 12640
rect 24400 12588 24452 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 4528 12384 4580 12436
rect 6092 12384 6144 12436
rect 6368 12384 6420 12436
rect 7380 12384 7432 12436
rect 7472 12384 7524 12436
rect 7748 12384 7800 12436
rect 10692 12384 10744 12436
rect 11980 12384 12032 12436
rect 15752 12384 15804 12436
rect 18420 12384 18472 12436
rect 21824 12427 21876 12436
rect 21824 12393 21833 12427
rect 21833 12393 21867 12427
rect 21867 12393 21876 12427
rect 21824 12384 21876 12393
rect 3424 12359 3476 12368
rect 3424 12325 3433 12359
rect 3433 12325 3467 12359
rect 3467 12325 3476 12359
rect 3424 12316 3476 12325
rect 1584 12291 1636 12300
rect 1584 12257 1593 12291
rect 1593 12257 1627 12291
rect 1627 12257 1636 12291
rect 1584 12248 1636 12257
rect 5356 12316 5408 12368
rect 4712 12291 4764 12300
rect 4712 12257 4721 12291
rect 4721 12257 4755 12291
rect 4755 12257 4764 12291
rect 4712 12248 4764 12257
rect 7656 12248 7708 12300
rect 2872 12180 2924 12232
rect 3148 12180 3200 12232
rect 4344 12180 4396 12232
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 4804 12180 4856 12232
rect 10416 12316 10468 12368
rect 8576 12248 8628 12300
rect 9312 12248 9364 12300
rect 15292 12316 15344 12368
rect 8392 12180 8444 12232
rect 8852 12180 8904 12232
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 10784 12291 10836 12300
rect 10784 12257 10793 12291
rect 10793 12257 10827 12291
rect 10827 12257 10836 12291
rect 10784 12248 10836 12257
rect 12348 12291 12400 12300
rect 12348 12257 12357 12291
rect 12357 12257 12391 12291
rect 12391 12257 12400 12291
rect 12348 12248 12400 12257
rect 14832 12248 14884 12300
rect 15844 12248 15896 12300
rect 16672 12248 16724 12300
rect 17316 12248 17368 12300
rect 2780 12155 2832 12164
rect 2780 12121 2789 12155
rect 2789 12121 2823 12155
rect 2823 12121 2832 12155
rect 2780 12112 2832 12121
rect 2044 12044 2096 12096
rect 5724 12112 5776 12164
rect 6644 12112 6696 12164
rect 6920 12112 6972 12164
rect 11980 12180 12032 12232
rect 16120 12180 16172 12232
rect 9680 12112 9732 12164
rect 15016 12112 15068 12164
rect 15108 12155 15160 12164
rect 15108 12121 15117 12155
rect 15117 12121 15151 12155
rect 15151 12121 15160 12155
rect 15108 12112 15160 12121
rect 15384 12112 15436 12164
rect 16488 12112 16540 12164
rect 17040 12112 17092 12164
rect 20076 12291 20128 12300
rect 20076 12257 20085 12291
rect 20085 12257 20119 12291
rect 20119 12257 20128 12291
rect 20076 12248 20128 12257
rect 21916 12248 21968 12300
rect 22192 12180 22244 12232
rect 7196 12044 7248 12096
rect 12440 12044 12492 12096
rect 12624 12044 12676 12096
rect 13360 12087 13412 12096
rect 13360 12053 13369 12087
rect 13369 12053 13403 12087
rect 13403 12053 13412 12087
rect 13360 12044 13412 12053
rect 16856 12044 16908 12096
rect 17316 12044 17368 12096
rect 20720 12044 20772 12096
rect 21640 12044 21692 12096
rect 23940 12112 23992 12164
rect 24032 12087 24084 12096
rect 24032 12053 24041 12087
rect 24041 12053 24075 12087
rect 24075 12053 24084 12087
rect 24032 12044 24084 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 3148 11840 3200 11892
rect 4620 11840 4672 11892
rect 6920 11840 6972 11892
rect 7380 11840 7432 11892
rect 7932 11840 7984 11892
rect 8484 11840 8536 11892
rect 11980 11883 12032 11892
rect 11980 11849 11989 11883
rect 11989 11849 12023 11883
rect 12023 11849 12032 11883
rect 11980 11840 12032 11849
rect 12164 11840 12216 11892
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 16948 11840 17000 11892
rect 17868 11840 17920 11892
rect 18512 11883 18564 11892
rect 18512 11849 18521 11883
rect 18521 11849 18555 11883
rect 18555 11849 18564 11883
rect 18512 11840 18564 11849
rect 20260 11840 20312 11892
rect 7288 11772 7340 11824
rect 9680 11772 9732 11824
rect 12532 11772 12584 11824
rect 20812 11840 20864 11892
rect 20720 11772 20772 11824
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 2412 11747 2464 11756
rect 2412 11713 2421 11747
rect 2421 11713 2455 11747
rect 2455 11713 2464 11747
rect 2412 11704 2464 11713
rect 4344 11747 4396 11756
rect 4344 11713 4353 11747
rect 4353 11713 4387 11747
rect 4387 11713 4396 11747
rect 4344 11704 4396 11713
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 6920 11704 6972 11756
rect 7196 11704 7248 11756
rect 8760 11704 8812 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11980 11704 12032 11756
rect 12164 11704 12216 11756
rect 12808 11704 12860 11756
rect 15936 11747 15988 11756
rect 15936 11713 15945 11747
rect 15945 11713 15979 11747
rect 15979 11713 15988 11747
rect 15936 11704 15988 11713
rect 16120 11704 16172 11756
rect 19064 11704 19116 11756
rect 7288 11679 7340 11688
rect 5724 11568 5776 11620
rect 7288 11645 7297 11679
rect 7297 11645 7331 11679
rect 7331 11645 7340 11679
rect 7288 11636 7340 11645
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 7196 11568 7248 11620
rect 3700 11500 3752 11552
rect 6644 11500 6696 11552
rect 7380 11500 7432 11552
rect 11520 11636 11572 11688
rect 11888 11636 11940 11688
rect 12164 11568 12216 11620
rect 9864 11500 9916 11552
rect 10140 11500 10192 11552
rect 12348 11500 12400 11552
rect 15660 11636 15712 11688
rect 17408 11636 17460 11688
rect 16856 11568 16908 11620
rect 17224 11568 17276 11620
rect 17592 11636 17644 11688
rect 19708 11679 19760 11688
rect 19708 11645 19717 11679
rect 19717 11645 19751 11679
rect 19751 11645 19760 11679
rect 19708 11636 19760 11645
rect 24032 11840 24084 11892
rect 22652 11815 22704 11824
rect 22652 11781 22661 11815
rect 22661 11781 22695 11815
rect 22695 11781 22704 11815
rect 22652 11772 22704 11781
rect 23940 11772 23992 11824
rect 22192 11636 22244 11688
rect 23296 11636 23348 11688
rect 25136 11840 25188 11892
rect 14556 11500 14608 11552
rect 14740 11500 14792 11552
rect 17040 11500 17092 11552
rect 21456 11543 21508 11552
rect 21456 11509 21465 11543
rect 21465 11509 21499 11543
rect 21499 11509 21508 11543
rect 21456 11500 21508 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 2596 11339 2648 11348
rect 2596 11305 2605 11339
rect 2605 11305 2639 11339
rect 2639 11305 2648 11339
rect 2596 11296 2648 11305
rect 2504 11228 2556 11280
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 3976 11092 4028 11144
rect 5540 11296 5592 11348
rect 5724 11296 5776 11348
rect 7748 11296 7800 11348
rect 10232 11296 10284 11348
rect 11888 11296 11940 11348
rect 12256 11296 12308 11348
rect 14740 11296 14792 11348
rect 6644 11228 6696 11280
rect 4804 11203 4856 11212
rect 4804 11169 4813 11203
rect 4813 11169 4847 11203
rect 4847 11169 4856 11203
rect 4804 11160 4856 11169
rect 5816 11160 5868 11212
rect 7840 11160 7892 11212
rect 9312 11228 9364 11280
rect 8392 11092 8444 11144
rect 6552 11024 6604 11076
rect 7288 10956 7340 11008
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 9220 11092 9272 11144
rect 10140 10956 10192 11008
rect 11152 11228 11204 11280
rect 16488 11339 16540 11348
rect 16488 11305 16497 11339
rect 16497 11305 16531 11339
rect 16531 11305 16540 11339
rect 16488 11296 16540 11305
rect 18788 11296 18840 11348
rect 18880 11339 18932 11348
rect 18880 11305 18889 11339
rect 18889 11305 18923 11339
rect 18923 11305 18932 11339
rect 18880 11296 18932 11305
rect 10784 11067 10836 11076
rect 10784 11033 10793 11067
rect 10793 11033 10827 11067
rect 10827 11033 10836 11067
rect 10784 11024 10836 11033
rect 11060 11024 11112 11076
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 12256 11160 12308 11212
rect 14556 11160 14608 11212
rect 15108 11160 15160 11212
rect 22652 11203 22704 11212
rect 22652 11169 22661 11203
rect 22661 11169 22695 11203
rect 22695 11169 22704 11203
rect 22652 11160 22704 11169
rect 26884 11160 26936 11212
rect 16856 11092 16908 11144
rect 19156 11092 19208 11144
rect 11888 11024 11940 11076
rect 11980 10956 12032 11008
rect 12532 11024 12584 11076
rect 15016 11067 15068 11076
rect 15016 11033 15025 11067
rect 15025 11033 15059 11067
rect 15059 11033 15068 11067
rect 15016 11024 15068 11033
rect 15292 11024 15344 11076
rect 17868 11024 17920 11076
rect 19708 11024 19760 11076
rect 21180 11067 21232 11076
rect 21180 11033 21189 11067
rect 21189 11033 21223 11067
rect 21223 11033 21232 11067
rect 21180 11024 21232 11033
rect 15200 10956 15252 11008
rect 15660 10956 15712 11008
rect 19340 10956 19392 11008
rect 20720 10956 20772 11008
rect 28356 11024 28408 11076
rect 30104 11024 30156 11076
rect 31668 11024 31720 11076
rect 47860 11024 47912 11076
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 3884 10795 3936 10804
rect 3884 10761 3893 10795
rect 3893 10761 3927 10795
rect 3927 10761 3936 10795
rect 3884 10752 3936 10761
rect 4344 10752 4396 10804
rect 6920 10752 6972 10804
rect 4252 10684 4304 10736
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 4436 10616 4488 10668
rect 4528 10659 4580 10668
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 4712 10727 4764 10736
rect 4712 10693 4721 10727
rect 4721 10693 4755 10727
rect 4755 10693 4764 10727
rect 4712 10684 4764 10693
rect 7196 10752 7248 10804
rect 11520 10752 11572 10804
rect 12164 10752 12216 10804
rect 15568 10752 15620 10804
rect 5264 10616 5316 10668
rect 5908 10591 5960 10600
rect 5908 10557 5917 10591
rect 5917 10557 5951 10591
rect 5951 10557 5960 10591
rect 5908 10548 5960 10557
rect 6920 10480 6972 10532
rect 6736 10455 6788 10464
rect 6736 10421 6745 10455
rect 6745 10421 6779 10455
rect 6779 10421 6788 10455
rect 6736 10412 6788 10421
rect 9404 10727 9456 10736
rect 9404 10693 9413 10727
rect 9413 10693 9447 10727
rect 9447 10693 9456 10727
rect 9404 10684 9456 10693
rect 8760 10616 8812 10668
rect 9588 10616 9640 10668
rect 11244 10616 11296 10668
rect 12348 10684 12400 10736
rect 12624 10684 12676 10736
rect 15752 10684 15804 10736
rect 14280 10616 14332 10668
rect 17408 10752 17460 10804
rect 17868 10684 17920 10736
rect 7380 10591 7432 10600
rect 7380 10557 7389 10591
rect 7389 10557 7423 10591
rect 7423 10557 7432 10591
rect 7380 10548 7432 10557
rect 7380 10412 7432 10464
rect 10324 10548 10376 10600
rect 11152 10548 11204 10600
rect 9680 10480 9732 10532
rect 7840 10412 7892 10464
rect 8024 10412 8076 10464
rect 15660 10480 15712 10532
rect 11980 10412 12032 10464
rect 15200 10412 15252 10464
rect 16028 10412 16080 10464
rect 16304 10548 16356 10600
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 17500 10659 17552 10668
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 17316 10548 17368 10600
rect 17040 10480 17092 10532
rect 21456 10752 21508 10804
rect 20720 10684 20772 10736
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 22652 10548 22704 10600
rect 18788 10480 18840 10532
rect 19432 10412 19484 10464
rect 24860 10412 24912 10464
rect 32864 10412 32916 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 1124 10140 1176 10192
rect 940 10072 992 10124
rect 2228 10072 2280 10124
rect 7840 10072 7892 10124
rect 2780 10004 2832 10056
rect 6460 10004 6512 10056
rect 8760 10004 8812 10056
rect 9036 10004 9088 10056
rect 12808 10208 12860 10260
rect 14188 10140 14240 10192
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 7196 9936 7248 9988
rect 8392 9936 8444 9988
rect 9496 9936 9548 9988
rect 11244 10115 11296 10124
rect 11244 10081 11253 10115
rect 11253 10081 11287 10115
rect 11287 10081 11296 10115
rect 11244 10072 11296 10081
rect 11520 10115 11572 10124
rect 11520 10081 11529 10115
rect 11529 10081 11563 10115
rect 11563 10081 11572 10115
rect 11520 10072 11572 10081
rect 12256 10072 12308 10124
rect 12900 10072 12952 10124
rect 12624 10004 12676 10056
rect 13084 10072 13136 10124
rect 15016 10208 15068 10260
rect 17592 10208 17644 10260
rect 19248 10208 19300 10260
rect 15844 10140 15896 10192
rect 16948 10140 17000 10192
rect 14556 10115 14608 10124
rect 14556 10081 14565 10115
rect 14565 10081 14599 10115
rect 14599 10081 14608 10115
rect 14556 10072 14608 10081
rect 14832 10115 14884 10124
rect 14832 10081 14841 10115
rect 14841 10081 14875 10115
rect 14875 10081 14884 10115
rect 14832 10072 14884 10081
rect 14924 10072 14976 10124
rect 17040 10072 17092 10124
rect 13176 10004 13228 10056
rect 16856 10004 16908 10056
rect 19708 10072 19760 10124
rect 13452 9936 13504 9988
rect 6736 9868 6788 9920
rect 8484 9868 8536 9920
rect 9680 9868 9732 9920
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 12348 9868 12400 9920
rect 14740 9936 14792 9988
rect 15292 9936 15344 9988
rect 13728 9868 13780 9920
rect 17408 9979 17460 9988
rect 17408 9945 17417 9979
rect 17417 9945 17451 9979
rect 17451 9945 17460 9979
rect 17408 9936 17460 9945
rect 17868 9936 17920 9988
rect 20720 9936 20772 9988
rect 23296 10208 23348 10260
rect 22100 10072 22152 10124
rect 23848 10072 23900 10124
rect 21180 9911 21232 9920
rect 21180 9877 21189 9911
rect 21189 9877 21223 9911
rect 21223 9877 21232 9911
rect 21180 9868 21232 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 6920 9707 6972 9716
rect 6920 9673 6929 9707
rect 6929 9673 6963 9707
rect 6963 9673 6972 9707
rect 6920 9664 6972 9673
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 3424 9528 3476 9580
rect 6092 9596 6144 9648
rect 6276 9596 6328 9648
rect 5632 9528 5684 9580
rect 7012 9528 7064 9580
rect 5908 9460 5960 9512
rect 6736 9460 6788 9512
rect 8392 9639 8444 9648
rect 8392 9605 8401 9639
rect 8401 9605 8435 9639
rect 8435 9605 8444 9639
rect 8392 9596 8444 9605
rect 9036 9596 9088 9648
rect 9864 9664 9916 9716
rect 10324 9707 10376 9716
rect 10324 9673 10333 9707
rect 10333 9673 10367 9707
rect 10367 9673 10376 9707
rect 10324 9664 10376 9673
rect 12164 9664 12216 9716
rect 10784 9639 10836 9648
rect 10784 9605 10793 9639
rect 10793 9605 10827 9639
rect 10827 9605 10836 9639
rect 10784 9596 10836 9605
rect 3792 9392 3844 9444
rect 7840 9460 7892 9512
rect 9864 9528 9916 9580
rect 11244 9528 11296 9580
rect 13452 9528 13504 9580
rect 13176 9460 13228 9512
rect 13636 9460 13688 9512
rect 17224 9596 17276 9648
rect 17408 9596 17460 9648
rect 18420 9596 18472 9648
rect 23572 9596 23624 9648
rect 14464 9571 14516 9580
rect 14464 9537 14473 9571
rect 14473 9537 14507 9571
rect 14507 9537 14516 9571
rect 14464 9528 14516 9537
rect 16120 9528 16172 9580
rect 19432 9571 19484 9580
rect 19432 9537 19441 9571
rect 19441 9537 19475 9571
rect 19475 9537 19484 9571
rect 19432 9528 19484 9537
rect 27436 9528 27488 9580
rect 14832 9460 14884 9512
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 18328 9460 18380 9512
rect 19248 9460 19300 9512
rect 21180 9460 21232 9512
rect 22560 9460 22612 9512
rect 11428 9392 11480 9444
rect 19616 9392 19668 9444
rect 10140 9324 10192 9376
rect 10324 9324 10376 9376
rect 14740 9324 14792 9376
rect 16304 9324 16356 9376
rect 31668 9324 31720 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 4068 9120 4120 9172
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 5172 9163 5224 9172
rect 5172 9129 5181 9163
rect 5181 9129 5215 9163
rect 5215 9129 5224 9163
rect 5172 9120 5224 9129
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 4528 9052 4580 9104
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 4988 8984 5040 9036
rect 940 8916 992 8968
rect 3332 8916 3384 8968
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 8392 9052 8444 9104
rect 9864 9052 9916 9104
rect 7104 8984 7156 9036
rect 9128 9027 9180 9036
rect 9128 8993 9137 9027
rect 9137 8993 9171 9027
rect 9171 8993 9180 9027
rect 9128 8984 9180 8993
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 9680 8984 9732 9036
rect 12256 9027 12308 9036
rect 12256 8993 12265 9027
rect 12265 8993 12299 9027
rect 12299 8993 12308 9027
rect 12256 8984 12308 8993
rect 15476 9052 15528 9104
rect 17408 9052 17460 9104
rect 22100 9052 22152 9104
rect 13820 8984 13872 9036
rect 14740 9027 14792 9036
rect 14740 8993 14749 9027
rect 14749 8993 14783 9027
rect 14783 8993 14792 9027
rect 14740 8984 14792 8993
rect 14924 9027 14976 9036
rect 14924 8993 14933 9027
rect 14933 8993 14967 9027
rect 14967 8993 14976 9027
rect 14924 8984 14976 8993
rect 16856 8984 16908 9036
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 10232 8916 10284 8968
rect 12072 8916 12124 8968
rect 12440 8916 12492 8968
rect 18420 8916 18472 8968
rect 8852 8848 8904 8900
rect 6460 8780 6512 8832
rect 6736 8780 6788 8832
rect 10324 8848 10376 8900
rect 9864 8780 9916 8832
rect 13084 8848 13136 8900
rect 11980 8823 12032 8832
rect 11980 8789 11989 8823
rect 11989 8789 12023 8823
rect 12023 8789 12032 8823
rect 11980 8780 12032 8789
rect 12072 8823 12124 8832
rect 12072 8789 12081 8823
rect 12081 8789 12115 8823
rect 12115 8789 12124 8823
rect 12072 8780 12124 8789
rect 12624 8780 12676 8832
rect 13636 8780 13688 8832
rect 15936 8780 15988 8832
rect 16304 8891 16356 8900
rect 16304 8857 16313 8891
rect 16313 8857 16347 8891
rect 16347 8857 16356 8891
rect 16304 8848 16356 8857
rect 19432 8848 19484 8900
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 3608 8576 3660 8628
rect 4436 8576 4488 8628
rect 11796 8576 11848 8628
rect 12808 8576 12860 8628
rect 13084 8619 13136 8628
rect 13084 8585 13093 8619
rect 13093 8585 13127 8619
rect 13127 8585 13136 8619
rect 13084 8576 13136 8585
rect 7564 8508 7616 8560
rect 2872 8440 2924 8492
rect 3516 8440 3568 8492
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 8944 8483 8996 8492
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 11336 8508 11388 8560
rect 9956 8440 10008 8492
rect 2044 8372 2096 8424
rect 1676 8304 1728 8356
rect 4252 8304 4304 8356
rect 9220 8372 9272 8424
rect 13360 8440 13412 8492
rect 15384 8440 15436 8492
rect 16948 8440 17000 8492
rect 11244 8372 11296 8424
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12440 8372 12492 8381
rect 11152 8304 11204 8356
rect 13728 8415 13780 8424
rect 13728 8381 13737 8415
rect 13737 8381 13771 8415
rect 13771 8381 13780 8415
rect 13728 8372 13780 8381
rect 18328 8372 18380 8424
rect 14280 8347 14332 8356
rect 14280 8313 14289 8347
rect 14289 8313 14323 8347
rect 14323 8313 14332 8347
rect 14280 8304 14332 8313
rect 10232 8236 10284 8288
rect 11060 8236 11112 8288
rect 14004 8236 14056 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 2136 8032 2188 8084
rect 8668 8032 8720 8084
rect 9588 8075 9640 8084
rect 9588 8041 9597 8075
rect 9597 8041 9631 8075
rect 9631 8041 9640 8075
rect 9588 8032 9640 8041
rect 11060 8032 11112 8084
rect 12716 8075 12768 8084
rect 12716 8041 12725 8075
rect 12725 8041 12759 8075
rect 12759 8041 12768 8075
rect 12716 8032 12768 8041
rect 13360 8075 13412 8084
rect 13360 8041 13369 8075
rect 13369 8041 13403 8075
rect 13403 8041 13412 8075
rect 13360 8032 13412 8041
rect 23940 8075 23992 8084
rect 23940 8041 23949 8075
rect 23949 8041 23983 8075
rect 23983 8041 23992 8075
rect 23940 8032 23992 8041
rect 28356 8032 28408 8084
rect 1308 7896 1360 7948
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 2780 7828 2832 7880
rect 8484 7896 8536 7948
rect 12440 7964 12492 8016
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 10968 7939 11020 7948
rect 10968 7905 10977 7939
rect 10977 7905 11011 7939
rect 11011 7905 11020 7939
rect 10968 7896 11020 7905
rect 11520 7896 11572 7948
rect 15200 8007 15252 8016
rect 15200 7973 15209 8007
rect 15209 7973 15243 8007
rect 15243 7973 15252 8007
rect 15200 7964 15252 7973
rect 22192 7939 22244 7948
rect 22192 7905 22201 7939
rect 22201 7905 22235 7939
rect 22235 7905 22244 7939
rect 22192 7896 22244 7905
rect 8300 7760 8352 7812
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 16672 7760 16724 7812
rect 13452 7692 13504 7744
rect 22468 7803 22520 7812
rect 22468 7769 22477 7803
rect 22477 7769 22511 7803
rect 22511 7769 22520 7803
rect 22468 7760 22520 7769
rect 23848 7760 23900 7812
rect 22560 7692 22612 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 8392 7488 8444 7540
rect 9864 7488 9916 7540
rect 10048 7488 10100 7540
rect 3700 7420 3752 7472
rect 1400 7352 1452 7404
rect 2780 7352 2832 7404
rect 9312 7352 9364 7404
rect 11980 7352 12032 7404
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 10140 7327 10192 7336
rect 10140 7293 10149 7327
rect 10149 7293 10183 7327
rect 10183 7293 10192 7327
rect 10140 7284 10192 7293
rect 7656 7216 7708 7268
rect 15568 7216 15620 7268
rect 16488 7148 16540 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 23940 6944 23992 6996
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 1216 6672 1268 6724
rect 2872 6740 2924 6792
rect 20904 6740 20956 6792
rect 27436 6740 27488 6792
rect 1676 6604 1728 6656
rect 6644 6672 6696 6724
rect 7288 6604 7340 6656
rect 22100 6604 22152 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 22560 6264 22612 6316
rect 940 6196 992 6248
rect 11704 6196 11756 6248
rect 24768 6060 24820 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 22468 5856 22520 5908
rect 12624 5788 12676 5840
rect 15476 5720 15528 5772
rect 16856 5720 16908 5772
rect 22100 5720 22152 5772
rect 24768 5763 24820 5772
rect 24768 5729 24777 5763
rect 24777 5729 24811 5763
rect 24811 5729 24820 5763
rect 24768 5720 24820 5729
rect 28908 5720 28960 5772
rect 940 5652 992 5704
rect 10600 5652 10652 5704
rect 20904 5695 20956 5704
rect 20904 5661 20913 5695
rect 20913 5661 20947 5695
rect 20947 5661 20956 5695
rect 20904 5652 20956 5661
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 18420 5584 18472 5636
rect 25504 5584 25556 5636
rect 17040 5516 17092 5568
rect 21364 5559 21416 5568
rect 21364 5525 21373 5559
rect 21373 5525 21407 5559
rect 21407 5525 21416 5559
rect 21364 5516 21416 5525
rect 27068 5627 27120 5636
rect 27068 5593 27077 5627
rect 27077 5593 27111 5627
rect 27111 5593 27120 5627
rect 27068 5584 27120 5593
rect 28724 5627 28776 5636
rect 28724 5593 28733 5627
rect 28733 5593 28767 5627
rect 28767 5593 28776 5627
rect 28724 5584 28776 5593
rect 27620 5516 27672 5568
rect 28356 5516 28408 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 27068 5312 27120 5364
rect 940 5176 992 5228
rect 7380 5176 7432 5228
rect 15568 5219 15620 5228
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 16488 5176 16540 5228
rect 15476 5108 15528 5160
rect 21364 5176 21416 5228
rect 22100 5219 22152 5228
rect 22100 5185 22144 5219
rect 22144 5185 22152 5219
rect 22100 5176 22152 5185
rect 17684 5151 17736 5160
rect 17684 5117 17693 5151
rect 17693 5117 17727 5151
rect 17727 5117 17736 5151
rect 17684 5108 17736 5117
rect 28816 5151 28868 5160
rect 28816 5117 28825 5151
rect 28825 5117 28859 5151
rect 28859 5117 28868 5151
rect 28816 5108 28868 5117
rect 30380 5108 30432 5160
rect 31392 5108 31444 5160
rect 33508 5040 33560 5092
rect 17868 4972 17920 5024
rect 20536 4972 20588 5024
rect 25964 4972 26016 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 17408 4768 17460 4820
rect 28816 4768 28868 4820
rect 940 4632 992 4684
rect 27804 4632 27856 4684
rect 11612 4564 11664 4616
rect 20904 4564 20956 4616
rect 17684 4428 17736 4480
rect 25964 4539 26016 4548
rect 25964 4505 25973 4539
rect 25973 4505 26007 4539
rect 26007 4505 26016 4539
rect 25964 4496 26016 4505
rect 27344 4496 27396 4548
rect 27528 4496 27580 4548
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 1308 4088 1360 4140
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 940 4020 992 4072
rect 9220 4020 9272 4072
rect 10324 3952 10376 4004
rect 2780 3884 2832 3936
rect 6736 3884 6788 3936
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 2780 3680 2832 3732
rect 11152 3680 11204 3732
rect 30380 3680 30432 3732
rect 41420 3680 41472 3732
rect 12072 3612 12124 3664
rect 28724 3612 28776 3664
rect 44088 3612 44140 3664
rect 27528 3544 27580 3596
rect 46756 3544 46808 3596
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 1216 3408 1268 3460
rect 2872 3476 2924 3528
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 28356 3476 28408 3528
rect 49424 3476 49476 3528
rect 17132 3408 17184 3460
rect 38752 3408 38804 3460
rect 2964 3340 3016 3392
rect 11244 3340 11296 3392
rect 11612 3383 11664 3392
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 2964 3136 3016 3188
rect 9772 3136 9824 3188
rect 7196 3068 7248 3120
rect 9036 3068 9088 3120
rect 12624 3111 12676 3120
rect 12624 3077 12633 3111
rect 12633 3077 12667 3111
rect 12667 3077 12676 3111
rect 12624 3068 12676 3077
rect 15476 3068 15528 3120
rect 17684 3068 17736 3120
rect 2780 3000 2832 3052
rect 7840 3000 7892 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 17868 3000 17920 3052
rect 20536 3043 20588 3052
rect 20536 3009 20545 3043
rect 20545 3009 20579 3043
rect 20579 3009 20588 3043
rect 20536 3000 20588 3009
rect 940 2932 992 2984
rect 8024 2932 8076 2984
rect 17408 2932 17460 2984
rect 12532 2864 12584 2916
rect 8300 2796 8352 2848
rect 17500 2796 17552 2848
rect 20076 2796 20128 2848
rect 22008 2796 22060 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 9680 2592 9732 2644
rect 25504 2635 25556 2644
rect 25504 2601 25513 2635
rect 25513 2601 25547 2635
rect 25547 2601 25556 2635
rect 25504 2592 25556 2601
rect 27804 2592 27856 2644
rect 28908 2592 28960 2644
rect 33508 2635 33560 2644
rect 33508 2601 33517 2635
rect 33517 2601 33551 2635
rect 33551 2601 33560 2635
rect 33508 2592 33560 2601
rect 4068 2456 4120 2508
rect 6736 2456 6788 2508
rect 9404 2456 9456 2508
rect 12072 2456 12124 2508
rect 14740 2456 14792 2508
rect 17408 2456 17460 2508
rect 20168 2456 20220 2508
rect 22744 2456 22796 2508
rect 27436 2456 27488 2508
rect 940 2388 992 2440
rect 1768 2388 1820 2440
rect 8300 2388 8352 2440
rect 9772 2388 9824 2440
rect 12532 2388 12584 2440
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 22008 2388 22060 2440
rect 25412 2388 25464 2440
rect 28356 2431 28408 2440
rect 28356 2397 28365 2431
rect 28365 2397 28399 2431
rect 28399 2397 28408 2431
rect 28356 2388 28408 2397
rect 30748 2388 30800 2440
rect 33416 2388 33468 2440
rect 36084 2431 36136 2440
rect 36084 2397 36093 2431
rect 36093 2397 36127 2431
rect 36127 2397 36136 2431
rect 36084 2388 36136 2397
rect 11612 2320 11664 2372
rect 8024 2252 8076 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
<< metal2 >>
rect 2226 26200 2282 27000
rect 2870 26200 2926 27000
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26330 4858 27000
rect 4802 26302 5120 26330
rect 4802 26200 4858 26302
rect 1490 24440 1546 24449
rect 1490 24375 1546 24384
rect 1124 23656 1176 23662
rect 1124 23598 1176 23604
rect 938 10976 994 10985
rect 938 10911 994 10920
rect 952 10130 980 10911
rect 1136 10198 1164 23598
rect 1308 22092 1360 22098
rect 1308 22034 1360 22040
rect 1320 20777 1348 22034
rect 1504 21350 1532 24375
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1492 21344 1544 21350
rect 1492 21286 1544 21292
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1412 18737 1440 19858
rect 1398 18728 1454 18737
rect 1398 18663 1454 18672
rect 1596 18170 1624 23802
rect 1860 23520 1912 23526
rect 1860 23462 1912 23468
rect 1676 23316 1728 23322
rect 1676 23258 1728 23264
rect 1688 22642 1716 23258
rect 1768 23112 1820 23118
rect 1768 23054 1820 23060
rect 1780 22710 1808 23054
rect 1768 22704 1820 22710
rect 1768 22646 1820 22652
rect 1676 22636 1728 22642
rect 1676 22578 1728 22584
rect 1768 21684 1820 21690
rect 1768 21626 1820 21632
rect 1780 19854 1808 21626
rect 1872 20466 1900 23462
rect 2136 21616 2188 21622
rect 2136 21558 2188 21564
rect 2044 21480 2096 21486
rect 2044 21422 2096 21428
rect 1952 21412 2004 21418
rect 1952 21354 2004 21360
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1766 19272 1822 19281
rect 1766 19207 1822 19216
rect 1596 18142 1716 18170
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1216 17740 1268 17746
rect 1216 17682 1268 17688
rect 1228 17105 1256 17682
rect 1308 17128 1360 17134
rect 1214 17096 1270 17105
rect 1308 17070 1360 17076
rect 1214 17031 1270 17040
rect 1320 16697 1348 17070
rect 1306 16688 1362 16697
rect 1306 16623 1362 16632
rect 1596 16574 1624 18022
rect 1688 17882 1716 18142
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1780 17678 1808 19207
rect 1964 18290 1992 21354
rect 2056 19961 2084 21422
rect 2042 19952 2098 19961
rect 2042 19887 2098 19896
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 2056 18329 2084 19246
rect 2042 18320 2098 18329
rect 1952 18284 2004 18290
rect 2042 18255 2098 18264
rect 1952 18226 2004 18232
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1858 17640 1914 17649
rect 1858 17575 1914 17584
rect 1596 16546 1716 16574
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15881 1348 15982
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15473 1348 15506
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1306 15056 1362 15065
rect 1306 14991 1362 15000
rect 1320 14958 1348 14991
rect 1308 14952 1360 14958
rect 1308 14894 1360 14900
rect 1492 14884 1544 14890
rect 1492 14826 1544 14832
rect 1306 14648 1362 14657
rect 1306 14583 1362 14592
rect 1320 14482 1348 14583
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 1124 10192 1176 10198
rect 1124 10134 1176 10140
rect 940 10124 992 10130
rect 940 10066 992 10072
rect 940 8968 992 8974
rect 940 8910 992 8916
rect 1398 8936 1454 8945
rect 952 8537 980 8910
rect 1398 8871 1454 8880
rect 938 8528 994 8537
rect 938 8463 994 8472
rect 1306 8120 1362 8129
rect 1306 8055 1362 8064
rect 1320 7954 1348 8055
rect 1308 7948 1360 7954
rect 1308 7890 1360 7896
rect 1412 7410 1440 8871
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1504 6914 1532 14826
rect 1582 13424 1638 13433
rect 1582 13359 1638 13368
rect 1596 12306 1624 13359
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1596 9586 1624 9687
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1688 8362 1716 16546
rect 1872 15026 1900 17575
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1858 14512 1914 14521
rect 1858 14447 1914 14456
rect 1766 12880 1822 12889
rect 1766 12815 1768 12824
rect 1820 12815 1822 12824
rect 1768 12786 1820 12792
rect 1766 12608 1822 12617
rect 1766 12543 1822 12552
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1780 7886 1808 12543
rect 1872 9042 1900 14447
rect 1964 11762 1992 17818
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 2056 10674 2084 12038
rect 2148 11762 2176 21558
rect 2240 18358 2268 26200
rect 2412 24200 2464 24206
rect 2412 24142 2464 24148
rect 2320 23588 2372 23594
rect 2320 23530 2372 23536
rect 2332 22030 2360 23530
rect 2320 22024 2372 22030
rect 2320 21966 2372 21972
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 2228 18352 2280 18358
rect 2228 18294 2280 18300
rect 2332 17270 2360 21490
rect 2320 17264 2372 17270
rect 2320 17206 2372 17212
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 2056 8430 2084 10610
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2148 8090 2176 11698
rect 2240 10130 2268 16594
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2332 10674 2360 14894
rect 2424 11762 2452 24142
rect 2884 23254 2912 26200
rect 3330 25664 3386 25673
rect 3330 25599 3386 25608
rect 3344 24886 3372 25599
rect 3422 25256 3478 25265
rect 3422 25191 3478 25200
rect 3332 24880 3384 24886
rect 3332 24822 3384 24828
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 3436 23497 3464 25191
rect 3528 24274 3556 26200
rect 3882 24848 3938 24857
rect 3882 24783 3938 24792
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3792 23792 3844 23798
rect 3792 23734 3844 23740
rect 3422 23488 3478 23497
rect 2950 23420 3258 23429
rect 3422 23423 3478 23432
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2872 23248 2924 23254
rect 2872 23190 2924 23196
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2502 22808 2558 22817
rect 2502 22743 2558 22752
rect 2516 20058 2544 22743
rect 2792 22250 2820 22986
rect 2872 22568 2924 22574
rect 3700 22568 3752 22574
rect 2872 22510 2924 22516
rect 3606 22536 3662 22545
rect 2700 22222 2820 22250
rect 2700 21593 2728 22222
rect 2686 21584 2742 21593
rect 2686 21519 2742 21528
rect 2778 21176 2834 21185
rect 2884 21162 2912 22510
rect 3516 22500 3568 22506
rect 3700 22510 3752 22516
rect 3606 22471 3662 22480
rect 3516 22442 3568 22448
rect 3424 22432 3476 22438
rect 3424 22374 3476 22380
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3436 22273 3464 22374
rect 3422 22264 3478 22273
rect 3422 22199 3478 22208
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2834 21134 2912 21162
rect 2778 21111 2834 21120
rect 2872 20868 2924 20874
rect 2872 20810 2924 20816
rect 2594 20496 2650 20505
rect 2594 20431 2650 20440
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 2504 18692 2556 18698
rect 2504 18634 2556 18640
rect 2516 17921 2544 18634
rect 2502 17912 2558 17921
rect 2502 17847 2558 17856
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2516 11286 2544 15438
rect 2608 11354 2636 20431
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2792 19145 2820 20334
rect 2884 19553 2912 20810
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2870 19544 2926 19553
rect 2870 19479 2926 19488
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3344 18834 3372 21286
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2792 17513 2820 18158
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2870 17776 2926 17785
rect 2870 17711 2926 17720
rect 2778 17504 2834 17513
rect 2778 17439 2834 17448
rect 2884 14414 2912 17711
rect 3344 17202 3372 18566
rect 3436 18290 3464 19246
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3330 16960 3386 16969
rect 2950 16892 3258 16901
rect 3330 16895 3386 16904
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2778 14240 2834 14249
rect 3344 14226 3372 16895
rect 2778 14175 2834 14184
rect 2884 14198 3372 14226
rect 2686 13832 2742 13841
rect 2686 13767 2742 13776
rect 2700 13274 2728 13767
rect 2792 13394 2820 14175
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2700 13246 2820 13274
rect 2792 12918 2820 13246
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2884 12238 2912 14198
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3330 13016 3386 13025
rect 3330 12951 3386 12960
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2872 12232 2924 12238
rect 2778 12200 2834 12209
rect 2872 12174 2924 12180
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2778 12135 2780 12144
rect 2832 12135 2834 12144
rect 2780 12106 2832 12112
rect 2870 12064 2926 12073
rect 2870 11999 2926 12008
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2778 11248 2834 11257
rect 2778 11183 2780 11192
rect 2832 11183 2834 11192
rect 2780 11154 2832 11160
rect 2884 11098 2912 11999
rect 3160 11898 3188 12174
rect 3148 11892 3200 11898
rect 3344 11880 3372 12951
rect 3436 12374 3464 17138
rect 3528 12986 3556 22442
rect 3620 22438 3648 22471
rect 3608 22432 3660 22438
rect 3608 22374 3660 22380
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3620 21729 3648 22170
rect 3606 21720 3662 21729
rect 3606 21655 3662 21664
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3620 14958 3648 21490
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 3712 14090 3740 22510
rect 3804 22234 3832 23734
rect 3896 22982 3924 24783
rect 3974 24032 4030 24041
rect 3974 23967 4030 23976
rect 3884 22976 3936 22982
rect 3884 22918 3936 22924
rect 3792 22228 3844 22234
rect 3792 22170 3844 22176
rect 3790 22128 3846 22137
rect 3790 22063 3846 22072
rect 3804 17134 3832 22063
rect 3988 22012 4016 23967
rect 4068 23792 4120 23798
rect 4172 23780 4200 26200
rect 4804 24200 4856 24206
rect 4802 24168 4804 24177
rect 4856 24168 4858 24177
rect 4802 24103 4858 24112
rect 4712 24064 4764 24070
rect 4712 24006 4764 24012
rect 4120 23752 4200 23780
rect 4068 23734 4120 23740
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 4066 23624 4122 23633
rect 4066 23559 4122 23568
rect 4080 22137 4108 23559
rect 4160 23248 4212 23254
rect 4160 23190 4212 23196
rect 4066 22128 4122 22137
rect 4066 22063 4122 22072
rect 3988 21984 4108 22012
rect 3884 20392 3936 20398
rect 3882 20360 3884 20369
rect 4080 20380 4108 21984
rect 4172 21486 4200 23190
rect 4252 22568 4304 22574
rect 4252 22510 4304 22516
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4160 20800 4212 20806
rect 4158 20768 4160 20777
rect 4212 20768 4214 20777
rect 4158 20703 4214 20712
rect 3936 20360 3938 20369
rect 3882 20295 3938 20304
rect 3988 20352 4108 20380
rect 3882 17368 3938 17377
rect 3882 17303 3938 17312
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3712 14062 3832 14090
rect 3698 13968 3754 13977
rect 3698 13903 3700 13912
rect 3752 13903 3754 13912
rect 3700 13874 3752 13880
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3804 12918 3832 14062
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3344 11852 3648 11880
rect 3148 11834 3200 11840
rect 3422 11792 3478 11801
rect 3422 11727 3478 11736
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2792 11070 2912 11098
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 2792 10062 2820 11070
rect 2870 10568 2926 10577
rect 2870 10503 2926 10512
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2778 9344 2834 9353
rect 2778 9279 2834 9288
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2792 7886 2820 9279
rect 2884 8498 2912 10503
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 3330 10160 3386 10169
rect 3330 10095 3386 10104
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3344 8974 3372 10095
rect 3436 9586 3464 11727
rect 3514 11112 3570 11121
rect 3514 11047 3570 11056
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3528 8498 3556 11047
rect 3620 8634 3648 11852
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 1766 7712 1822 7721
rect 1766 7647 1822 7656
rect 1504 6886 1716 6914
rect 1216 6724 1268 6730
rect 1216 6666 1268 6672
rect 1228 6497 1256 6666
rect 1688 6662 1716 6886
rect 1780 6798 1808 7647
rect 3712 7478 3740 11494
rect 3804 9450 3832 12854
rect 3896 10810 3924 17303
rect 3988 16522 4016 20352
rect 4264 19334 4292 22510
rect 4528 22432 4580 22438
rect 4528 22374 4580 22380
rect 4436 22092 4488 22098
rect 4436 22034 4488 22040
rect 4448 22001 4476 22034
rect 4434 21992 4490 22001
rect 4434 21927 4490 21936
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4172 19306 4292 19334
rect 4172 18222 4200 19306
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4066 17232 4122 17241
rect 4066 17167 4122 17176
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 4080 16402 4108 17167
rect 3988 16374 4108 16402
rect 3988 11150 4016 16374
rect 4172 15881 4200 17614
rect 4158 15872 4214 15881
rect 4158 15807 4214 15816
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 4080 14618 4108 15302
rect 4172 15026 4200 15807
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3792 9444 3844 9450
rect 3792 9386 3844 9392
rect 4080 9178 4108 14350
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 4172 9194 4200 14282
rect 4264 10742 4292 19110
rect 4356 17882 4384 20878
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4342 16552 4398 16561
rect 4342 16487 4398 16496
rect 4356 16182 4384 16487
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 4448 15570 4476 21286
rect 4540 19446 4568 22374
rect 4528 19440 4580 19446
rect 4528 19382 4580 19388
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4434 15328 4490 15337
rect 4434 15263 4490 15272
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4356 12238 4384 14214
rect 4448 12918 4476 15263
rect 4632 14414 4660 23666
rect 4724 18766 4752 24006
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 4804 22976 4856 22982
rect 4908 22953 4936 23666
rect 4986 23216 5042 23225
rect 4986 23151 5042 23160
rect 5000 22982 5028 23151
rect 4988 22976 5040 22982
rect 4804 22918 4856 22924
rect 4894 22944 4950 22953
rect 4816 22094 4844 22918
rect 4988 22918 5040 22924
rect 4894 22879 4950 22888
rect 5092 22574 5120 26302
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26200 7434 27000
rect 8022 26330 8078 27000
rect 7852 26302 8078 26330
rect 5460 23662 5488 26200
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 6104 23186 6132 26200
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 6656 23497 6684 24142
rect 6642 23488 6698 23497
rect 6642 23423 6698 23432
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5356 22500 5408 22506
rect 5356 22442 5408 22448
rect 4816 22066 4936 22094
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 4816 18766 4844 20878
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4804 18760 4856 18766
rect 4908 18737 4936 22066
rect 4988 21072 5040 21078
rect 4988 21014 5040 21020
rect 5000 20874 5028 21014
rect 5172 21004 5224 21010
rect 5172 20946 5224 20952
rect 4988 20868 5040 20874
rect 4988 20810 5040 20816
rect 4804 18702 4856 18708
rect 4894 18728 4950 18737
rect 4816 17678 4844 18702
rect 4894 18663 4950 18672
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4894 16008 4950 16017
rect 4710 15600 4766 15609
rect 4710 15535 4712 15544
rect 4764 15535 4766 15544
rect 4712 15506 4764 15512
rect 4816 15162 4844 15982
rect 4894 15943 4950 15952
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4540 14006 4568 14214
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4540 12918 4568 13194
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4528 12912 4580 12918
rect 4528 12854 4580 12860
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4540 12442 4568 12718
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4434 12336 4490 12345
rect 4434 12271 4490 12280
rect 4448 12238 4476 12271
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4632 11898 4660 14010
rect 4724 12617 4752 15030
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4816 13394 4844 14350
rect 4908 14346 4936 15943
rect 4896 14340 4948 14346
rect 4896 14282 4948 14288
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4710 12608 4766 12617
rect 4710 12543 4766 12552
rect 4724 12306 4752 12543
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4816 12238 4844 13330
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4356 10810 4384 11698
rect 4710 11384 4766 11393
rect 4710 11319 4766 11328
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4724 10742 4752 11319
rect 4816 11218 4844 12174
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4068 9172 4120 9178
rect 4172 9166 4292 9194
rect 4068 9114 4120 9120
rect 4158 9072 4214 9081
rect 4158 9007 4214 9016
rect 4172 8974 4200 9007
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4264 8362 4292 9166
rect 4448 8634 4476 10610
rect 4540 9110 4568 10610
rect 5000 9178 5028 20810
rect 5184 18698 5212 20946
rect 5172 18692 5224 18698
rect 5172 18634 5224 18640
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5092 18086 5120 18362
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 5184 17882 5212 18634
rect 5368 18272 5396 22442
rect 5276 18244 5396 18272
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 5092 15745 5120 17546
rect 5276 17377 5304 18244
rect 5460 18170 5488 23054
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6552 22228 6604 22234
rect 6552 22170 6604 22176
rect 6460 21956 6512 21962
rect 6460 21898 6512 21904
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 5540 21480 5592 21486
rect 5540 21422 5592 21428
rect 5368 18142 5488 18170
rect 5262 17368 5318 17377
rect 5262 17303 5318 17312
rect 5172 17264 5224 17270
rect 5368 17241 5396 18142
rect 5172 17206 5224 17212
rect 5354 17232 5410 17241
rect 5184 16522 5212 17206
rect 5354 17167 5410 17176
rect 5356 17128 5408 17134
rect 5354 17096 5356 17105
rect 5408 17096 5410 17105
rect 5354 17031 5410 17040
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 16658 5304 16934
rect 5354 16688 5410 16697
rect 5264 16652 5316 16658
rect 5354 16623 5410 16632
rect 5264 16594 5316 16600
rect 5172 16516 5224 16522
rect 5172 16458 5224 16464
rect 5078 15736 5134 15745
rect 5078 15671 5134 15680
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5184 13938 5212 15302
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5170 11112 5226 11121
rect 5170 11047 5226 11056
rect 5184 9178 5212 11047
rect 5276 10674 5304 12582
rect 5368 12374 5396 16623
rect 5552 15570 5580 21422
rect 6012 21146 6040 21830
rect 6288 21690 6316 21830
rect 6276 21684 6328 21690
rect 6276 21626 6328 21632
rect 6092 21616 6144 21622
rect 6092 21558 6144 21564
rect 6366 21584 6422 21593
rect 6000 21140 6052 21146
rect 6000 21082 6052 21088
rect 6104 20754 6132 21558
rect 6366 21519 6422 21528
rect 6182 21312 6238 21321
rect 6182 21247 6238 21256
rect 6012 20726 6132 20754
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5816 20392 5868 20398
rect 5816 20334 5868 20340
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5644 19514 5672 20198
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5630 18320 5686 18329
rect 5630 18255 5632 18264
rect 5684 18255 5686 18264
rect 5632 18226 5684 18232
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5552 14482 5580 15506
rect 5644 14482 5672 16934
rect 5736 16114 5764 20334
rect 5828 18873 5856 20334
rect 5920 20058 5948 20334
rect 5908 20052 5960 20058
rect 5908 19994 5960 20000
rect 5814 18864 5870 18873
rect 5814 18799 5870 18808
rect 5828 17864 5856 18799
rect 5828 17836 5948 17864
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5828 15434 5856 17682
rect 5920 17134 5948 17836
rect 6012 17270 6040 20726
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 6000 17264 6052 17270
rect 6000 17206 6052 17212
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 6012 16998 6040 17206
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 5816 15428 5868 15434
rect 5816 15370 5868 15376
rect 6012 15094 6040 16458
rect 6104 16250 6132 20538
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5736 12986 5764 13806
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5446 11792 5502 11801
rect 5446 11727 5448 11736
rect 5500 11727 5502 11736
rect 5448 11698 5500 11704
rect 5552 11354 5580 12718
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5644 9586 5672 12786
rect 5828 12714 5856 14826
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5920 13190 5948 13738
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5816 12708 5868 12714
rect 5816 12650 5868 12656
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5736 11626 5764 12106
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5736 11354 5764 11562
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5920 11234 5948 13126
rect 5828 11218 5948 11234
rect 5816 11212 5948 11218
rect 5868 11206 5948 11212
rect 5816 11154 5868 11160
rect 5920 10606 5948 11206
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 6012 9738 6040 14418
rect 6104 12442 6132 15370
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6196 12288 6224 21247
rect 6276 20868 6328 20874
rect 6276 20810 6328 20816
rect 6288 19786 6316 20810
rect 6276 19780 6328 19786
rect 6276 19722 6328 19728
rect 6288 18834 6316 19722
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6288 17678 6316 18770
rect 6380 18290 6408 21519
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 6288 15026 6316 17614
rect 6380 15502 6408 18022
rect 6472 17218 6500 21898
rect 6564 20466 6592 22170
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6552 19712 6604 19718
rect 6552 19654 6604 19660
rect 6564 18834 6592 19654
rect 6656 19417 6684 22374
rect 6748 22166 6776 26200
rect 7392 24274 7420 26200
rect 7472 24336 7524 24342
rect 7472 24278 7524 24284
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6840 23089 6868 24142
rect 7484 23730 7512 24278
rect 7472 23724 7524 23730
rect 7472 23666 7524 23672
rect 7852 23186 7880 26302
rect 8022 26200 8078 26302
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26330 10010 27000
rect 9692 26302 10010 26330
rect 8576 24880 8628 24886
rect 8576 24822 8628 24828
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8114 23760 8170 23769
rect 8114 23695 8116 23704
rect 8168 23695 8170 23704
rect 8116 23666 8168 23672
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 8220 23174 8432 23202
rect 7288 23112 7340 23118
rect 6826 23080 6882 23089
rect 7288 23054 7340 23060
rect 6826 23015 6882 23024
rect 6920 22704 6972 22710
rect 6920 22646 6972 22652
rect 6828 22432 6880 22438
rect 6828 22374 6880 22380
rect 6840 22234 6868 22374
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6736 22160 6788 22166
rect 6736 22102 6788 22108
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6748 20058 6776 21558
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 6840 21457 6868 21490
rect 6826 21448 6882 21457
rect 6826 21383 6882 21392
rect 6828 21072 6880 21078
rect 6828 21014 6880 21020
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6642 19408 6698 19417
rect 6748 19378 6776 19654
rect 6840 19514 6868 21014
rect 6932 20641 6960 22646
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 7024 22234 7052 22578
rect 7012 22228 7064 22234
rect 7012 22170 7064 22176
rect 7012 22024 7064 22030
rect 7010 21992 7012 22001
rect 7064 21992 7066 22001
rect 7010 21927 7066 21936
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7116 21350 7144 21422
rect 7104 21344 7156 21350
rect 7024 21304 7104 21332
rect 6918 20632 6974 20641
rect 6918 20567 6974 20576
rect 6920 20528 6972 20534
rect 6918 20496 6920 20505
rect 6972 20496 6974 20505
rect 6918 20431 6974 20440
rect 7024 19922 7052 21304
rect 7104 21286 7156 21292
rect 7196 20800 7248 20806
rect 7300 20777 7328 23054
rect 8220 22982 8248 23174
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7392 21622 7420 22510
rect 7380 21616 7432 21622
rect 7380 21558 7432 21564
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7472 20868 7524 20874
rect 7472 20810 7524 20816
rect 7380 20800 7432 20806
rect 7196 20742 7248 20748
rect 7286 20768 7342 20777
rect 7208 20482 7236 20742
rect 7380 20742 7432 20748
rect 7286 20703 7342 20712
rect 7208 20454 7328 20482
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 6642 19343 6698 19352
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6932 17882 6960 19382
rect 7024 19378 7052 19858
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 7010 18728 7066 18737
rect 7010 18663 7066 18672
rect 7024 18222 7052 18663
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6472 17190 6868 17218
rect 6460 17060 6512 17066
rect 6460 17002 6512 17008
rect 6472 16454 6500 17002
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6368 15496 6420 15502
rect 6368 15438 6420 15444
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6288 14346 6316 14962
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 6288 13258 6316 14282
rect 6380 14074 6408 15302
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6276 13252 6328 13258
rect 6276 13194 6328 13200
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 5920 9710 6040 9738
rect 6104 12260 6224 12288
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5920 9518 5948 9710
rect 6104 9654 6132 12260
rect 6288 9654 6316 12718
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6092 9648 6144 9654
rect 5998 9616 6054 9625
rect 6092 9590 6144 9596
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6380 9602 6408 12378
rect 6472 10062 6500 16050
rect 6564 16046 6592 16526
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6564 14482 6592 15846
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6642 15464 6698 15473
rect 6642 15399 6644 15408
rect 6696 15399 6698 15408
rect 6644 15370 6696 15376
rect 6748 15026 6776 15506
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6656 14550 6684 14962
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6734 13696 6790 13705
rect 6734 13631 6790 13640
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6656 12170 6684 13194
rect 6748 12850 6776 13631
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6656 11558 6684 12106
rect 6644 11552 6696 11558
rect 6564 11512 6644 11540
rect 6564 11082 6592 11512
rect 6644 11494 6696 11500
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6380 9574 6500 9602
rect 5998 9551 6054 9560
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 5000 9042 5028 9114
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 6012 8498 6040 9551
rect 6366 9480 6422 9489
rect 6366 9415 6422 9424
rect 6380 8974 6408 9415
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6472 8838 6500 9574
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 3700 7472 3752 7478
rect 3700 7414 3752 7420
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2792 6905 2820 7346
rect 2870 7304 2926 7313
rect 2870 7239 2926 7248
rect 2778 6896 2834 6905
rect 2778 6831 2834 6840
rect 2884 6798 2912 7239
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 6656 6730 6684 11222
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6748 9926 6776 10406
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6748 8838 6776 9454
rect 6840 9178 6868 17190
rect 6932 15042 6960 17614
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 7024 17218 7052 17546
rect 7116 17338 7144 20334
rect 7196 20324 7248 20330
rect 7196 20266 7248 20272
rect 7208 17338 7236 20266
rect 7300 19174 7328 20454
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7300 17338 7328 18566
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7024 17190 7144 17218
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 15706 7052 16390
rect 7116 16153 7144 17190
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7208 16658 7236 17070
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 7392 16522 7420 20742
rect 7484 20398 7512 20810
rect 7472 20392 7524 20398
rect 7472 20334 7524 20340
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7484 19786 7512 19858
rect 7472 19780 7524 19786
rect 7472 19722 7524 19728
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 7102 16144 7158 16153
rect 7102 16079 7158 16088
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 7024 15144 7052 15506
rect 7116 15473 7144 16079
rect 7378 15600 7434 15609
rect 7378 15535 7380 15544
rect 7432 15535 7434 15544
rect 7380 15506 7432 15512
rect 7196 15496 7248 15502
rect 7102 15464 7158 15473
rect 7196 15438 7248 15444
rect 7102 15399 7158 15408
rect 7024 15116 7144 15144
rect 6932 15014 7052 15042
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6932 11898 6960 12106
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6932 10810 6960 11698
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6932 9722 6960 10474
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 7024 9586 7052 15014
rect 7116 14890 7144 15116
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7116 13258 7144 13806
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7208 12102 7236 15438
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 14074 7328 14758
rect 7392 14414 7420 15506
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7208 11762 7236 12038
rect 7300 11830 7328 13738
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12986 7420 13126
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7484 12442 7512 18022
rect 7576 16250 7604 20878
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7668 17134 7696 19246
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7760 16250 7788 17546
rect 7852 17338 7880 22578
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8404 21010 8432 23174
rect 8484 23112 8536 23118
rect 8484 23054 8536 23060
rect 8496 21350 8524 23054
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8392 21004 8444 21010
rect 8392 20946 8444 20952
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8392 20460 8444 20466
rect 8496 20448 8524 21286
rect 8444 20420 8524 20448
rect 8392 20402 8444 20408
rect 8404 19990 8432 20402
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8496 19394 8524 19858
rect 8588 19446 8616 24822
rect 8680 22574 8708 26200
rect 9128 24676 9180 24682
rect 9128 24618 9180 24624
rect 9140 24410 9168 24618
rect 9128 24404 9180 24410
rect 9128 24346 9180 24352
rect 9324 24342 9352 26200
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 9312 24336 9364 24342
rect 9312 24278 9364 24284
rect 9600 24206 9628 24686
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9692 23798 9720 26302
rect 9954 26200 10010 26302
rect 10598 26330 10654 27000
rect 10598 26302 10732 26330
rect 10598 26200 10654 26302
rect 9956 25152 10008 25158
rect 9956 25094 10008 25100
rect 9968 24206 9996 25094
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 10048 24132 10100 24138
rect 10048 24074 10100 24080
rect 9680 23792 9732 23798
rect 9680 23734 9732 23740
rect 10060 23730 10088 24074
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 9956 23724 10008 23730
rect 9956 23666 10008 23672
rect 10048 23724 10100 23730
rect 10048 23666 10100 23672
rect 9968 23633 9996 23666
rect 9954 23624 10010 23633
rect 9954 23559 10010 23568
rect 9036 23248 9088 23254
rect 9036 23190 9088 23196
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8760 20936 8812 20942
rect 8760 20878 8812 20884
rect 8772 19514 8800 20878
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8404 19378 8524 19394
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8392 19372 8524 19378
rect 8444 19366 8524 19372
rect 8668 19372 8720 19378
rect 8392 19314 8444 19320
rect 8668 19314 8720 19320
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 8298 18864 8354 18873
rect 8298 18799 8300 18808
rect 8352 18799 8354 18808
rect 8300 18770 8352 18776
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8496 18329 8524 19178
rect 8576 18692 8628 18698
rect 8576 18634 8628 18640
rect 8482 18320 8538 18329
rect 8024 18284 8076 18290
rect 8482 18255 8538 18264
rect 8024 18226 8076 18232
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 7944 17542 7972 17682
rect 8036 17649 8064 18226
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8022 17640 8078 17649
rect 8022 17575 8078 17584
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8128 16522 8156 16730
rect 8208 16584 8260 16590
rect 8206 16552 8208 16561
rect 8260 16552 8262 16561
rect 8116 16516 8168 16522
rect 8206 16487 8262 16496
rect 8116 16458 8168 16464
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7562 15600 7618 15609
rect 7562 15535 7618 15544
rect 7576 14890 7604 15535
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7576 13870 7604 14350
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7576 12986 7604 13670
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7668 12866 7696 16050
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7760 15473 7788 15982
rect 7746 15464 7802 15473
rect 7746 15399 7802 15408
rect 7852 15094 7880 16390
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7944 16114 7972 16186
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7944 15706 7972 15914
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 8036 15570 8064 15982
rect 8206 15736 8262 15745
rect 8206 15671 8262 15680
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8220 15366 8248 15671
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7840 15088 7892 15094
rect 7746 15056 7802 15065
rect 7840 15030 7892 15036
rect 7746 14991 7802 15000
rect 7760 14958 7788 14991
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7944 14822 7972 14894
rect 7932 14816 7984 14822
rect 7576 12838 7696 12866
rect 7760 14776 7932 14804
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7392 11898 7420 12378
rect 7470 12336 7526 12345
rect 7470 12271 7526 12280
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7288 11688 7340 11694
rect 7286 11656 7288 11665
rect 7380 11688 7432 11694
rect 7340 11656 7342 11665
rect 7196 11620 7248 11626
rect 7380 11630 7432 11636
rect 7286 11591 7342 11600
rect 7196 11562 7248 11568
rect 7102 11112 7158 11121
rect 7102 11047 7158 11056
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 7116 9042 7144 11047
rect 7208 10810 7236 11562
rect 7392 11558 7420 11630
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7300 10146 7328 10950
rect 7392 10606 7420 11494
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7208 10118 7328 10146
rect 7208 9994 7236 10118
rect 7392 10010 7420 10406
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7300 9982 7420 10010
rect 7194 9888 7250 9897
rect 7194 9823 7250 9832
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1214 6488 1270 6497
rect 1214 6423 1270 6432
rect 940 6248 992 6254
rect 940 6190 992 6196
rect 952 6089 980 6190
rect 938 6080 994 6089
rect 938 6015 994 6024
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 940 5704 992 5710
rect 938 5672 940 5681
rect 992 5672 994 5681
rect 938 5607 994 5616
rect 938 5264 994 5273
rect 938 5199 940 5208
rect 992 5199 994 5208
rect 940 5170 992 5176
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 938 4856 994 4865
rect 2950 4859 3258 4868
rect 938 4791 994 4800
rect 952 4690 980 4791
rect 940 4684 992 4690
rect 940 4626 992 4632
rect 1766 4448 1822 4457
rect 1766 4383 1822 4392
rect 1308 4140 1360 4146
rect 1308 4082 1360 4088
rect 940 4072 992 4078
rect 1320 4049 1348 4082
rect 940 4014 992 4020
rect 1306 4040 1362 4049
rect 952 3641 980 4014
rect 1306 3975 1362 3984
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 1780 3534 1808 4383
rect 6748 3942 6776 8774
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 2792 3738 2820 3878
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 1216 3460 1268 3466
rect 1216 3402 1268 3408
rect 1228 3233 1256 3402
rect 1214 3224 1270 3233
rect 1214 3159 1270 3168
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 940 2984 992 2990
rect 940 2926 992 2932
rect 952 2825 980 2926
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 940 2440 992 2446
rect 938 2408 940 2417
rect 1768 2440 1820 2446
rect 992 2408 994 2417
rect 1768 2382 1820 2388
rect 938 2343 994 2352
rect 1412 870 1532 898
rect 1412 800 1440 870
rect 1398 0 1454 800
rect 1504 762 1532 870
rect 1780 762 1808 2382
rect 2792 2009 2820 2994
rect 2778 2000 2834 2009
rect 2778 1935 2834 1944
rect 2884 1601 2912 3470
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 3194 3004 3334
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 7208 3126 7236 9823
rect 7300 6662 7328 9982
rect 7484 9058 7512 12271
rect 7576 10826 7604 12838
rect 7760 12594 7788 14776
rect 7932 14758 7984 14764
rect 8312 14770 8340 17138
rect 8404 16114 8432 18158
rect 8484 17264 8536 17270
rect 8482 17232 8484 17241
rect 8536 17232 8538 17241
rect 8482 17167 8538 17176
rect 8588 17134 8616 18634
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8484 16516 8536 16522
rect 8484 16458 8536 16464
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8404 15881 8432 16050
rect 8390 15872 8446 15881
rect 8390 15807 8446 15816
rect 8312 14742 8432 14770
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7668 12566 7788 12594
rect 7668 12306 7696 12566
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7760 11354 7788 12378
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7852 11218 7880 14214
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8220 13462 8248 13738
rect 8300 13728 8352 13734
rect 8298 13696 8300 13705
rect 8352 13696 8354 13705
rect 8298 13631 8354 13640
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8312 12986 8340 13330
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8404 12434 8432 14742
rect 8496 14414 8524 16458
rect 8588 15434 8616 16934
rect 8680 16182 8708 19314
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8772 17218 8800 18770
rect 8864 17610 8892 19654
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8772 17190 8892 17218
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8668 15632 8720 15638
rect 8668 15574 8720 15580
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8496 13002 8524 13806
rect 8588 13190 8616 15098
rect 8680 14074 8708 15574
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8772 13546 8800 17070
rect 8864 16182 8892 17190
rect 8852 16176 8904 16182
rect 8852 16118 8904 16124
rect 8864 15570 8892 16118
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8680 13518 8800 13546
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8496 12974 8616 13002
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8496 12646 8524 12854
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8312 12406 8432 12434
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7746 11112 7802 11121
rect 7944 11098 7972 11834
rect 7746 11047 7802 11056
rect 7852 11070 7972 11098
rect 7576 10798 7696 10826
rect 7562 10704 7618 10713
rect 7562 10639 7618 10648
rect 7392 9030 7512 9058
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7392 5234 7420 9030
rect 7472 8968 7524 8974
rect 7470 8936 7472 8945
rect 7524 8936 7526 8945
rect 7470 8871 7526 8880
rect 7576 8566 7604 10639
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7668 7274 7696 10798
rect 7760 8498 7788 11047
rect 7852 10690 7880 11070
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7852 10662 7972 10690
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7944 10418 7972 10662
rect 8024 10464 8076 10470
rect 7944 10412 8024 10418
rect 7944 10406 8076 10412
rect 7852 10130 7880 10406
rect 7944 10390 8064 10406
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7852 9518 7880 10066
rect 7944 10033 7972 10390
rect 7930 10024 7986 10033
rect 7930 9959 7986 9968
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7852 3058 7880 9454
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 8312 7818 8340 12406
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 11150 8432 12174
rect 8496 11898 8524 12582
rect 8588 12306 8616 12974
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8404 9654 8432 9930
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8404 7546 8432 9046
rect 8496 7954 8524 9862
rect 8680 8090 8708 13518
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8772 11762 8800 12854
rect 8864 12238 8892 15098
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8772 10674 8800 11698
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8772 10062 8800 10610
rect 8850 10568 8906 10577
rect 8850 10503 8906 10512
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8864 8906 8892 10503
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8956 8498 8984 21830
rect 9048 15502 9076 23190
rect 9496 23044 9548 23050
rect 9496 22986 9548 22992
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9312 21548 9364 21554
rect 9312 21490 9364 21496
rect 9324 21350 9352 21490
rect 9312 21344 9364 21350
rect 9310 21312 9312 21321
rect 9364 21312 9366 21321
rect 9310 21247 9366 21256
rect 9416 20942 9444 21830
rect 9508 21418 9536 22986
rect 9954 22672 10010 22681
rect 9954 22607 9956 22616
rect 10008 22607 10010 22616
rect 9956 22578 10008 22584
rect 9588 21616 9640 21622
rect 9640 21564 9720 21570
rect 9588 21558 9720 21564
rect 9600 21542 9720 21558
rect 9496 21412 9548 21418
rect 9496 21354 9548 21360
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9692 20466 9720 21542
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 9968 21350 9996 21422
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9220 19984 9272 19990
rect 9220 19926 9272 19932
rect 9232 19334 9260 19926
rect 9692 19922 9720 20402
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9312 19780 9364 19786
rect 9312 19722 9364 19728
rect 9324 19689 9352 19722
rect 9404 19712 9456 19718
rect 9310 19680 9366 19689
rect 9404 19654 9456 19660
rect 9310 19615 9366 19624
rect 9232 19306 9352 19334
rect 9128 18352 9180 18358
rect 9128 18294 9180 18300
rect 9140 17678 9168 18294
rect 9324 17746 9352 19306
rect 9416 19281 9444 19654
rect 9402 19272 9458 19281
rect 9402 19207 9458 19216
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9508 18086 9536 18226
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9312 17740 9364 17746
rect 9312 17682 9364 17688
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 9034 15192 9090 15201
rect 9034 15127 9090 15136
rect 9048 14414 9076 15127
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9140 12646 9168 17614
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9232 15337 9260 15370
rect 9218 15328 9274 15337
rect 9218 15263 9274 15272
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9140 12238 9168 12582
rect 9232 12481 9260 15263
rect 9324 15094 9352 16934
rect 9416 16454 9444 17138
rect 9508 17134 9536 17274
rect 9600 17134 9628 18090
rect 9692 17626 9720 18566
rect 9784 17814 9812 19790
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9692 17598 9812 17626
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9402 15600 9458 15609
rect 9402 15535 9458 15544
rect 9416 15162 9444 15535
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 9508 14958 9536 15642
rect 9600 15201 9628 17070
rect 9692 15314 9720 17478
rect 9784 16697 9812 17598
rect 9876 16969 9904 21286
rect 10060 20262 10088 21422
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 10060 20058 10088 20198
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9968 17746 9996 19450
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 10046 17368 10102 17377
rect 10046 17303 10102 17312
rect 10060 17270 10088 17303
rect 10048 17264 10100 17270
rect 10048 17206 10100 17212
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9862 16960 9918 16969
rect 9862 16895 9918 16904
rect 9770 16688 9826 16697
rect 9770 16623 9826 16632
rect 9784 16590 9812 16623
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9692 15286 9904 15314
rect 9586 15192 9642 15201
rect 9586 15127 9642 15136
rect 9770 15192 9826 15201
rect 9770 15127 9826 15136
rect 9586 15056 9642 15065
rect 9784 15042 9812 15127
rect 9642 15014 9812 15042
rect 9586 14991 9642 15000
rect 9496 14952 9548 14958
rect 9772 14952 9824 14958
rect 9692 14912 9772 14940
rect 9692 14906 9720 14912
rect 9496 14894 9548 14900
rect 9646 14878 9720 14906
rect 9772 14894 9824 14900
rect 9646 14498 9674 14878
rect 9876 14550 9904 15286
rect 9496 14476 9548 14482
rect 9600 14470 9674 14498
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9600 14464 9628 14470
rect 9548 14436 9628 14464
rect 9496 14418 9548 14424
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9324 12986 9352 13806
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9218 12472 9274 12481
rect 9218 12407 9274 12416
rect 9324 12306 9352 12922
rect 9416 12617 9444 14350
rect 9600 13870 9628 14436
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9784 14113 9812 14350
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9770 14104 9826 14113
rect 9770 14039 9826 14048
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9402 12608 9458 12617
rect 9402 12543 9458 12552
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9048 9654 9076 9998
rect 9036 9648 9088 9654
rect 9036 9590 9088 9596
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 9048 3126 9076 9590
rect 9126 9480 9182 9489
rect 9126 9415 9182 9424
rect 9140 9042 9168 9415
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9232 8430 9260 11086
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9232 4078 9260 8366
rect 9324 7410 9352 11222
rect 9416 10742 9444 12543
rect 9600 11234 9628 13806
rect 9770 13424 9826 13433
rect 9770 13359 9826 13368
rect 9784 13326 9812 13359
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9876 12850 9904 14214
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12170 9720 12582
rect 9876 12434 9904 12786
rect 9784 12406 9904 12434
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 11830 9720 12106
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9508 11218 9720 11234
rect 9508 11212 9732 11218
rect 9508 11206 9680 11212
rect 9404 10736 9456 10742
rect 9404 10678 9456 10684
rect 9508 9994 9536 11206
rect 9680 11154 9732 11160
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9402 9616 9458 9625
rect 9402 9551 9458 9560
rect 9416 9042 9444 9551
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9600 8090 9628 10610
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9692 9926 9720 10474
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 9042 9720 9862
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9784 7562 9812 12406
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9876 9722 9904 11494
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9876 9110 9904 9522
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9692 7534 9812 7562
rect 9876 7546 9904 8774
rect 9968 8498 9996 17138
rect 10152 16590 10180 24006
rect 10704 22710 10732 26302
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26330 12586 27000
rect 12452 26302 12586 26330
rect 10876 25424 10928 25430
rect 10876 25366 10928 25372
rect 10784 23044 10836 23050
rect 10784 22986 10836 22992
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10796 22506 10824 22986
rect 10508 22500 10560 22506
rect 10508 22442 10560 22448
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 10324 22228 10376 22234
rect 10324 22170 10376 22176
rect 10232 20528 10284 20534
rect 10232 20470 10284 20476
rect 10244 17610 10272 20470
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10336 17202 10364 22170
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10428 20262 10456 20538
rect 10520 20466 10548 22442
rect 10598 22128 10654 22137
rect 10598 22063 10600 22072
rect 10652 22063 10654 22072
rect 10600 22034 10652 22040
rect 10784 21480 10836 21486
rect 10888 21457 10916 25366
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 10968 23112 11020 23118
rect 10968 23054 11020 23060
rect 10980 22982 11008 23054
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 10980 22166 11008 22918
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10784 21422 10836 21428
rect 10874 21448 10930 21457
rect 10796 21350 10824 21422
rect 10874 21383 10930 21392
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10796 21049 10824 21286
rect 10782 21040 10838 21049
rect 10782 20975 10838 20984
rect 10888 20777 10916 21383
rect 10874 20768 10930 20777
rect 10874 20703 10930 20712
rect 11072 20466 11100 25230
rect 11150 24848 11206 24857
rect 11150 24783 11206 24792
rect 11164 22030 11192 24783
rect 11256 22030 11284 26200
rect 11428 25016 11480 25022
rect 11428 24958 11480 24964
rect 11334 24712 11390 24721
rect 11334 24647 11390 24656
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11348 20874 11376 24647
rect 11336 20868 11388 20874
rect 11336 20810 11388 20816
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 10874 18728 10930 18737
rect 10414 18592 10470 18601
rect 10414 18527 10470 18536
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10244 16522 10272 16662
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 10060 14249 10088 16118
rect 10152 16028 10180 16390
rect 10232 16040 10284 16046
rect 10152 16000 10232 16028
rect 10152 14482 10180 16000
rect 10232 15982 10284 15988
rect 10232 15632 10284 15638
rect 10230 15600 10232 15609
rect 10284 15600 10286 15609
rect 10230 15535 10286 15544
rect 10232 15496 10284 15502
rect 10230 15464 10232 15473
rect 10284 15464 10286 15473
rect 10230 15399 10286 15408
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 10140 14272 10192 14278
rect 10046 14240 10102 14249
rect 10140 14214 10192 14220
rect 10046 14175 10102 14184
rect 10060 14006 10088 14175
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 10152 11558 10180 14214
rect 10244 12918 10272 15399
rect 10336 14657 10364 16662
rect 10428 16046 10456 18527
rect 10520 18465 10548 18702
rect 10874 18663 10930 18672
rect 10888 18630 10916 18663
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10506 18456 10562 18465
rect 10968 18420 11020 18426
rect 10506 18391 10562 18400
rect 10520 16454 10548 18391
rect 10888 18380 10968 18408
rect 10888 17134 10916 18380
rect 10968 18362 11020 18368
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10598 16688 10654 16697
rect 10598 16623 10654 16632
rect 10612 16590 10640 16623
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10520 15978 10548 16390
rect 10508 15972 10560 15978
rect 10508 15914 10560 15920
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10416 14884 10468 14890
rect 10416 14826 10468 14832
rect 10322 14648 10378 14657
rect 10322 14583 10378 14592
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10336 14113 10364 14418
rect 10322 14104 10378 14113
rect 10322 14039 10378 14048
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10428 12374 10456 14826
rect 10508 14544 10560 14550
rect 10508 14486 10560 14492
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 10060 7546 10088 9862
rect 10152 9382 10180 10950
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 9864 7540 9916 7546
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 4080 800 4108 2450
rect 6748 800 6776 2450
rect 8036 2310 8064 2926
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8312 2446 8340 2790
rect 9692 2650 9720 7534
rect 9864 7482 9916 7488
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10152 7342 10180 9318
rect 10244 8974 10272 11290
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10336 9722 10364 10542
rect 10520 10130 10548 14486
rect 10612 13734 10640 15846
rect 10704 15706 10732 16934
rect 10888 16726 10916 17070
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 10980 16658 11008 17070
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10796 15434 10824 15642
rect 10876 15632 10928 15638
rect 10876 15574 10928 15580
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10782 15192 10838 15201
rect 10782 15127 10838 15136
rect 10796 15094 10824 15127
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10888 14414 10916 15574
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10704 13546 10732 14214
rect 10612 13518 10732 13546
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10336 8906 10364 9318
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10244 7886 10272 8230
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10336 4010 10364 7686
rect 10612 5710 10640 13518
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12442 10732 13126
rect 10980 12986 11008 15438
rect 11072 15348 11100 20402
rect 11164 16640 11192 20742
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11256 19174 11284 19654
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11256 18834 11284 19110
rect 11244 18828 11296 18834
rect 11244 18770 11296 18776
rect 11348 17338 11376 20810
rect 11440 19689 11468 24958
rect 11796 24336 11848 24342
rect 11796 24278 11848 24284
rect 11808 24206 11836 24278
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 11900 22710 11928 26200
rect 12256 25356 12308 25362
rect 12256 25298 12308 25304
rect 12164 25220 12216 25226
rect 12164 25162 12216 25168
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 11992 22817 12020 24142
rect 11978 22808 12034 22817
rect 11978 22743 12034 22752
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11888 21956 11940 21962
rect 11888 21898 11940 21904
rect 11900 21690 11928 21898
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11900 20505 11928 20538
rect 11886 20496 11942 20505
rect 11612 20460 11664 20466
rect 11886 20431 11942 20440
rect 11612 20402 11664 20408
rect 11520 19712 11572 19718
rect 11426 19680 11482 19689
rect 11520 19654 11572 19660
rect 11426 19615 11482 19624
rect 11428 19236 11480 19242
rect 11428 19178 11480 19184
rect 11440 18816 11468 19178
rect 11532 18970 11560 19654
rect 11520 18964 11572 18970
rect 11520 18906 11572 18912
rect 11520 18828 11572 18834
rect 11440 18788 11520 18816
rect 11520 18770 11572 18776
rect 11428 18692 11480 18698
rect 11428 18634 11480 18640
rect 11440 18290 11468 18634
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11624 17377 11652 20402
rect 11704 20392 11756 20398
rect 11704 20334 11756 20340
rect 11716 20058 11744 20334
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 11702 19272 11758 19281
rect 11702 19207 11758 19216
rect 11610 17368 11666 17377
rect 11336 17332 11388 17338
rect 11610 17303 11666 17312
rect 11336 17274 11388 17280
rect 11610 17096 11666 17105
rect 11610 17031 11666 17040
rect 11520 16652 11572 16658
rect 11164 16612 11376 16640
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11164 16114 11192 16458
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11150 15736 11206 15745
rect 11348 15722 11376 16612
rect 11520 16594 11572 16600
rect 11532 15910 11560 16594
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11348 15694 11560 15722
rect 11150 15671 11206 15680
rect 11164 15502 11192 15671
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11152 15496 11204 15502
rect 11440 15473 11468 15506
rect 11152 15438 11204 15444
rect 11426 15464 11482 15473
rect 11336 15428 11388 15434
rect 11256 15388 11336 15416
rect 11072 15320 11192 15348
rect 11058 15192 11114 15201
rect 11058 15127 11114 15136
rect 11072 14550 11100 15127
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10782 12336 10838 12345
rect 10782 12271 10784 12280
rect 10836 12271 10838 12280
rect 10784 12242 10836 12248
rect 10782 11112 10838 11121
rect 11072 11082 11100 14010
rect 11164 14006 11192 15320
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11256 13938 11284 15388
rect 11426 15399 11482 15408
rect 11336 15370 11388 15376
rect 11532 15314 11560 15694
rect 11348 15286 11560 15314
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11164 11762 11192 13670
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 10782 11047 10784 11056
rect 10836 11047 10838 11056
rect 11060 11076 11112 11082
rect 10784 11018 10836 11024
rect 11060 11018 11112 11024
rect 11164 10606 11192 11222
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11256 10130 11284 10610
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 10784 9648 10836 9654
rect 10782 9616 10784 9625
rect 10836 9616 10838 9625
rect 11256 9586 11284 10066
rect 10782 9551 10838 9560
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11348 8566 11376 15286
rect 11520 15088 11572 15094
rect 11518 15056 11520 15065
rect 11572 15056 11574 15065
rect 11428 15020 11480 15026
rect 11518 14991 11574 15000
rect 11428 14962 11480 14968
rect 11440 14929 11468 14962
rect 11426 14920 11482 14929
rect 11426 14855 11482 14864
rect 11624 14822 11652 17031
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11716 14634 11744 19207
rect 11532 14606 11744 14634
rect 11532 12434 11560 14606
rect 11808 14414 11836 19722
rect 11992 19530 12020 22578
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 11900 19502 12020 19530
rect 11900 18834 11928 19502
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11900 17338 11928 18566
rect 11992 17678 12020 19382
rect 12084 18970 12112 21490
rect 12176 19786 12204 25162
rect 12268 23866 12296 25298
rect 12348 24608 12400 24614
rect 12348 24550 12400 24556
rect 12360 23866 12388 24550
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12452 23798 12480 26302
rect 12530 26200 12586 26302
rect 13174 26330 13230 27000
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12530 24304 12586 24313
rect 12530 24239 12586 24248
rect 12544 24206 12572 24239
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 12440 23792 12492 23798
rect 12440 23734 12492 23740
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12268 21146 12296 22374
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12360 21078 12388 23462
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12806 23216 12862 23225
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12716 23180 12768 23186
rect 12806 23151 12862 23160
rect 12716 23122 12768 23128
rect 12452 22574 12480 23122
rect 12728 23066 12756 23122
rect 12636 23038 12756 23066
rect 12636 22982 12664 23038
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12530 22536 12586 22545
rect 12452 21536 12480 22510
rect 12530 22471 12586 22480
rect 12544 22030 12572 22471
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12532 21548 12584 21554
rect 12452 21508 12532 21536
rect 12348 21072 12400 21078
rect 12348 21014 12400 21020
rect 12254 20496 12310 20505
rect 12254 20431 12256 20440
rect 12308 20431 12310 20440
rect 12256 20402 12308 20408
rect 12452 19990 12480 21508
rect 12532 21490 12584 21496
rect 12636 21010 12664 22646
rect 12820 22250 12848 23151
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 13188 22438 13216 22918
rect 13176 22432 13228 22438
rect 13176 22374 13228 22380
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12728 22222 12848 22250
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12728 20942 12756 22222
rect 13372 22098 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15750 26200 15806 27000
rect 16394 26330 16450 27000
rect 16132 26302 16450 26330
rect 13452 25492 13504 25498
rect 13452 25434 13504 25440
rect 13464 23730 13492 25434
rect 13832 24342 13860 26200
rect 14476 24970 14504 26200
rect 13912 24948 13964 24954
rect 13912 24890 13964 24896
rect 14292 24942 14504 24970
rect 13820 24336 13872 24342
rect 13820 24278 13872 24284
rect 13452 23724 13504 23730
rect 13452 23666 13504 23672
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12820 21350 12848 21626
rect 13464 21486 13492 22374
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12530 20360 12586 20369
rect 12530 20295 12532 20304
rect 12584 20295 12586 20304
rect 12532 20266 12584 20272
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12544 19836 12572 19994
rect 12452 19808 12572 19836
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 12452 18834 12480 19808
rect 12820 19258 12848 21082
rect 13360 20528 13412 20534
rect 13360 20470 13412 20476
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13268 19848 13320 19854
rect 12990 19816 13046 19825
rect 13372 19836 13400 20470
rect 13464 20398 13492 21422
rect 13556 21321 13584 23598
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13832 22642 13860 22986
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13832 21486 13860 22578
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 13820 21344 13872 21350
rect 13542 21312 13598 21321
rect 13820 21286 13872 21292
rect 13542 21247 13598 21256
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13740 19990 13768 20334
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13320 19808 13400 19836
rect 13268 19790 13320 19796
rect 12990 19751 13046 19760
rect 13004 19718 13032 19751
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 13372 19446 13400 19808
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 13360 19440 13412 19446
rect 13360 19382 13412 19388
rect 12636 19242 13032 19258
rect 12636 19236 13044 19242
rect 12636 19230 12992 19236
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12084 18426 12112 18566
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12070 18184 12126 18193
rect 12070 18119 12126 18128
rect 12084 18086 12112 18119
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 15162 11928 16390
rect 11992 16114 12020 17614
rect 12070 17368 12126 17377
rect 12070 17303 12126 17312
rect 12084 16590 12112 17303
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 12070 16144 12126 16153
rect 11980 16108 12032 16114
rect 12070 16079 12126 16088
rect 11980 16050 12032 16056
rect 12084 15706 12112 16079
rect 12268 16017 12296 18770
rect 12438 18456 12494 18465
rect 12438 18391 12440 18400
rect 12492 18391 12494 18400
rect 12440 18362 12492 18368
rect 12544 18306 12572 18838
rect 12452 18278 12572 18306
rect 12452 18154 12480 18278
rect 12440 18148 12492 18154
rect 12440 18090 12492 18096
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12346 18048 12402 18057
rect 12346 17983 12402 17992
rect 12360 17882 12388 17983
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12438 17504 12494 17513
rect 12438 17439 12494 17448
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12254 16008 12310 16017
rect 12254 15943 12310 15952
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11978 15056 12034 15065
rect 11978 14991 11980 15000
rect 12032 14991 12034 15000
rect 11980 14962 12032 14968
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11440 12406 11560 12434
rect 11440 9450 11468 12406
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11532 11218 11560 11630
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11532 10130 11560 10746
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11060 8288 11112 8294
rect 10966 8256 11022 8265
rect 11060 8230 11112 8236
rect 10966 8191 11022 8200
rect 10980 7954 11008 8191
rect 11072 8090 11100 8230
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 11164 3738 11192 8298
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11256 3398 11284 8366
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11532 3534 11560 7890
rect 11624 4622 11652 13874
rect 11716 6254 11744 13874
rect 11992 13394 12020 14350
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 12084 13002 12112 15438
rect 12176 13802 12204 15846
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12268 15366 12296 15642
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12360 14958 12388 16730
rect 12452 16658 12480 17439
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12544 15994 12572 18090
rect 12636 18057 12664 19230
rect 12992 19178 13044 19184
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12714 18320 12770 18329
rect 12714 18255 12770 18264
rect 12808 18284 12860 18290
rect 12622 18048 12678 18057
rect 12622 17983 12678 17992
rect 12728 17610 12756 18255
rect 12808 18226 12860 18232
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12636 16182 12664 17002
rect 12728 16250 12756 17546
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 12544 15966 12664 15994
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12268 14278 12296 14554
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12452 13734 12480 15302
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 11992 12974 12112 13002
rect 11992 12442 12020 12974
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11992 11898 12020 12174
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11900 11354 11928 11630
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 11796 8628 11848 8634
rect 11900 8616 11928 11018
rect 11992 11014 12020 11698
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11992 10470 12020 10950
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 12084 8974 12112 12854
rect 12360 12306 12388 13194
rect 12348 12300 12400 12306
rect 12268 12260 12348 12288
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12176 11762 12204 11834
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12176 10810 12204 11562
rect 12268 11354 12296 12260
rect 12348 12242 12400 12248
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12268 10690 12296 11154
rect 12360 10742 12388 11494
rect 12176 10662 12296 10690
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12176 9722 12204 10662
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12268 9042 12296 10066
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 11848 8588 11928 8616
rect 11796 8570 11848 8576
rect 11992 7410 12020 8774
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 12084 3670 12112 8774
rect 12360 8514 12388 9862
rect 12452 8974 12480 12038
rect 12544 11830 12572 13194
rect 12636 12753 12664 15966
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12728 14482 12756 15506
rect 12820 15162 12848 18226
rect 12912 18086 12940 18770
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13188 18086 13216 18702
rect 13372 18329 13400 19382
rect 13556 18834 13584 19722
rect 13740 19446 13768 19926
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13358 18320 13414 18329
rect 13358 18255 13414 18264
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13268 17740 13320 17746
rect 13372 17728 13400 18158
rect 13320 17700 13400 17728
rect 13268 17682 13320 17688
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13280 15892 13308 16390
rect 13372 16250 13400 17700
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13464 16289 13492 16594
rect 13556 16522 13584 18226
rect 13648 17814 13676 19246
rect 13740 18358 13768 19246
rect 13832 18873 13860 21286
rect 13818 18864 13874 18873
rect 13818 18799 13874 18808
rect 13924 18766 13952 24890
rect 14292 24274 14320 24942
rect 14280 24268 14332 24274
rect 14280 24210 14332 24216
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14830 24168 14886 24177
rect 14476 23866 14504 24142
rect 14830 24103 14886 24112
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14476 22234 14504 22714
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 14004 20800 14056 20806
rect 14004 20742 14056 20748
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13820 17876 13872 17882
rect 13740 17836 13820 17864
rect 13636 17808 13688 17814
rect 13740 17785 13768 17836
rect 13820 17818 13872 17824
rect 13636 17750 13688 17756
rect 13726 17776 13782 17785
rect 13648 17134 13676 17750
rect 13726 17711 13782 17720
rect 13726 17640 13782 17649
rect 13726 17575 13782 17584
rect 13740 17542 13768 17575
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13924 17270 13952 18702
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13634 16960 13690 16969
rect 13634 16895 13690 16904
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13450 16280 13506 16289
rect 13360 16244 13412 16250
rect 13450 16215 13506 16224
rect 13360 16186 13412 16192
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13280 15864 13400 15892
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12728 14249 12756 14282
rect 12714 14240 12770 14249
rect 12714 14175 12770 14184
rect 12728 13297 12756 14175
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12714 13288 12770 13297
rect 12714 13223 12716 13232
rect 12768 13223 12770 13232
rect 12716 13194 12768 13200
rect 12820 12850 12848 13874
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12622 12744 12678 12753
rect 12622 12679 12678 12688
rect 12806 12744 12862 12753
rect 12806 12679 12862 12688
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 12102 12664 12582
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12820 11880 12848 12679
rect 13372 12646 13400 15864
rect 13556 14958 13584 15982
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13464 14657 13492 14894
rect 13450 14648 13506 14657
rect 13450 14583 13506 14592
rect 13556 14550 13584 14894
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13464 13530 13492 14418
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13648 13190 13676 16895
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13832 12646 13860 15098
rect 13924 14278 13952 15846
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 12728 11852 12848 11880
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12544 11082 12572 11766
rect 12532 11076 12584 11082
rect 12584 11036 12664 11064
rect 12532 11018 12584 11024
rect 12636 10742 12664 11036
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12636 10062 12664 10678
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12360 8486 12480 8514
rect 12452 8430 12480 8486
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12440 8016 12492 8022
rect 12636 7970 12664 8774
rect 12728 8090 12756 11852
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12820 10266 12848 11698
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12806 10160 12862 10169
rect 12806 10095 12862 10104
rect 12900 10124 12952 10130
rect 12820 8634 12848 10095
rect 13084 10124 13136 10130
rect 12952 10084 13084 10112
rect 12900 10066 12952 10072
rect 13084 10066 13136 10072
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13188 9518 13216 9998
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 13372 8956 13400 12038
rect 13450 10024 13506 10033
rect 13450 9959 13452 9968
rect 13504 9959 13506 9968
rect 13452 9930 13504 9936
rect 13464 9586 13492 9930
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13372 8928 13492 8956
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8634 13124 8842
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 13372 8090 13400 8434
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 12492 7964 12664 7970
rect 12440 7958 12664 7964
rect 12452 7942 12664 7958
rect 13464 7750 13492 8928
rect 13648 8838 13676 9454
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13740 8430 13768 9862
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13832 7410 13860 8978
rect 14016 8294 14044 20742
rect 14108 20398 14136 21286
rect 14292 20534 14320 21422
rect 14384 21049 14412 21898
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14370 21040 14426 21049
rect 14370 20975 14426 20984
rect 14752 20806 14780 21286
rect 14844 21010 14872 24103
rect 15120 22166 15148 26200
rect 15764 23798 15792 26200
rect 15844 25084 15896 25090
rect 15844 25026 15896 25032
rect 15752 23792 15804 23798
rect 15752 23734 15804 23740
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 15212 23186 15240 23666
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 15200 23180 15252 23186
rect 15200 23122 15252 23128
rect 15304 23050 15332 23530
rect 15292 23044 15344 23050
rect 15292 22986 15344 22992
rect 15750 22808 15806 22817
rect 15750 22743 15806 22752
rect 15108 22160 15160 22166
rect 15108 22102 15160 22108
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 14936 21622 14964 21830
rect 14924 21616 14976 21622
rect 14924 21558 14976 21564
rect 15028 21554 15056 21830
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 14108 18902 14136 20334
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14568 19514 14596 19790
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14476 18154 14504 18566
rect 14568 18358 14596 19450
rect 14660 18902 14688 20198
rect 15028 19281 15056 21490
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15212 20806 15240 21422
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15488 20874 15516 21286
rect 15476 20868 15528 20874
rect 15476 20810 15528 20816
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15292 20460 15344 20466
rect 15120 20420 15292 20448
rect 15120 20262 15148 20420
rect 15292 20402 15344 20408
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 15304 19786 15332 20266
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15396 19802 15424 19994
rect 15488 19922 15516 20198
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15292 19780 15344 19786
rect 15396 19774 15516 19802
rect 15292 19722 15344 19728
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15014 19272 15070 19281
rect 15014 19207 15070 19216
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 14648 18896 14700 18902
rect 14648 18838 14700 18844
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 14556 18352 14608 18358
rect 14556 18294 14608 18300
rect 14464 18148 14516 18154
rect 14464 18090 14516 18096
rect 15028 17513 15056 18634
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 15120 18329 15148 18362
rect 15106 18320 15162 18329
rect 15106 18255 15162 18264
rect 15304 17649 15332 19110
rect 15290 17640 15346 17649
rect 15396 17610 15424 19382
rect 15488 18698 15516 19774
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15488 18465 15516 18634
rect 15580 18630 15608 20198
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15474 18456 15530 18465
rect 15474 18391 15530 18400
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15290 17575 15346 17584
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15014 17504 15070 17513
rect 15014 17439 15070 17448
rect 14094 17096 14150 17105
rect 14094 17031 14150 17040
rect 14924 17060 14976 17066
rect 14108 13462 14136 17031
rect 14924 17002 14976 17008
rect 14188 16992 14240 16998
rect 14186 16960 14188 16969
rect 14832 16992 14884 16998
rect 14240 16960 14242 16969
rect 14832 16934 14884 16940
rect 14186 16895 14242 16904
rect 14186 16824 14242 16833
rect 14186 16759 14242 16768
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 14200 10198 14228 16759
rect 14844 16250 14872 16934
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14936 16130 14964 17002
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15396 16454 15424 16594
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 14844 16102 14964 16130
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14476 13870 14504 15982
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14556 14952 14608 14958
rect 14608 14912 14688 14940
rect 14556 14894 14608 14900
rect 14660 14414 14688 14912
rect 14752 14618 14780 15302
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14462 13696 14518 13705
rect 14462 13631 14518 13640
rect 14476 12782 14504 13631
rect 14660 13394 14688 14350
rect 14844 14074 14872 16102
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14936 14958 14964 15506
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 15028 13530 15056 15982
rect 15106 15736 15162 15745
rect 15106 15671 15162 15680
rect 15120 15450 15148 15671
rect 15120 15434 15240 15450
rect 15120 15428 15252 15434
rect 15120 15422 15200 15428
rect 15200 15370 15252 15376
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 15120 14278 15148 15030
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15304 14618 15332 14894
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 15014 13288 15070 13297
rect 15120 13274 15148 14214
rect 15212 13870 15240 14214
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15070 13246 15148 13274
rect 15014 13223 15016 13232
rect 15068 13223 15070 13232
rect 15016 13194 15068 13200
rect 15212 13190 15240 13806
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14752 11558 14780 12786
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14568 11218 14596 11494
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14188 10192 14240 10198
rect 14188 10134 14240 10140
rect 14292 8362 14320 10610
rect 14568 10130 14596 11154
rect 14556 10124 14608 10130
rect 14476 10084 14556 10112
rect 14476 9586 14504 10084
rect 14556 10066 14608 10072
rect 14752 9994 14780 11290
rect 14844 10130 14872 12242
rect 15028 12170 15056 12854
rect 15304 12374 15332 13942
rect 15396 13938 15424 16186
rect 15488 15638 15516 16390
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14482 15516 14894
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15396 13190 15424 13670
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 15292 12368 15344 12374
rect 15292 12310 15344 12316
rect 15396 12170 15424 12650
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15120 11218 15148 12106
rect 15290 12064 15346 12073
rect 15290 11999 15346 12008
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15304 11082 15332 11999
rect 15488 11200 15516 12582
rect 15580 11898 15608 17614
rect 15672 16833 15700 19314
rect 15764 17762 15792 22743
rect 15856 19446 15884 25026
rect 16132 22710 16160 26302
rect 16394 26200 16450 26302
rect 17038 26200 17094 27000
rect 17682 26330 17738 27000
rect 17420 26302 17738 26330
rect 16212 24132 16264 24138
rect 16212 24074 16264 24080
rect 16224 23322 16252 24074
rect 16212 23316 16264 23322
rect 16212 23258 16264 23264
rect 16948 23112 17000 23118
rect 16578 23080 16634 23089
rect 16948 23054 17000 23060
rect 16578 23015 16634 23024
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 16592 22642 16620 23015
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16672 21956 16724 21962
rect 16672 21898 16724 21904
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16396 20800 16448 20806
rect 16396 20742 16448 20748
rect 16408 20466 16436 20742
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 15936 20324 15988 20330
rect 15936 20266 15988 20272
rect 15844 19440 15896 19446
rect 15844 19382 15896 19388
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15856 18601 15884 19246
rect 15948 19174 15976 20266
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 16120 18828 16172 18834
rect 16316 18816 16344 19246
rect 16172 18788 16344 18816
rect 16120 18770 16172 18776
rect 15842 18592 15898 18601
rect 15842 18527 15898 18536
rect 16118 17912 16174 17921
rect 16118 17847 16174 17856
rect 15764 17734 15976 17762
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15658 16824 15714 16833
rect 15658 16759 15714 16768
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15672 15201 15700 16390
rect 15658 15192 15714 15201
rect 15658 15127 15714 15136
rect 15660 13456 15712 13462
rect 15660 13398 15712 13404
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15672 11694 15700 13398
rect 15764 12442 15792 17614
rect 15948 17610 15976 17734
rect 15936 17604 15988 17610
rect 15936 17546 15988 17552
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15948 16794 15976 16934
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15856 14958 15884 16594
rect 16040 15638 16068 17070
rect 16132 16561 16160 17847
rect 16316 17746 16344 18788
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16118 16552 16174 16561
rect 16118 16487 16174 16496
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16132 15706 16160 15846
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16028 15632 16080 15638
rect 16028 15574 16080 15580
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16132 14482 16160 14758
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16224 14362 16252 17478
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16316 14929 16344 15302
rect 16302 14920 16358 14929
rect 16302 14855 16358 14864
rect 16132 14334 16252 14362
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15856 12782 15884 13330
rect 16040 12986 16068 13806
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15856 12306 15884 12718
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15948 11880 15976 12718
rect 16132 12434 16160 14334
rect 16408 14006 16436 20402
rect 16486 18048 16542 18057
rect 16486 17983 16542 17992
rect 16500 15570 16528 17983
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 15764 11852 15976 11880
rect 16040 12406 16160 12434
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15396 11172 15516 11200
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15028 10266 15056 11018
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15212 10470 15240 10950
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14740 9988 14792 9994
rect 14740 9930 14792 9936
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14844 9518 14872 10066
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14752 9042 14780 9318
rect 14936 9042 14964 10066
rect 15304 10033 15332 11018
rect 15290 10024 15346 10033
rect 15290 9959 15292 9968
rect 15344 9959 15346 9968
rect 15292 9930 15344 9936
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 15396 8498 15424 11172
rect 15764 11098 15792 11852
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15580 11070 15792 11098
rect 15580 10810 15608 11070
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15672 10538 15700 10950
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15764 10554 15792 10678
rect 15660 10532 15712 10538
rect 15764 10526 15884 10554
rect 15660 10474 15712 10480
rect 15856 10198 15884 10526
rect 15844 10192 15896 10198
rect 15844 10134 15896 10140
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9416 800 9444 2450
rect 9784 2446 9812 3130
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 11624 2378 11652 3334
rect 12636 3126 12664 5782
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 15212 4146 15240 7958
rect 15488 5778 15516 9046
rect 15948 8838 15976 11698
rect 16040 10470 16068 12406
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16132 11762 16160 12174
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 16224 10169 16252 13874
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16316 12782 16344 13806
rect 16486 13288 16542 13297
rect 16486 13223 16542 13232
rect 16500 13190 16528 13223
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11354 16528 12106
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16592 10713 16620 21490
rect 16684 21010 16712 21898
rect 16672 21004 16724 21010
rect 16672 20946 16724 20952
rect 16960 20913 16988 23054
rect 17052 21486 17080 26200
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17132 24268 17184 24274
rect 17132 24210 17184 24216
rect 17144 23118 17172 24210
rect 17236 24138 17264 24754
rect 17224 24132 17276 24138
rect 17224 24074 17276 24080
rect 17420 23186 17448 26302
rect 17682 26200 17738 26302
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26200 20958 27000
rect 21546 26200 21602 27000
rect 22190 26200 22246 27000
rect 22834 26330 22890 27000
rect 22834 26302 23336 26330
rect 22834 26200 22890 26302
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 17144 22098 17172 23054
rect 17512 23050 17540 24006
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23662 18368 26200
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18512 24132 18564 24138
rect 18512 24074 18564 24080
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 17776 23588 17828 23594
rect 17776 23530 17828 23536
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17224 22568 17276 22574
rect 17224 22510 17276 22516
rect 17132 22092 17184 22098
rect 17132 22034 17184 22040
rect 17236 21894 17264 22510
rect 17406 21992 17462 22001
rect 17406 21927 17462 21936
rect 17500 21956 17552 21962
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 17040 21480 17092 21486
rect 17040 21422 17092 21428
rect 17236 21418 17264 21830
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17314 21312 17370 21321
rect 17314 21247 17370 21256
rect 17040 20936 17092 20942
rect 16946 20904 17002 20913
rect 16856 20868 16908 20874
rect 17040 20878 17092 20884
rect 16946 20839 17002 20848
rect 16856 20810 16908 20816
rect 16868 20754 16896 20810
rect 17052 20754 17080 20878
rect 17132 20868 17184 20874
rect 17132 20810 17184 20816
rect 16868 20726 17080 20754
rect 17144 19922 17172 20810
rect 17328 20602 17356 21247
rect 17420 20942 17448 21927
rect 17500 21898 17552 21904
rect 17512 21350 17540 21898
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17316 20596 17368 20602
rect 17316 20538 17368 20544
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 17132 19440 17184 19446
rect 16854 19408 16910 19417
rect 16764 19372 16816 19378
rect 17132 19382 17184 19388
rect 16854 19343 16910 19352
rect 16764 19314 16816 19320
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16684 18766 16712 19110
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16684 18222 16712 18566
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16684 17746 16712 18158
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16776 16590 16804 19314
rect 16868 19174 16896 19343
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 17144 17746 17172 19382
rect 17236 18902 17264 20538
rect 17420 20466 17448 20742
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17316 20256 17368 20262
rect 17316 20198 17368 20204
rect 17224 18896 17276 18902
rect 17224 18838 17276 18844
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17130 17368 17186 17377
rect 17130 17303 17186 17312
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16868 16794 16896 17138
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 16960 16794 16988 17002
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16684 13326 16712 15846
rect 17052 15502 17080 17002
rect 17144 16998 17172 17303
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16960 15162 16988 15438
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 16946 14376 17002 14385
rect 17052 14346 17080 15438
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 16946 14311 17002 14320
rect 17040 14340 17092 14346
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16578 10704 16634 10713
rect 16578 10639 16634 10648
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16210 10160 16266 10169
rect 16210 10095 16266 10104
rect 16118 10024 16174 10033
rect 16118 9959 16174 9968
rect 16132 9586 16160 9959
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16316 9382 16344 10542
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 8906 16344 9318
rect 16304 8900 16356 8906
rect 16304 8842 16356 8848
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 16684 7818 16712 12242
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16868 11626 16896 12038
rect 16960 11898 16988 14311
rect 17040 14282 17092 14288
rect 17052 13870 17080 14282
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17052 13394 17080 13806
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 17052 12073 17080 12106
rect 17038 12064 17094 12073
rect 17038 11999 17094 12008
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16868 10062 16896 11086
rect 17052 10674 17080 11494
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 17040 10532 17092 10538
rect 17040 10474 17092 10480
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16868 9518 16896 9998
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16868 9042 16896 9454
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15580 5234 15608 7210
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16500 5234 16528 7142
rect 16868 5778 16896 8978
rect 16960 8498 16988 10134
rect 17052 10130 17080 10474
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 12084 800 12112 2450
rect 12544 2446 12572 2858
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 14752 800 14780 2450
rect 15028 2446 15056 3878
rect 15488 3126 15516 5102
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 17052 3058 17080 5510
rect 17144 3466 17172 14962
rect 17236 14346 17264 15302
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 17328 12306 17356 20198
rect 17788 19145 17816 23530
rect 18524 23118 18552 24074
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18524 22710 18552 23054
rect 18512 22704 18564 22710
rect 18512 22646 18564 22652
rect 18524 22438 18552 22646
rect 18616 22574 18644 24754
rect 18788 24676 18840 24682
rect 18788 24618 18840 24624
rect 18800 24206 18828 24618
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18984 23322 19012 26200
rect 19064 24676 19116 24682
rect 19064 24618 19116 24624
rect 19076 23662 19104 24618
rect 19628 24426 19656 26200
rect 19352 24398 19656 24426
rect 19352 23798 19380 24398
rect 19800 24200 19852 24206
rect 19800 24142 19852 24148
rect 19522 23896 19578 23905
rect 19522 23831 19578 23840
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 18972 23316 19024 23322
rect 18972 23258 19024 23264
rect 19076 23254 19104 23598
rect 19536 23322 19564 23831
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19064 23248 19116 23254
rect 19064 23190 19116 23196
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 19064 22432 19116 22438
rect 19064 22374 19116 22380
rect 18524 22030 18552 22374
rect 18880 22160 18932 22166
rect 18880 22102 18932 22108
rect 18696 22092 18748 22098
rect 18696 22034 18748 22040
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18602 21720 18658 21729
rect 18602 21655 18658 21664
rect 18328 21412 18380 21418
rect 18328 21354 18380 21360
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17880 19961 17908 21082
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18340 20584 18368 21354
rect 18616 21010 18644 21655
rect 18708 21486 18736 22034
rect 18788 21956 18840 21962
rect 18788 21898 18840 21904
rect 18800 21690 18828 21898
rect 18788 21684 18840 21690
rect 18788 21626 18840 21632
rect 18696 21480 18748 21486
rect 18696 21422 18748 21428
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18420 20800 18472 20806
rect 18418 20768 18420 20777
rect 18472 20768 18474 20777
rect 18418 20703 18474 20712
rect 18248 20556 18368 20584
rect 17866 19952 17922 19961
rect 18248 19922 18276 20556
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18432 19922 18460 20402
rect 17866 19887 17922 19896
rect 18236 19916 18288 19922
rect 18236 19858 18288 19864
rect 18420 19916 18472 19922
rect 18420 19858 18472 19864
rect 18248 19786 18276 19858
rect 18236 19780 18288 19786
rect 18236 19722 18288 19728
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17774 19136 17830 19145
rect 17774 19071 17830 19080
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17498 18456 17554 18465
rect 17498 18391 17554 18400
rect 17512 18358 17540 18391
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17696 17678 17724 18634
rect 17788 18154 17816 18702
rect 18064 18698 18092 19246
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18156 18970 18184 19110
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18340 18834 18368 19178
rect 18328 18828 18380 18834
rect 18328 18770 18380 18776
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17776 18148 17828 18154
rect 17776 18090 17828 18096
rect 18340 18057 18368 18566
rect 18432 18358 18460 19654
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18326 18048 18382 18057
rect 18326 17983 18382 17992
rect 18432 17882 18460 18158
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17696 17270 17724 17614
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17420 14006 17448 15982
rect 17512 15366 17540 17070
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17880 15978 17908 16526
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 18340 16046 18368 17818
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18432 17542 18460 17682
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18432 17134 18460 17478
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18432 16726 18460 17070
rect 18420 16720 18472 16726
rect 18420 16662 18472 16668
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 18432 15688 18460 16526
rect 18524 16114 18552 20402
rect 18708 19446 18736 21422
rect 18892 20398 18920 22102
rect 19076 22030 19104 22374
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18984 20534 19012 21830
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 19076 21010 19104 21422
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 18604 19304 18656 19310
rect 18602 19272 18604 19281
rect 18656 19272 18658 19281
rect 18602 19207 18658 19216
rect 18602 18864 18658 18873
rect 18602 18799 18658 18808
rect 18616 18465 18644 18799
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18602 18456 18658 18465
rect 18602 18391 18658 18400
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18616 17649 18644 18294
rect 18602 17640 18658 17649
rect 18602 17575 18658 17584
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18340 15660 18460 15688
rect 17684 15428 17736 15434
rect 17604 15388 17684 15416
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17604 14346 17632 15388
rect 17684 15370 17736 15376
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17604 13988 17632 14282
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18340 14074 18368 15660
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18432 14074 18460 15506
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 17684 14000 17736 14006
rect 17604 13960 17684 13988
rect 17420 13530 17448 13942
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17512 12714 17540 13330
rect 17604 13240 17632 13960
rect 17684 13942 17736 13948
rect 17684 13252 17736 13258
rect 17604 13212 17684 13240
rect 17500 12708 17552 12714
rect 17500 12650 17552 12656
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17224 11620 17276 11626
rect 17224 11562 17276 11568
rect 17236 9654 17264 11562
rect 17328 10606 17356 12038
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17420 10810 17448 11630
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17420 9994 17448 10746
rect 17512 10674 17540 12650
rect 17604 12073 17632 13212
rect 17684 13194 17736 13200
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17590 12064 17646 12073
rect 17590 11999 17646 12008
rect 17880 11898 17908 12786
rect 18432 12442 18460 13126
rect 18616 12481 18644 17575
rect 18708 15008 18736 18702
rect 18800 16794 18828 19790
rect 18892 19378 18920 19994
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18972 19304 19024 19310
rect 18970 19272 18972 19281
rect 19024 19272 19026 19281
rect 18970 19207 19026 19216
rect 18970 19136 19026 19145
rect 18970 19071 19026 19080
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18892 17542 18920 18634
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18892 17134 18920 17478
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18892 15042 18920 16730
rect 18984 16114 19012 19071
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 18892 15014 19012 15042
rect 18708 14980 18828 15008
rect 18694 14648 18750 14657
rect 18694 14583 18750 14592
rect 18708 14006 18736 14583
rect 18800 14550 18828 14980
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18602 12472 18658 12481
rect 18420 12436 18472 12442
rect 18602 12407 18658 12416
rect 18420 12378 18472 12384
rect 18708 12356 18736 13942
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18800 13190 18828 13874
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18892 12918 18920 14894
rect 18984 13938 19012 15014
rect 19076 14958 19104 20198
rect 19168 16454 19196 22578
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19352 22166 19380 22374
rect 19522 22264 19578 22273
rect 19522 22199 19524 22208
rect 19576 22199 19578 22208
rect 19524 22170 19576 22176
rect 19340 22160 19392 22166
rect 19340 22102 19392 22108
rect 19628 22094 19656 23598
rect 19708 23520 19760 23526
rect 19708 23462 19760 23468
rect 19720 23186 19748 23462
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 19720 22778 19748 23122
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19628 22066 19748 22094
rect 19294 22024 19346 22030
rect 19616 22024 19668 22030
rect 19346 21984 19616 22012
rect 19294 21966 19346 21972
rect 19616 21966 19668 21972
rect 19340 21888 19392 21894
rect 19338 21856 19340 21865
rect 19392 21856 19394 21865
rect 19338 21791 19394 21800
rect 19720 21690 19748 22066
rect 19708 21684 19760 21690
rect 19708 21626 19760 21632
rect 19524 21140 19576 21146
rect 19576 21100 19656 21128
rect 19524 21082 19576 21088
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19260 18358 19288 20742
rect 19352 19378 19380 20742
rect 19522 20632 19578 20641
rect 19522 20567 19578 20576
rect 19536 19990 19564 20567
rect 19524 19984 19576 19990
rect 19524 19926 19576 19932
rect 19524 19712 19576 19718
rect 19522 19680 19524 19689
rect 19576 19680 19578 19689
rect 19522 19615 19578 19624
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19628 19242 19656 21100
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19720 20466 19748 20946
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19720 19922 19748 20402
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19616 19236 19668 19242
rect 19616 19178 19668 19184
rect 19720 18834 19748 19246
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19248 18352 19300 18358
rect 19248 18294 19300 18300
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19156 16448 19208 16454
rect 19156 16390 19208 16396
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19064 14544 19116 14550
rect 19064 14486 19116 14492
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18984 13258 19012 13670
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18788 12776 18840 12782
rect 18984 12764 19012 13194
rect 18788 12718 18840 12724
rect 18892 12736 19012 12764
rect 18524 12328 18736 12356
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18524 11898 18552 12328
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17604 10266 17632 11630
rect 18800 11354 18828 12718
rect 18892 11354 18920 12736
rect 19076 12594 19104 14486
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19168 13444 19196 14282
rect 19260 14074 19288 17614
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19536 16810 19564 16934
rect 19444 16794 19564 16810
rect 19432 16788 19564 16794
rect 19484 16782 19564 16788
rect 19432 16730 19484 16736
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19352 15502 19380 16458
rect 19444 15570 19472 16526
rect 19522 16008 19578 16017
rect 19522 15943 19578 15952
rect 19536 15706 19564 15943
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19168 13416 19288 13444
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 18984 12566 19104 12594
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17880 10742 17908 11018
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17880 10033 17908 10678
rect 18800 10538 18828 11290
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 17866 10024 17922 10033
rect 17408 9988 17460 9994
rect 17866 9959 17868 9968
rect 17408 9930 17460 9936
rect 17920 9959 17922 9968
rect 18418 10024 18474 10033
rect 18418 9959 18474 9968
rect 17868 9930 17920 9936
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 18432 9654 18460 9959
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 18420 9648 18472 9654
rect 18984 9625 19012 12566
rect 19062 12472 19118 12481
rect 19062 12407 19118 12416
rect 19076 11762 19104 12407
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 19168 11150 19196 12854
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19260 10266 19288 13416
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19352 11014 19380 13262
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19444 10470 19472 14214
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19536 11121 19564 13670
rect 19522 11112 19578 11121
rect 19522 11047 19578 11056
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 18420 9590 18472 9596
rect 18970 9616 19026 9625
rect 17420 9110 17448 9590
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 17408 9104 17460 9110
rect 17408 9046 17460 9052
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18340 8430 18368 9454
rect 18432 8974 18460 9590
rect 18970 9551 19026 9560
rect 19260 9518 19288 10202
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18432 5642 18460 8910
rect 19444 8906 19472 9522
rect 19628 9450 19656 17614
rect 19720 15366 19748 18634
rect 19812 18290 19840 24142
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19890 23216 19946 23225
rect 19890 23151 19946 23160
rect 19904 19854 19932 23151
rect 20088 22710 20116 23462
rect 20076 22704 20128 22710
rect 20076 22646 20128 22652
rect 19982 22264 20038 22273
rect 19982 22199 19984 22208
rect 20036 22199 20038 22208
rect 19984 22170 20036 22176
rect 20088 22094 20116 22646
rect 20272 22098 20300 26200
rect 20812 25560 20864 25566
rect 20812 25502 20864 25508
rect 20824 24070 20852 25502
rect 20916 24274 20944 26200
rect 21560 24410 21588 26200
rect 21548 24404 21600 24410
rect 21548 24346 21600 24352
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 21916 24200 21968 24206
rect 21968 24148 22140 24154
rect 21916 24142 22140 24148
rect 20812 24064 20864 24070
rect 20812 24006 20864 24012
rect 21456 23792 21508 23798
rect 21456 23734 21508 23740
rect 20352 23656 20404 23662
rect 20352 23598 20404 23604
rect 20364 23186 20392 23598
rect 20352 23180 20404 23186
rect 20404 23140 20484 23168
rect 20352 23122 20404 23128
rect 20352 23044 20404 23050
rect 20352 22986 20404 22992
rect 20364 22778 20392 22986
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 19996 22066 20116 22094
rect 20168 22092 20220 22098
rect 19996 20874 20024 22066
rect 20168 22034 20220 22040
rect 20260 22092 20312 22098
rect 20260 22034 20312 22040
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 20088 21593 20116 21830
rect 20180 21604 20208 22034
rect 20456 21672 20484 23140
rect 21468 23118 21496 23734
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 21468 22642 21496 23054
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 20536 21956 20588 21962
rect 20536 21898 20588 21904
rect 20548 21865 20576 21898
rect 20534 21856 20590 21865
rect 20534 21791 20590 21800
rect 20364 21644 20484 21672
rect 20536 21684 20588 21690
rect 20260 21616 20312 21622
rect 20074 21584 20130 21593
rect 20180 21576 20260 21604
rect 20260 21558 20312 21564
rect 20074 21519 20130 21528
rect 20364 21010 20392 21644
rect 20536 21626 20588 21632
rect 20548 21418 20576 21626
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 20536 21412 20588 21418
rect 20456 21372 20536 21400
rect 20456 21146 20484 21372
rect 20536 21354 20588 21360
rect 20904 21412 20956 21418
rect 20904 21354 20956 21360
rect 20444 21140 20496 21146
rect 20720 21140 20772 21146
rect 20444 21082 20496 21088
rect 20548 21100 20720 21128
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 20074 20768 20130 20777
rect 20074 20703 20130 20712
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19800 18284 19852 18290
rect 19800 18226 19852 18232
rect 19904 17105 19932 19654
rect 19996 19174 20024 20334
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 19996 18970 20024 19110
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19890 17096 19946 17105
rect 19890 17031 19946 17040
rect 19798 16552 19854 16561
rect 19798 16487 19854 16496
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19812 13802 19840 16487
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19996 15434 20024 15642
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 19800 13796 19852 13802
rect 19800 13738 19852 13744
rect 19996 13705 20024 15370
rect 20088 13938 20116 20703
rect 20548 20262 20576 21100
rect 20720 21082 20772 21088
rect 20812 21072 20864 21078
rect 20640 21020 20812 21026
rect 20640 21014 20864 21020
rect 20640 20998 20852 21014
rect 20640 20806 20668 20998
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 20618 20760 20742
rect 20640 20590 20760 20618
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 19922 20576 20198
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20640 19514 20668 20590
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20180 18426 20208 19110
rect 20364 18426 20392 19246
rect 20640 18698 20668 19450
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 20180 17626 20208 18158
rect 20180 17598 20300 17626
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20180 17338 20208 17478
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20272 17134 20300 17598
rect 20350 17232 20406 17241
rect 20350 17167 20406 17176
rect 20260 17128 20312 17134
rect 20260 17070 20312 17076
rect 20272 16794 20300 17070
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 20166 16688 20222 16697
rect 20166 16623 20222 16632
rect 20180 16114 20208 16623
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19982 13696 20038 13705
rect 19982 13631 20038 13640
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 20088 12306 20116 12718
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20260 11892 20312 11898
rect 20364 11880 20392 17167
rect 20732 16538 20760 20198
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20824 19514 20852 19722
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20812 18896 20864 18902
rect 20812 18838 20864 18844
rect 20824 18222 20852 18838
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20640 16510 20760 16538
rect 20640 15910 20668 16510
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20640 15162 20668 15506
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20442 13424 20498 13433
rect 20442 13359 20498 13368
rect 20456 12345 20484 13359
rect 20732 12850 20760 16390
rect 20824 16250 20852 16662
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20916 15994 20944 21354
rect 21100 20942 21128 21558
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21100 20466 21128 20878
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 21192 18834 21220 20946
rect 21468 20602 21496 21286
rect 21560 20942 21588 24142
rect 21928 24126 22140 24142
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21548 19984 21600 19990
rect 21468 19944 21548 19972
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21272 18080 21324 18086
rect 21270 18048 21272 18057
rect 21324 18048 21326 18057
rect 21270 17983 21326 17992
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 21008 17105 21036 17478
rect 20994 17096 21050 17105
rect 20994 17031 21050 17040
rect 20996 16516 21048 16522
rect 20996 16458 21048 16464
rect 20824 15966 20944 15994
rect 20824 14414 20852 15966
rect 20902 15872 20958 15881
rect 20902 15807 20958 15816
rect 20916 15026 20944 15807
rect 21008 15502 21036 16458
rect 21100 16250 21128 17614
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21192 16794 21220 17478
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20902 14784 20958 14793
rect 20902 14719 20958 14728
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20916 12889 20944 14719
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21100 12918 21128 14010
rect 21192 13734 21220 16730
rect 21284 16658 21312 17070
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 21376 15910 21404 19654
rect 21468 18834 21496 19944
rect 21548 19926 21600 19932
rect 21652 19854 21680 20266
rect 21640 19848 21692 19854
rect 21640 19790 21692 19796
rect 21652 19446 21680 19790
rect 21744 19446 21772 23666
rect 21824 23588 21876 23594
rect 21824 23530 21876 23536
rect 21836 22982 21864 23530
rect 21824 22976 21876 22982
rect 21824 22918 21876 22924
rect 21836 22438 21864 22918
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21928 21146 21956 23802
rect 21916 21140 21968 21146
rect 21916 21082 21968 21088
rect 21640 19440 21692 19446
rect 21640 19382 21692 19388
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21456 18828 21508 18834
rect 21456 18770 21508 18776
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21468 17338 21496 18022
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 21560 16726 21588 17274
rect 21548 16720 21600 16726
rect 21548 16662 21600 16668
rect 21456 16516 21508 16522
rect 21456 16458 21508 16464
rect 21468 16182 21496 16458
rect 21456 16176 21508 16182
rect 21456 16118 21508 16124
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21468 14890 21496 15302
rect 21560 15094 21588 15302
rect 21548 15088 21600 15094
rect 21548 15030 21600 15036
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21468 14346 21496 14826
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21652 14278 21680 18158
rect 21744 17921 21772 19382
rect 22112 18834 22140 24126
rect 22204 22273 22232 26200
rect 22560 24880 22612 24886
rect 22560 24822 22612 24828
rect 22284 24812 22336 24818
rect 22284 24754 22336 24760
rect 22296 23254 22324 24754
rect 22572 24410 22600 24822
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22284 23248 22336 23254
rect 22284 23190 22336 23196
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 23308 23066 23336 26302
rect 23478 26200 23534 27000
rect 24122 26200 24178 27000
rect 24766 26200 24822 27000
rect 25410 26200 25466 27000
rect 26054 26200 26110 27000
rect 26698 26200 26754 27000
rect 27342 26200 27398 27000
rect 27986 26330 28042 27000
rect 27986 26302 28580 26330
rect 27986 26200 28042 26302
rect 23492 24750 23520 26200
rect 24136 25566 24164 26200
rect 24124 25560 24176 25566
rect 24124 25502 24176 25508
rect 23480 24744 23532 24750
rect 23480 24686 23532 24692
rect 23940 24064 23992 24070
rect 23940 24006 23992 24012
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23768 23254 23796 23462
rect 23756 23248 23808 23254
rect 23756 23190 23808 23196
rect 23848 23112 23900 23118
rect 23308 23060 23848 23066
rect 23308 23054 23900 23060
rect 22296 22574 22324 23054
rect 23308 23038 23888 23054
rect 23388 22976 23440 22982
rect 23388 22918 23440 22924
rect 23400 22574 23428 22918
rect 23664 22704 23716 22710
rect 23664 22646 23716 22652
rect 22284 22568 22336 22574
rect 23388 22568 23440 22574
rect 22284 22510 22336 22516
rect 23308 22516 23388 22522
rect 23308 22510 23440 22516
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23308 22494 23428 22510
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22190 22264 22246 22273
rect 22950 22267 23258 22276
rect 22190 22199 22246 22208
rect 22836 22160 22888 22166
rect 23308 22114 23336 22494
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 22836 22102 22888 22108
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22480 21350 22508 21490
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22848 20602 22876 22102
rect 23216 22086 23336 22114
rect 23216 21554 23244 22086
rect 23400 22030 23428 22374
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23204 21548 23256 21554
rect 23204 21490 23256 21496
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23202 21040 23258 21049
rect 23202 20975 23204 20984
rect 23256 20975 23258 20984
rect 23204 20946 23256 20952
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22204 19417 22232 20198
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22560 19984 22612 19990
rect 22560 19926 22612 19932
rect 22928 19984 22980 19990
rect 22928 19926 22980 19932
rect 22572 19514 22600 19926
rect 22650 19544 22706 19553
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22560 19508 22612 19514
rect 22650 19479 22706 19488
rect 22560 19450 22612 19456
rect 22190 19408 22246 19417
rect 22190 19343 22246 19352
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21730 17912 21786 17921
rect 21730 17847 21786 17856
rect 21836 16561 21864 18566
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22190 18048 22246 18057
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 21822 16552 21878 16561
rect 21822 16487 21878 16496
rect 21928 15162 21956 17614
rect 22112 15570 22140 18022
rect 22190 17983 22246 17992
rect 22204 16250 22232 17983
rect 22282 17776 22338 17785
rect 22282 17711 22338 17720
rect 22296 17202 22324 17711
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22296 17105 22324 17138
rect 22282 17096 22338 17105
rect 22282 17031 22338 17040
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22204 15638 22232 16186
rect 22192 15632 22244 15638
rect 22192 15574 22244 15580
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22008 15496 22060 15502
rect 22060 15444 22140 15450
rect 22008 15438 22140 15444
rect 22020 15422 22140 15438
rect 22112 15366 22140 15422
rect 22100 15360 22152 15366
rect 22296 15314 22324 17031
rect 22100 15302 22152 15308
rect 22204 15286 22324 15314
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 22112 14006 22140 14214
rect 22204 14006 22232 15286
rect 22284 15156 22336 15162
rect 22284 15098 22336 15104
rect 22296 14482 22324 15098
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 21376 13530 21404 13874
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21640 13252 21692 13258
rect 21640 13194 21692 13200
rect 21088 12912 21140 12918
rect 20902 12880 20958 12889
rect 20720 12844 20772 12850
rect 21088 12854 21140 12860
rect 20902 12815 20958 12824
rect 20720 12786 20772 12792
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 12434 20760 12582
rect 20732 12406 20852 12434
rect 20442 12336 20498 12345
rect 20442 12271 20498 12280
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20312 11852 20392 11880
rect 20260 11834 20312 11840
rect 20732 11830 20760 12038
rect 20824 11898 20852 12406
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19720 11082 19748 11630
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19720 10606 19748 11018
rect 20732 11014 20760 11766
rect 21468 11558 21496 12718
rect 21652 12102 21680 13194
rect 21836 12442 21864 13738
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 21824 12436 21876 12442
rect 22020 12434 22048 12922
rect 22112 12850 22140 13670
rect 22388 13569 22416 19450
rect 22664 19446 22692 19479
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 22940 19334 22968 19926
rect 22756 19306 22968 19334
rect 22466 18864 22522 18873
rect 22466 18799 22522 18808
rect 22480 18465 22508 18799
rect 22466 18456 22522 18465
rect 22466 18391 22522 18400
rect 22480 18358 22508 18391
rect 22468 18352 22520 18358
rect 22468 18294 22520 18300
rect 22652 18216 22704 18222
rect 22480 18176 22652 18204
rect 22480 17542 22508 18176
rect 22652 18158 22704 18164
rect 22756 18154 22784 19306
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22928 18624 22980 18630
rect 22928 18566 22980 18572
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 22744 18148 22796 18154
rect 22744 18090 22796 18096
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22480 14822 22508 17478
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22756 17066 22784 17274
rect 22848 17202 22876 18294
rect 22940 18290 22968 18566
rect 22928 18284 22980 18290
rect 22928 18226 22980 18232
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 22744 17060 22796 17066
rect 22744 17002 22796 17008
rect 22836 17060 22888 17066
rect 22836 17002 22888 17008
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22560 15972 22612 15978
rect 22560 15914 22612 15920
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22374 13560 22430 13569
rect 22374 13495 22430 13504
rect 22480 13462 22508 14758
rect 22468 13456 22520 13462
rect 22468 13398 22520 13404
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22204 12850 22232 13330
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 21824 12378 21876 12384
rect 21928 12406 22048 12434
rect 21928 12306 21956 12406
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 22204 12238 22232 12786
rect 22572 12714 22600 15914
rect 22664 15745 22692 16186
rect 22650 15736 22706 15745
rect 22650 15671 22706 15680
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22560 12708 22612 12714
rect 22560 12650 22612 12656
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 22204 11694 22232 12174
rect 22664 11830 22692 14418
rect 22756 13870 22784 16594
rect 22848 15502 22876 17002
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22928 16720 22980 16726
rect 22928 16662 22980 16668
rect 22940 16250 22968 16662
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22836 15496 22888 15502
rect 22836 15438 22888 15444
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22928 14612 22980 14618
rect 22928 14554 22980 14560
rect 22940 14006 22968 14554
rect 22928 14000 22980 14006
rect 22928 13942 22980 13948
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22652 11824 22704 11830
rect 22652 11766 22704 11772
rect 22192 11688 22244 11694
rect 22756 11642 22784 13806
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 23032 12850 23060 13262
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23308 11778 23336 21830
rect 23400 21554 23428 21966
rect 23492 21962 23520 22510
rect 23676 21962 23704 22646
rect 23952 22522 23980 24006
rect 24492 23792 24544 23798
rect 24492 23734 24544 23740
rect 24504 23050 24532 23734
rect 24688 23730 24716 24006
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 24780 23322 24808 26200
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25240 24274 25268 24686
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25424 24206 25452 26200
rect 26068 24818 26096 26200
rect 25964 24812 26016 24818
rect 25964 24754 26016 24760
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 25976 24682 26004 24754
rect 25872 24676 25924 24682
rect 25872 24618 25924 24624
rect 25964 24676 26016 24682
rect 25964 24618 26016 24624
rect 25780 24608 25832 24614
rect 25780 24550 25832 24556
rect 25792 24410 25820 24550
rect 25884 24410 25912 24618
rect 25780 24404 25832 24410
rect 25780 24346 25832 24352
rect 25872 24404 25924 24410
rect 25872 24346 25924 24352
rect 26712 24206 26740 26200
rect 27252 24404 27304 24410
rect 27252 24346 27304 24352
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 26700 24200 26752 24206
rect 26700 24142 26752 24148
rect 27158 24168 27214 24177
rect 27158 24103 27214 24112
rect 27172 24070 27200 24103
rect 25044 24064 25096 24070
rect 25044 24006 25096 24012
rect 25688 24064 25740 24070
rect 25688 24006 25740 24012
rect 26240 24064 26292 24070
rect 26240 24006 26292 24012
rect 27160 24064 27212 24070
rect 27160 24006 27212 24012
rect 25056 23866 25084 24006
rect 25044 23860 25096 23866
rect 25044 23802 25096 23808
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24872 23526 24900 23598
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24492 23044 24544 23050
rect 24492 22986 24544 22992
rect 24504 22642 24532 22986
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 24596 22574 24624 22918
rect 24676 22704 24728 22710
rect 24676 22646 24728 22652
rect 23768 22494 23980 22522
rect 24584 22568 24636 22574
rect 24584 22510 24636 22516
rect 23480 21956 23532 21962
rect 23480 21898 23532 21904
rect 23664 21956 23716 21962
rect 23664 21898 23716 21904
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23386 21040 23442 21049
rect 23386 20975 23442 20984
rect 23400 20534 23428 20975
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23386 20088 23442 20097
rect 23386 20023 23442 20032
rect 23400 19854 23428 20023
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23386 19680 23442 19689
rect 23492 19666 23520 20878
rect 23584 20398 23612 21830
rect 23662 21176 23718 21185
rect 23662 21111 23718 21120
rect 23676 21010 23704 21111
rect 23664 21004 23716 21010
rect 23664 20946 23716 20952
rect 23664 20800 23716 20806
rect 23662 20768 23664 20777
rect 23716 20768 23718 20777
rect 23662 20703 23718 20712
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23442 19638 23520 19666
rect 23386 19615 23442 19624
rect 23400 16726 23428 19615
rect 23584 19514 23612 19994
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23572 19304 23624 19310
rect 23572 19246 23624 19252
rect 23584 18766 23612 19246
rect 23676 18970 23704 19654
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23570 17640 23626 17649
rect 23570 17575 23626 17584
rect 23584 17202 23612 17575
rect 23768 17218 23796 22494
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23952 21622 23980 22374
rect 24688 21962 24716 22646
rect 24872 22030 24900 23462
rect 25700 23186 25728 24006
rect 26252 23905 26280 24006
rect 26238 23896 26294 23905
rect 27264 23866 27292 24346
rect 27356 23866 27384 26200
rect 28078 24712 28134 24721
rect 28078 24647 28134 24656
rect 28092 24342 28120 24647
rect 28080 24336 28132 24342
rect 28080 24278 28132 24284
rect 28356 24268 28408 24274
rect 28356 24210 28408 24216
rect 27436 24064 27488 24070
rect 27436 24006 27488 24012
rect 27712 24064 27764 24070
rect 27712 24006 27764 24012
rect 26238 23831 26294 23840
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 27344 23860 27396 23866
rect 27344 23802 27396 23808
rect 26608 23792 26660 23798
rect 27448 23746 27476 24006
rect 26608 23734 26660 23740
rect 25872 23656 25924 23662
rect 25872 23598 25924 23604
rect 25884 23322 25912 23598
rect 26240 23588 26292 23594
rect 26240 23530 26292 23536
rect 26252 23474 26280 23530
rect 26620 23526 26648 23734
rect 27068 23724 27120 23730
rect 27068 23666 27120 23672
rect 27356 23718 27476 23746
rect 26884 23656 26936 23662
rect 26884 23598 26936 23604
rect 26160 23446 26280 23474
rect 26608 23520 26660 23526
rect 26608 23462 26660 23468
rect 25872 23316 25924 23322
rect 25872 23258 25924 23264
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 25688 23180 25740 23186
rect 25688 23122 25740 23128
rect 25872 23180 25924 23186
rect 25872 23122 25924 23128
rect 24952 22976 25004 22982
rect 24952 22918 25004 22924
rect 24964 22094 24992 22918
rect 25148 22778 25176 23122
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 24964 22066 25084 22094
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24950 21992 25006 22001
rect 24676 21956 24728 21962
rect 24676 21898 24728 21904
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23860 19922 23888 20946
rect 24688 20398 24716 21422
rect 24872 20534 24900 21966
rect 24950 21927 25006 21936
rect 24964 20942 24992 21927
rect 25056 21865 25084 22066
rect 25136 22092 25188 22098
rect 25136 22034 25188 22040
rect 25042 21856 25098 21865
rect 25042 21791 25098 21800
rect 25056 21593 25084 21791
rect 25148 21690 25176 22034
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25240 21622 25268 22578
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25412 22432 25464 22438
rect 25412 22374 25464 22380
rect 25228 21616 25280 21622
rect 25042 21584 25098 21593
rect 25228 21558 25280 21564
rect 25042 21519 25098 21528
rect 24952 20936 25004 20942
rect 24952 20878 25004 20884
rect 24860 20528 24912 20534
rect 24860 20470 24912 20476
rect 25240 20398 25268 21558
rect 25332 21350 25360 22374
rect 25424 22166 25452 22374
rect 25412 22160 25464 22166
rect 25412 22102 25464 22108
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 25516 20618 25544 22578
rect 25700 21962 25728 23122
rect 25780 22976 25832 22982
rect 25780 22918 25832 22924
rect 25792 22094 25820 22918
rect 25884 22522 25912 23122
rect 25964 23112 26016 23118
rect 25964 23054 26016 23060
rect 25976 22658 26004 23054
rect 26160 22778 26188 23446
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 25976 22630 26188 22658
rect 26160 22574 26188 22630
rect 26056 22568 26108 22574
rect 25884 22516 26056 22522
rect 25884 22510 26108 22516
rect 26148 22568 26200 22574
rect 26148 22510 26200 22516
rect 25884 22494 26096 22510
rect 26620 22438 26648 23462
rect 26896 23168 26924 23598
rect 27080 23186 27108 23666
rect 27068 23180 27120 23186
rect 26896 23140 27068 23168
rect 27068 23122 27120 23128
rect 27356 23066 27384 23718
rect 27436 23316 27488 23322
rect 27436 23258 27488 23264
rect 27620 23316 27672 23322
rect 27620 23258 27672 23264
rect 27172 23038 27384 23066
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 27068 22160 27120 22166
rect 26712 22120 27068 22148
rect 25792 22066 25912 22094
rect 25780 22024 25832 22030
rect 25780 21966 25832 21972
rect 25688 21956 25740 21962
rect 25688 21898 25740 21904
rect 25594 21448 25650 21457
rect 25594 21383 25596 21392
rect 25648 21383 25650 21392
rect 25596 21354 25648 21360
rect 25792 21010 25820 21966
rect 25884 21729 25912 22066
rect 25964 21956 26016 21962
rect 25964 21898 26016 21904
rect 25870 21720 25926 21729
rect 25870 21655 25926 21664
rect 25976 21570 26004 21898
rect 26712 21690 26740 22120
rect 27068 22102 27120 22108
rect 26792 21956 26844 21962
rect 26792 21898 26844 21904
rect 26804 21690 26832 21898
rect 26700 21684 26752 21690
rect 26700 21626 26752 21632
rect 26792 21684 26844 21690
rect 26792 21626 26844 21632
rect 25884 21542 26004 21570
rect 25780 21004 25832 21010
rect 25780 20946 25832 20952
rect 25516 20590 25820 20618
rect 25594 20496 25650 20505
rect 25594 20431 25650 20440
rect 24676 20392 24728 20398
rect 24676 20334 24728 20340
rect 25228 20392 25280 20398
rect 25228 20334 25280 20340
rect 25240 20097 25268 20334
rect 25608 20233 25636 20431
rect 25688 20324 25740 20330
rect 25688 20266 25740 20272
rect 25594 20224 25650 20233
rect 25594 20159 25650 20168
rect 25226 20088 25282 20097
rect 25226 20023 25282 20032
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 24032 19780 24084 19786
rect 24032 19722 24084 19728
rect 24044 19514 24072 19722
rect 24032 19508 24084 19514
rect 24032 19450 24084 19456
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23860 18358 23888 18634
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23572 17196 23624 17202
rect 23572 17138 23624 17144
rect 23676 17190 23796 17218
rect 23388 16720 23440 16726
rect 23440 16668 23520 16674
rect 23388 16662 23520 16668
rect 23400 16646 23520 16662
rect 23492 16590 23520 16646
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 23400 15144 23428 16458
rect 23572 15360 23624 15366
rect 23572 15302 23624 15308
rect 23400 15116 23520 15144
rect 23492 14906 23520 15116
rect 23584 15094 23612 15302
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23400 14878 23520 14906
rect 23400 13394 23428 14878
rect 23584 14346 23612 15030
rect 23572 14340 23624 14346
rect 23572 14282 23624 14288
rect 23572 14068 23624 14074
rect 23572 14010 23624 14016
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23492 12986 23520 13330
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23308 11750 23428 11778
rect 22192 11630 22244 11636
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 10742 20760 10950
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19720 10130 19748 10542
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 20732 9994 20760 10678
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 21192 9926 21220 11018
rect 21468 10810 21496 11494
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 22100 10124 22152 10130
rect 22100 10066 22152 10072
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 21192 9518 21220 9862
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 22112 9110 22140 10066
rect 22100 9104 22152 9110
rect 22100 9046 22152 9052
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 22204 7954 22232 11630
rect 22664 11614 22784 11642
rect 23296 11688 23348 11694
rect 23296 11630 23348 11636
rect 22664 11218 22692 11614
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22664 10606 22692 11154
rect 22652 10600 22704 10606
rect 22652 10542 22704 10548
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23308 10266 23336 11630
rect 23400 10577 23428 11750
rect 23386 10568 23442 10577
rect 23386 10503 23442 10512
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23584 9654 23612 14010
rect 23676 12434 23704 17190
rect 23860 17134 23888 17478
rect 23848 17128 23900 17134
rect 23848 17070 23900 17076
rect 24136 16590 24164 19314
rect 24952 19304 25004 19310
rect 24952 19246 25004 19252
rect 24858 19000 24914 19009
rect 24858 18935 24914 18944
rect 24492 18692 24544 18698
rect 24492 18634 24544 18640
rect 24504 17882 24532 18634
rect 24872 18630 24900 18935
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24492 17876 24544 17882
rect 24492 17818 24544 17824
rect 24504 17762 24532 17818
rect 24412 17734 24532 17762
rect 24412 17678 24440 17734
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 24490 17640 24546 17649
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24228 17241 24256 17478
rect 24214 17232 24270 17241
rect 24214 17167 24270 17176
rect 24124 16584 24176 16590
rect 24124 16526 24176 16532
rect 24228 16454 24256 17167
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 24216 16448 24268 16454
rect 24216 16390 24268 16396
rect 23768 16250 23796 16390
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23768 14958 23796 15506
rect 23756 14952 23808 14958
rect 23756 14894 23808 14900
rect 23860 13802 23888 15982
rect 23940 15428 23992 15434
rect 23940 15370 23992 15376
rect 23952 15162 23980 15370
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 23952 15026 23980 15098
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23940 14272 23992 14278
rect 23940 14214 23992 14220
rect 23848 13796 23900 13802
rect 23848 13738 23900 13744
rect 23952 12782 23980 14214
rect 24032 13796 24084 13802
rect 24032 13738 24084 13744
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 23940 12640 23992 12646
rect 23940 12582 23992 12588
rect 23676 12406 23888 12434
rect 23860 10130 23888 12406
rect 23952 12170 23980 12582
rect 23940 12164 23992 12170
rect 23940 12106 23992 12112
rect 23952 11830 23980 12106
rect 24044 12102 24072 13738
rect 24136 13258 24164 15302
rect 24412 15094 24440 17614
rect 24490 17575 24546 17584
rect 24504 17202 24532 17575
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24688 15910 24716 18226
rect 24768 18080 24820 18086
rect 24768 18022 24820 18028
rect 24780 17746 24808 18022
rect 24768 17740 24820 17746
rect 24768 17682 24820 17688
rect 24780 17202 24808 17682
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24780 17082 24808 17138
rect 24780 17054 24900 17082
rect 24872 16114 24900 17054
rect 24964 16250 24992 19246
rect 25056 18358 25084 19314
rect 25332 18630 25360 19858
rect 25504 19780 25556 19786
rect 25504 19722 25556 19728
rect 25410 19272 25466 19281
rect 25410 19207 25466 19216
rect 25424 19174 25452 19207
rect 25412 19168 25464 19174
rect 25412 19110 25464 19116
rect 25320 18624 25372 18630
rect 25320 18566 25372 18572
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 24676 15904 24728 15910
rect 24676 15846 24728 15852
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24400 15088 24452 15094
rect 24400 15030 24452 15036
rect 24124 13252 24176 13258
rect 24124 13194 24176 13200
rect 24412 12850 24440 15030
rect 24596 13258 24624 15438
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24872 14414 24900 15370
rect 24964 15162 24992 16186
rect 25056 15502 25084 18294
rect 25148 17270 25176 18362
rect 25332 18222 25360 18566
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 25228 17604 25280 17610
rect 25228 17546 25280 17552
rect 25136 17264 25188 17270
rect 25136 17206 25188 17212
rect 25240 16726 25268 17546
rect 25228 16720 25280 16726
rect 25134 16688 25190 16697
rect 25228 16662 25280 16668
rect 25134 16623 25136 16632
rect 25188 16623 25190 16632
rect 25136 16594 25188 16600
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24860 14408 24912 14414
rect 25148 14385 25176 16594
rect 25226 16552 25282 16561
rect 25226 16487 25228 16496
rect 25280 16487 25282 16496
rect 25228 16458 25280 16464
rect 25240 14414 25268 16458
rect 25424 15502 25452 19110
rect 25516 16522 25544 19722
rect 25700 18698 25728 20266
rect 25792 19854 25820 20590
rect 25884 20262 25912 21542
rect 25976 21486 26004 21542
rect 25964 21480 26016 21486
rect 25964 21422 26016 21428
rect 25976 21134 26464 21162
rect 25976 21078 26004 21134
rect 25964 21072 26016 21078
rect 25964 21014 26016 21020
rect 26056 21004 26108 21010
rect 26056 20946 26108 20952
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25872 19848 25924 19854
rect 25872 19790 25924 19796
rect 25792 19174 25820 19790
rect 25884 19310 25912 19790
rect 25872 19304 25924 19310
rect 25872 19246 25924 19252
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25884 18850 25912 19246
rect 25792 18834 25912 18850
rect 25780 18828 25912 18834
rect 25832 18822 25912 18828
rect 25780 18770 25832 18776
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25884 17746 25912 18822
rect 26068 18358 26096 20946
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26252 20074 26280 20810
rect 26436 20534 26464 21134
rect 26804 20856 26832 21626
rect 27068 20868 27120 20874
rect 26804 20828 27068 20856
rect 27068 20810 27120 20816
rect 26424 20528 26476 20534
rect 26424 20470 26476 20476
rect 26252 20046 26372 20074
rect 26238 19952 26294 19961
rect 26238 19887 26240 19896
rect 26292 19887 26294 19896
rect 26240 19858 26292 19864
rect 26148 19780 26200 19786
rect 26148 19722 26200 19728
rect 26160 19242 26188 19722
rect 26344 19310 26372 20046
rect 26332 19304 26384 19310
rect 26332 19246 26384 19252
rect 26436 19242 26464 20470
rect 27080 20466 27108 20810
rect 27172 20777 27200 23038
rect 27448 22710 27476 23258
rect 27526 22808 27582 22817
rect 27632 22778 27660 23258
rect 27724 22982 27752 24006
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 28368 23474 28396 24210
rect 28552 23644 28580 26302
rect 28630 26200 28686 27000
rect 29274 26330 29330 27000
rect 29918 26330 29974 27000
rect 29274 26302 29592 26330
rect 29274 26200 29330 26302
rect 28644 24970 28672 26200
rect 28644 24942 28764 24970
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 28644 24206 28672 24754
rect 28632 24200 28684 24206
rect 28632 24142 28684 24148
rect 28736 24138 28764 24942
rect 29092 24744 29144 24750
rect 29092 24686 29144 24692
rect 28724 24132 28776 24138
rect 28724 24074 28776 24080
rect 29000 24064 29052 24070
rect 29000 24006 29052 24012
rect 29012 23882 29040 24006
rect 28828 23854 29040 23882
rect 28632 23656 28684 23662
rect 28552 23616 28632 23644
rect 28632 23598 28684 23604
rect 28724 23520 28776 23526
rect 28368 23446 28488 23474
rect 28724 23462 28776 23468
rect 28262 23352 28318 23361
rect 28262 23287 28318 23296
rect 28276 23186 28304 23287
rect 28264 23180 28316 23186
rect 28264 23122 28316 23128
rect 28356 23180 28408 23186
rect 28356 23122 28408 23128
rect 27712 22976 27764 22982
rect 27712 22918 27764 22924
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27526 22743 27582 22752
rect 27620 22772 27672 22778
rect 27436 22704 27488 22710
rect 27436 22646 27488 22652
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27252 22092 27304 22098
rect 27252 22034 27304 22040
rect 27264 21690 27292 22034
rect 27252 21684 27304 21690
rect 27252 21626 27304 21632
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 27158 20768 27214 20777
rect 27158 20703 27214 20712
rect 27172 20466 27200 20703
rect 27264 20602 27292 21286
rect 27252 20596 27304 20602
rect 27252 20538 27304 20544
rect 27068 20460 27120 20466
rect 27068 20402 27120 20408
rect 27160 20460 27212 20466
rect 27160 20402 27212 20408
rect 27080 19836 27108 20402
rect 27356 20262 27384 22578
rect 27448 22098 27476 22646
rect 27436 22092 27488 22098
rect 27436 22034 27488 22040
rect 27540 21078 27568 22743
rect 27620 22714 27672 22720
rect 28368 22642 28396 23122
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 27804 22500 27856 22506
rect 27804 22442 27856 22448
rect 27816 22030 27844 22442
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 27894 21584 27950 21593
rect 27894 21519 27896 21528
rect 27948 21519 27950 21528
rect 27896 21490 27948 21496
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 27528 21072 27580 21078
rect 27528 21014 27580 21020
rect 27724 20942 27752 21422
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 27712 20800 27764 20806
rect 27816 20754 27844 21422
rect 27908 20806 27936 21490
rect 28368 21486 28396 22578
rect 28460 22094 28488 23446
rect 28632 22976 28684 22982
rect 28736 22964 28764 23462
rect 28828 23361 28856 23854
rect 28908 23792 28960 23798
rect 28908 23734 28960 23740
rect 28814 23352 28870 23361
rect 28814 23287 28870 23296
rect 28684 22936 28764 22964
rect 28632 22918 28684 22924
rect 28736 22574 28764 22936
rect 28724 22568 28776 22574
rect 28724 22510 28776 22516
rect 28460 22066 28764 22094
rect 28356 21480 28408 21486
rect 28356 21422 28408 21428
rect 28368 21010 28396 21422
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 27764 20748 27844 20754
rect 27712 20742 27844 20748
rect 27896 20800 27948 20806
rect 27896 20742 27948 20748
rect 27724 20726 27844 20742
rect 27528 20460 27580 20466
rect 27528 20402 27580 20408
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27172 20058 27200 20198
rect 27160 20052 27212 20058
rect 27160 19994 27212 20000
rect 27252 19848 27304 19854
rect 27080 19808 27252 19836
rect 27252 19790 27304 19796
rect 26148 19236 26200 19242
rect 26148 19178 26200 19184
rect 26424 19236 26476 19242
rect 26424 19178 26476 19184
rect 26160 18970 26188 19178
rect 26148 18964 26200 18970
rect 26148 18906 26200 18912
rect 27068 18896 27120 18902
rect 27068 18838 27120 18844
rect 26608 18624 26660 18630
rect 26608 18566 26660 18572
rect 26700 18624 26752 18630
rect 26700 18566 26752 18572
rect 26056 18352 26108 18358
rect 26056 18294 26108 18300
rect 26620 17882 26648 18566
rect 26712 18290 26740 18566
rect 26700 18284 26752 18290
rect 26700 18226 26752 18232
rect 26424 17876 26476 17882
rect 26424 17818 26476 17824
rect 26608 17876 26660 17882
rect 26608 17818 26660 17824
rect 25872 17740 25924 17746
rect 25872 17682 25924 17688
rect 26436 17610 26464 17818
rect 26424 17604 26476 17610
rect 26424 17546 26476 17552
rect 26700 17604 26752 17610
rect 26700 17546 26752 17552
rect 26436 17270 26464 17546
rect 26424 17264 26476 17270
rect 25778 17232 25834 17241
rect 26424 17206 26476 17212
rect 25778 17167 25834 17176
rect 25792 16794 25820 17167
rect 26712 17134 26740 17546
rect 26700 17128 26752 17134
rect 26700 17070 26752 17076
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25700 15570 25728 16594
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25228 14408 25280 14414
rect 24860 14350 24912 14356
rect 25134 14376 25190 14385
rect 25228 14350 25280 14356
rect 25700 14346 25728 15506
rect 25792 15434 25820 16730
rect 27080 16658 27108 18838
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 27172 17542 27200 18702
rect 27264 18698 27292 19790
rect 27252 18692 27304 18698
rect 27252 18634 27304 18640
rect 27160 17536 27212 17542
rect 27160 17478 27212 17484
rect 27160 17264 27212 17270
rect 27264 17218 27292 18634
rect 27212 17212 27292 17218
rect 27160 17206 27292 17212
rect 27172 17190 27292 17206
rect 27264 16810 27292 17190
rect 27172 16782 27292 16810
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27172 16182 27200 16782
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27160 16176 27212 16182
rect 27160 16118 27212 16124
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 25780 15428 25832 15434
rect 25780 15370 25832 15376
rect 25792 14414 25820 15370
rect 25780 14408 25832 14414
rect 25780 14350 25832 14356
rect 26160 14346 26188 15438
rect 27172 15094 27200 16118
rect 27264 16046 27292 16594
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 27160 15088 27212 15094
rect 27160 15030 27212 15036
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26620 14482 26648 14758
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 25134 14311 25190 14320
rect 25688 14340 25740 14346
rect 25148 14278 25176 14311
rect 25688 14282 25740 14288
rect 26148 14340 26200 14346
rect 26148 14282 26200 14288
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 24872 14006 24900 14214
rect 25792 14074 25820 14214
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 24860 14000 24912 14006
rect 24860 13942 24912 13948
rect 25136 13728 25188 13734
rect 25136 13670 25188 13676
rect 24584 13252 24636 13258
rect 24584 13194 24636 13200
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24412 12646 24440 12786
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 24044 11898 24072 12038
rect 25148 11898 25176 13670
rect 26884 13252 26936 13258
rect 26884 13194 26936 13200
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 25136 11892 25188 11898
rect 25136 11834 25188 11840
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22192 7948 22244 7954
rect 22192 7890 22244 7896
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20916 5710 20944 6734
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22112 5778 22140 6598
rect 22480 5914 22508 7754
rect 22572 7750 22600 9454
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23952 8242 23980 11766
rect 26896 11218 26924 13194
rect 26884 11212 26936 11218
rect 26884 11154 26936 11160
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 24872 8945 24900 10406
rect 24858 8936 24914 8945
rect 24858 8871 24914 8880
rect 23860 8214 23980 8242
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23860 7818 23888 8214
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 23848 7812 23900 7818
rect 23848 7754 23900 7760
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22572 6322 22600 7686
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 23952 7002 23980 8026
rect 23940 6996 23992 7002
rect 23940 6938 23992 6944
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 24780 5778 24808 6054
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 24768 5772 24820 5778
rect 24768 5714 24820 5720
rect 20904 5704 20956 5710
rect 20904 5646 20956 5652
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 17420 4826 17448 5578
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17420 2990 17448 4762
rect 17696 4486 17724 5102
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17696 3126 17724 4422
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17880 3058 17908 4966
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 20548 3058 20576 4966
rect 20916 4622 20944 5646
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21376 5234 21404 5510
rect 22112 5234 22140 5714
rect 25504 5636 25556 5642
rect 25504 5578 25556 5584
rect 27068 5636 27120 5642
rect 27068 5578 27120 5584
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 17420 800 17448 2450
rect 17512 2446 17540 2790
rect 20088 2446 20116 2790
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20180 1170 20208 2450
rect 22020 2446 22048 2790
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 25516 2650 25544 5578
rect 27080 5370 27108 5578
rect 27068 5364 27120 5370
rect 27068 5306 27120 5312
rect 25964 5024 26016 5030
rect 25964 4966 26016 4972
rect 25976 4554 26004 4966
rect 27356 4554 27384 20198
rect 27540 19990 27568 20402
rect 27816 20058 27844 20726
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 28368 20466 28396 20946
rect 28448 20936 28500 20942
rect 28540 20936 28592 20942
rect 28448 20878 28500 20884
rect 28538 20904 28540 20913
rect 28592 20904 28594 20913
rect 28356 20460 28408 20466
rect 28356 20402 28408 20408
rect 27804 20052 27856 20058
rect 27804 19994 27856 20000
rect 27528 19984 27580 19990
rect 27528 19926 27580 19932
rect 27436 19848 27488 19854
rect 27436 19790 27488 19796
rect 27448 18329 27476 19790
rect 27620 19712 27672 19718
rect 27620 19654 27672 19660
rect 27632 19553 27660 19654
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27618 19544 27674 19553
rect 27950 19547 28258 19556
rect 27618 19479 27674 19488
rect 27620 19372 27672 19378
rect 27620 19314 27672 19320
rect 27528 18828 27580 18834
rect 27528 18770 27580 18776
rect 27434 18320 27490 18329
rect 27434 18255 27490 18264
rect 27540 18086 27568 18770
rect 27632 18193 27660 19314
rect 28356 19304 28408 19310
rect 28356 19246 28408 19252
rect 28460 19258 28488 20878
rect 28538 20839 28594 20848
rect 28540 20800 28592 20806
rect 28540 20742 28592 20748
rect 28552 19394 28580 20742
rect 28552 19366 28672 19394
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 27724 18290 27752 18566
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 28368 18358 28396 19246
rect 28460 19230 28580 19258
rect 28448 19168 28500 19174
rect 28448 19110 28500 19116
rect 28356 18352 28408 18358
rect 28356 18294 28408 18300
rect 27712 18284 27764 18290
rect 27712 18226 27764 18232
rect 27804 18284 27856 18290
rect 27804 18226 27856 18232
rect 27618 18184 27674 18193
rect 27618 18119 27674 18128
rect 27528 18080 27580 18086
rect 27528 18022 27580 18028
rect 27540 17882 27568 18022
rect 27528 17876 27580 17882
rect 27528 17818 27580 17824
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27632 16590 27660 17818
rect 27816 17762 27844 18226
rect 27724 17746 27844 17762
rect 27712 17740 27844 17746
rect 27764 17734 27844 17740
rect 27712 17682 27764 17688
rect 27816 17202 27844 17734
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 28172 16992 28224 16998
rect 28172 16934 28224 16940
rect 28264 16992 28316 16998
rect 28264 16934 28316 16940
rect 28184 16590 28212 16934
rect 28276 16658 28304 16934
rect 28264 16652 28316 16658
rect 28264 16594 28316 16600
rect 27620 16584 27672 16590
rect 28172 16584 28224 16590
rect 27620 16526 27672 16532
rect 27816 16522 27936 16538
rect 28172 16526 28224 16532
rect 28460 16522 28488 19110
rect 27816 16516 27948 16522
rect 27816 16510 27896 16516
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 27540 12209 27568 14350
rect 27526 12200 27582 12209
rect 27526 12135 27582 12144
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 27448 6798 27476 9522
rect 27816 6914 27844 16510
rect 27896 16458 27948 16464
rect 28448 16516 28500 16522
rect 28448 16458 28500 16464
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 28552 13190 28580 19230
rect 28540 13184 28592 13190
rect 28540 13126 28592 13132
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 28644 12434 28672 19366
rect 28736 16561 28764 22066
rect 28814 20768 28870 20777
rect 28814 20703 28870 20712
rect 28828 18970 28856 20703
rect 28920 20602 28948 23734
rect 29000 23724 29052 23730
rect 29000 23666 29052 23672
rect 29012 23118 29040 23666
rect 29104 23254 29132 24686
rect 29564 24274 29592 26302
rect 29918 26302 30052 26330
rect 29918 26200 29974 26302
rect 29552 24268 29604 24274
rect 29552 24210 29604 24216
rect 29184 24064 29236 24070
rect 29184 24006 29236 24012
rect 29196 23798 29224 24006
rect 29736 23860 29788 23866
rect 29736 23802 29788 23808
rect 29184 23792 29236 23798
rect 29644 23792 29696 23798
rect 29184 23734 29236 23740
rect 29472 23752 29644 23780
rect 29092 23248 29144 23254
rect 29092 23190 29144 23196
rect 29184 23248 29236 23254
rect 29184 23190 29236 23196
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 29104 23050 29132 23190
rect 29196 23118 29224 23190
rect 29184 23112 29236 23118
rect 29184 23054 29236 23060
rect 29092 23044 29144 23050
rect 29092 22986 29144 22992
rect 29000 22432 29052 22438
rect 29000 22374 29052 22380
rect 29012 22094 29040 22374
rect 29196 22098 29224 23054
rect 29012 22066 29132 22094
rect 29000 21888 29052 21894
rect 29000 21830 29052 21836
rect 29012 21622 29040 21830
rect 29000 21616 29052 21622
rect 29000 21558 29052 21564
rect 29104 21486 29132 22066
rect 29184 22092 29236 22098
rect 29184 22034 29236 22040
rect 29184 21956 29236 21962
rect 29184 21898 29236 21904
rect 29092 21480 29144 21486
rect 29092 21422 29144 21428
rect 28998 20632 29054 20641
rect 28908 20596 28960 20602
rect 28998 20567 29054 20576
rect 28908 20538 28960 20544
rect 29012 20233 29040 20567
rect 29196 20505 29224 21898
rect 29368 20936 29420 20942
rect 29368 20878 29420 20884
rect 29182 20496 29238 20505
rect 29182 20431 29238 20440
rect 28998 20224 29054 20233
rect 28998 20159 29054 20168
rect 28816 18964 28868 18970
rect 28816 18906 28868 18912
rect 29090 18864 29146 18873
rect 29090 18799 29146 18808
rect 29104 18766 29132 18799
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 29092 18760 29144 18766
rect 29092 18702 29144 18708
rect 28816 17672 28868 17678
rect 28814 17640 28816 17649
rect 28868 17640 28870 17649
rect 28814 17575 28870 17584
rect 28722 16552 28778 16561
rect 28722 16487 28778 16496
rect 29012 16153 29040 18702
rect 28998 16144 29054 16153
rect 28998 16079 29054 16088
rect 29380 15609 29408 20878
rect 29472 19009 29500 23752
rect 29644 23734 29696 23740
rect 29748 23322 29776 23802
rect 30024 23730 30052 26302
rect 30562 26200 30618 27000
rect 31206 26200 31262 27000
rect 31850 26200 31906 27000
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26200 33838 27000
rect 34426 26200 34482 27000
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26330 36414 27000
rect 37002 26330 37058 27000
rect 36358 26302 36676 26330
rect 36358 26200 36414 26302
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30012 23724 30064 23730
rect 30012 23666 30064 23672
rect 30288 23656 30340 23662
rect 30288 23598 30340 23604
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 30012 23316 30064 23322
rect 30012 23258 30064 23264
rect 29552 22976 29604 22982
rect 29552 22918 29604 22924
rect 29564 20777 29592 22918
rect 30024 22710 30052 23258
rect 30012 22704 30064 22710
rect 30012 22646 30064 22652
rect 29920 22500 29972 22506
rect 29920 22442 29972 22448
rect 29644 22092 29696 22098
rect 29932 22094 29960 22442
rect 29932 22066 30052 22094
rect 29644 22034 29696 22040
rect 29656 21570 29684 22034
rect 29736 21616 29788 21622
rect 29656 21564 29736 21570
rect 29656 21558 29788 21564
rect 29656 21542 29776 21558
rect 29550 20768 29606 20777
rect 29550 20703 29606 20712
rect 29656 20534 29684 21542
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29644 20528 29696 20534
rect 29644 20470 29696 20476
rect 29656 19446 29684 20470
rect 29644 19440 29696 19446
rect 29840 19417 29868 20878
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 29644 19382 29696 19388
rect 29826 19408 29882 19417
rect 29458 19000 29514 19009
rect 29458 18935 29514 18944
rect 29472 18630 29500 18935
rect 29460 18624 29512 18630
rect 29460 18566 29512 18572
rect 29656 18290 29684 19382
rect 29826 19343 29882 19352
rect 29460 18284 29512 18290
rect 29460 18226 29512 18232
rect 29644 18284 29696 18290
rect 29644 18226 29696 18232
rect 29472 17746 29500 18226
rect 29460 17740 29512 17746
rect 29460 17682 29512 17688
rect 29472 17270 29500 17682
rect 29460 17264 29512 17270
rect 29460 17206 29512 17212
rect 29366 15600 29422 15609
rect 29366 15535 29422 15544
rect 28644 12406 28764 12434
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 28356 11076 28408 11082
rect 28356 11018 28408 11024
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 28368 8090 28396 11018
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27632 6886 27844 6914
rect 27436 6792 27488 6798
rect 27436 6734 27488 6740
rect 25964 4548 26016 4554
rect 25964 4490 26016 4496
rect 27344 4548 27396 4554
rect 27344 4490 27396 4496
rect 25504 2644 25556 2650
rect 25504 2586 25556 2592
rect 27448 2514 27476 6734
rect 27632 5574 27660 6886
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 28736 5642 28764 12406
rect 29932 11257 29960 19790
rect 30024 18834 30052 22066
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 30116 19174 30144 20402
rect 30208 20398 30236 21286
rect 30300 20641 30328 23598
rect 30392 22506 30420 24346
rect 30576 24206 30604 26200
rect 30564 24200 30616 24206
rect 30564 24142 30616 24148
rect 31220 23662 31248 26200
rect 31760 25492 31812 25498
rect 31760 25434 31812 25440
rect 31208 23656 31260 23662
rect 31208 23598 31260 23604
rect 31772 23610 31800 25434
rect 31864 23730 31892 26200
rect 32128 25356 32180 25362
rect 32128 25298 32180 25304
rect 32036 25152 32088 25158
rect 32036 25094 32088 25100
rect 31944 24268 31996 24274
rect 31944 24210 31996 24216
rect 31852 23724 31904 23730
rect 31852 23666 31904 23672
rect 31024 23588 31076 23594
rect 31772 23582 31892 23610
rect 31024 23530 31076 23536
rect 30564 23520 30616 23526
rect 30564 23462 30616 23468
rect 30380 22500 30432 22506
rect 30380 22442 30432 22448
rect 30576 21185 30604 23462
rect 31036 22710 31064 23530
rect 31760 23520 31812 23526
rect 31760 23462 31812 23468
rect 31116 23248 31168 23254
rect 31116 23190 31168 23196
rect 31128 22710 31156 23190
rect 31484 22976 31536 22982
rect 31484 22918 31536 22924
rect 31496 22778 31524 22918
rect 31484 22772 31536 22778
rect 31484 22714 31536 22720
rect 31024 22704 31076 22710
rect 31024 22646 31076 22652
rect 31116 22704 31168 22710
rect 31116 22646 31168 22652
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30656 21344 30708 21350
rect 30656 21286 30708 21292
rect 30562 21176 30618 21185
rect 30668 21146 30696 21286
rect 30562 21111 30618 21120
rect 30656 21140 30708 21146
rect 30656 21082 30708 21088
rect 30286 20632 30342 20641
rect 30286 20567 30342 20576
rect 30196 20392 30248 20398
rect 30196 20334 30248 20340
rect 30288 20256 30340 20262
rect 30288 20198 30340 20204
rect 30104 19168 30156 19174
rect 30104 19110 30156 19116
rect 30012 18828 30064 18834
rect 30012 18770 30064 18776
rect 30024 17746 30052 18770
rect 30116 18222 30144 19110
rect 30300 18698 30328 20198
rect 30944 19242 30972 22578
rect 31496 22166 31524 22714
rect 31668 22500 31720 22506
rect 31668 22442 31720 22448
rect 31576 22432 31628 22438
rect 31576 22374 31628 22380
rect 31588 22166 31616 22374
rect 31484 22160 31536 22166
rect 31484 22102 31536 22108
rect 31576 22160 31628 22166
rect 31680 22137 31708 22442
rect 31576 22102 31628 22108
rect 31666 22128 31722 22137
rect 31666 22063 31722 22072
rect 31300 21888 31352 21894
rect 31484 21888 31536 21894
rect 31352 21836 31432 21842
rect 31300 21830 31432 21836
rect 31484 21830 31536 21836
rect 31312 21814 31432 21830
rect 31024 21548 31076 21554
rect 31024 21490 31076 21496
rect 31036 20806 31064 21490
rect 31300 20936 31352 20942
rect 31300 20878 31352 20884
rect 31024 20800 31076 20806
rect 31024 20742 31076 20748
rect 30932 19236 30984 19242
rect 30932 19178 30984 19184
rect 30288 18692 30340 18698
rect 30288 18634 30340 18640
rect 30380 18692 30432 18698
rect 30380 18634 30432 18640
rect 30392 18578 30420 18634
rect 30300 18550 30420 18578
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 30300 17785 30328 18550
rect 30944 18358 30972 19178
rect 30932 18352 30984 18358
rect 30932 18294 30984 18300
rect 30840 18216 30892 18222
rect 30840 18158 30892 18164
rect 30286 17776 30342 17785
rect 30012 17740 30064 17746
rect 30286 17711 30342 17720
rect 30012 17682 30064 17688
rect 30024 17134 30052 17682
rect 30852 17610 30880 18158
rect 30840 17604 30892 17610
rect 30840 17546 30892 17552
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30208 17338 30236 17478
rect 30196 17332 30248 17338
rect 30196 17274 30248 17280
rect 30104 17264 30156 17270
rect 30104 17206 30156 17212
rect 30012 17128 30064 17134
rect 30012 17070 30064 17076
rect 29918 11248 29974 11257
rect 29918 11183 29974 11192
rect 30116 11082 30144 17206
rect 30104 11076 30156 11082
rect 30104 11018 30156 11024
rect 31312 9081 31340 20878
rect 31404 19990 31432 21814
rect 31392 19984 31444 19990
rect 31392 19926 31444 19932
rect 31404 19718 31432 19926
rect 31392 19712 31444 19718
rect 31392 19654 31444 19660
rect 31298 9072 31354 9081
rect 31298 9007 31354 9016
rect 28908 5772 28960 5778
rect 28908 5714 28960 5720
rect 28724 5636 28776 5642
rect 28724 5578 28776 5584
rect 27620 5568 27672 5574
rect 27620 5510 27672 5516
rect 28356 5568 28408 5574
rect 28356 5510 28408 5516
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27804 4684 27856 4690
rect 27804 4626 27856 4632
rect 27528 4548 27580 4554
rect 27528 4490 27580 4496
rect 27540 3602 27568 4490
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 27816 2650 27844 4626
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 28368 3534 28396 5510
rect 28736 3670 28764 5578
rect 28816 5160 28868 5166
rect 28816 5102 28868 5108
rect 28828 4826 28856 5102
rect 28816 4820 28868 4826
rect 28816 4762 28868 4768
rect 28724 3664 28776 3670
rect 28724 3606 28776 3612
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28920 2650 28948 5714
rect 31404 5166 31432 19654
rect 31496 15473 31524 21830
rect 31772 21554 31800 23462
rect 31760 21548 31812 21554
rect 31760 21490 31812 21496
rect 31864 21146 31892 23582
rect 31956 23225 31984 24210
rect 31942 23216 31998 23225
rect 31942 23151 31998 23160
rect 32048 21690 32076 25094
rect 32140 23322 32168 25298
rect 32312 24676 32364 24682
rect 32312 24618 32364 24624
rect 32324 24410 32352 24618
rect 32312 24404 32364 24410
rect 32312 24346 32364 24352
rect 32508 23780 32536 26200
rect 33152 25242 33180 26200
rect 33416 25288 33468 25294
rect 33152 25214 33364 25242
rect 33416 25230 33468 25236
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 33336 24206 33364 25214
rect 33428 24410 33456 25230
rect 33416 24404 33468 24410
rect 33416 24346 33468 24352
rect 33796 24206 33824 26200
rect 34152 25220 34204 25226
rect 34152 25162 34204 25168
rect 34164 24410 34192 25162
rect 34152 24404 34204 24410
rect 34152 24346 34204 24352
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 33784 24200 33836 24206
rect 34440 24188 34468 26200
rect 34520 25424 34572 25430
rect 34520 25366 34572 25372
rect 34532 24410 34560 25366
rect 34520 24404 34572 24410
rect 34520 24346 34572 24352
rect 34610 24304 34666 24313
rect 34610 24239 34666 24248
rect 34520 24200 34572 24206
rect 34440 24160 34520 24188
rect 33784 24142 33836 24148
rect 34520 24142 34572 24148
rect 34520 24064 34572 24070
rect 34520 24006 34572 24012
rect 32588 23792 32640 23798
rect 32508 23752 32588 23780
rect 32588 23734 32640 23740
rect 34060 23724 34112 23730
rect 34060 23666 34112 23672
rect 34428 23724 34480 23730
rect 34428 23666 34480 23672
rect 32494 23624 32550 23633
rect 32494 23559 32550 23568
rect 32128 23316 32180 23322
rect 32128 23258 32180 23264
rect 32508 22778 32536 23559
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 33506 23080 33562 23089
rect 32680 23044 32732 23050
rect 33506 23015 33562 23024
rect 32680 22986 32732 22992
rect 32496 22772 32548 22778
rect 32496 22714 32548 22720
rect 32404 22636 32456 22642
rect 32404 22578 32456 22584
rect 32036 21684 32088 21690
rect 32036 21626 32088 21632
rect 32220 21548 32272 21554
rect 32220 21490 32272 21496
rect 31852 21140 31904 21146
rect 31852 21082 31904 21088
rect 31576 19916 31628 19922
rect 31576 19858 31628 19864
rect 31588 16658 31616 19858
rect 31576 16652 31628 16658
rect 31576 16594 31628 16600
rect 31482 15464 31538 15473
rect 31482 15399 31538 15408
rect 32232 13977 32260 21490
rect 32312 20868 32364 20874
rect 32312 20810 32364 20816
rect 32218 13968 32274 13977
rect 32218 13903 32274 13912
rect 32324 13297 32352 20810
rect 32310 13288 32366 13297
rect 32310 13223 32366 13232
rect 32416 11801 32444 22578
rect 32588 22024 32640 22030
rect 32588 21966 32640 21972
rect 32600 19825 32628 21966
rect 32586 19816 32642 19825
rect 32586 19751 32642 19760
rect 32692 15065 32720 22986
rect 33520 22982 33548 23015
rect 32772 22976 32824 22982
rect 32772 22918 32824 22924
rect 33508 22976 33560 22982
rect 33508 22918 33560 22924
rect 32784 22234 32812 22918
rect 33324 22636 33376 22642
rect 33324 22578 33376 22584
rect 33508 22636 33560 22642
rect 33508 22578 33560 22584
rect 33230 22536 33286 22545
rect 33230 22471 33286 22480
rect 33244 22438 33272 22471
rect 33232 22432 33284 22438
rect 33232 22374 33284 22380
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 32772 22228 32824 22234
rect 32772 22170 32824 22176
rect 32864 22024 32916 22030
rect 32864 21966 32916 21972
rect 32678 15056 32734 15065
rect 32678 14991 32734 15000
rect 32402 11792 32458 11801
rect 32402 11727 32458 11736
rect 31668 11076 31720 11082
rect 31668 11018 31720 11024
rect 31680 9382 31708 11018
rect 32876 10470 32904 21966
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 33336 13433 33364 22578
rect 33416 21548 33468 21554
rect 33416 21490 33468 21496
rect 33428 18737 33456 21490
rect 33520 20369 33548 22578
rect 33506 20360 33562 20369
rect 33506 20295 33562 20304
rect 33414 18728 33470 18737
rect 33414 18663 33470 18672
rect 34072 16017 34100 23666
rect 34152 23044 34204 23050
rect 34152 22986 34204 22992
rect 34164 21690 34192 22986
rect 34244 22976 34296 22982
rect 34244 22918 34296 22924
rect 34256 22681 34284 22918
rect 34242 22672 34298 22681
rect 34242 22607 34298 22616
rect 34336 22432 34388 22438
rect 34336 22374 34388 22380
rect 34152 21684 34204 21690
rect 34152 21626 34204 21632
rect 34058 16008 34114 16017
rect 34058 15943 34114 15952
rect 33322 13424 33378 13433
rect 33322 13359 33378 13368
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32864 10464 32916 10470
rect 32864 10406 32916 10412
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 34348 9489 34376 22374
rect 34440 18902 34468 23666
rect 34532 22098 34560 24006
rect 34624 23798 34652 24239
rect 35084 24206 35112 26200
rect 35162 24848 35218 24857
rect 35162 24783 35218 24792
rect 35072 24200 35124 24206
rect 35072 24142 35124 24148
rect 34704 24132 34756 24138
rect 34704 24074 34756 24080
rect 34612 23792 34664 23798
rect 34612 23734 34664 23740
rect 34520 22092 34572 22098
rect 34520 22034 34572 22040
rect 34716 20602 34744 24074
rect 35176 23866 35204 24783
rect 35728 24188 35756 26200
rect 35900 25016 35952 25022
rect 35900 24958 35952 24964
rect 35912 24410 35940 24958
rect 35900 24404 35952 24410
rect 35900 24346 35952 24352
rect 35900 24200 35952 24206
rect 35728 24160 35900 24188
rect 35900 24142 35952 24148
rect 35164 23860 35216 23866
rect 35164 23802 35216 23808
rect 35992 23792 36044 23798
rect 35990 23760 35992 23769
rect 36044 23760 36046 23769
rect 35072 23724 35124 23730
rect 35072 23666 35124 23672
rect 35808 23724 35860 23730
rect 36648 23730 36676 26302
rect 37002 26302 37228 26330
rect 37002 26200 37058 26302
rect 37200 24188 37228 26302
rect 37646 26200 37702 27000
rect 38290 26330 38346 27000
rect 38934 26330 38990 27000
rect 39578 26330 39634 27000
rect 40222 26330 40278 27000
rect 40866 26330 40922 27000
rect 38290 26302 38516 26330
rect 38290 26200 38346 26302
rect 37280 24200 37332 24206
rect 37200 24160 37280 24188
rect 37280 24142 37332 24148
rect 37660 23730 37688 26200
rect 38488 24206 38516 26302
rect 38934 26302 39252 26330
rect 38934 26200 38990 26302
rect 38660 24948 38712 24954
rect 38660 24890 38712 24896
rect 38672 24206 38700 24890
rect 39224 24206 39252 26302
rect 39578 26302 39988 26330
rect 39578 26200 39634 26302
rect 39304 25084 39356 25090
rect 39304 25026 39356 25032
rect 39316 24410 39344 25026
rect 39960 24834 39988 26302
rect 40222 26302 40632 26330
rect 40222 26200 40278 26302
rect 39960 24806 40080 24834
rect 39304 24404 39356 24410
rect 39304 24346 39356 24352
rect 40052 24274 40080 24806
rect 40040 24268 40092 24274
rect 40040 24210 40092 24216
rect 40604 24206 40632 26302
rect 40866 26302 41184 26330
rect 40866 26200 40922 26302
rect 38476 24200 38528 24206
rect 38476 24142 38528 24148
rect 38660 24200 38712 24206
rect 38660 24142 38712 24148
rect 39212 24200 39264 24206
rect 39212 24142 39264 24148
rect 40592 24200 40644 24206
rect 40592 24142 40644 24148
rect 40040 24132 40092 24138
rect 40040 24074 40092 24080
rect 38660 24064 38712 24070
rect 38660 24006 38712 24012
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 35990 23695 36046 23704
rect 36636 23724 36688 23730
rect 35808 23666 35860 23672
rect 36636 23666 36688 23672
rect 37648 23724 37700 23730
rect 37648 23666 37700 23672
rect 34704 20596 34756 20602
rect 34704 20538 34756 20544
rect 35084 19514 35112 23666
rect 35256 23520 35308 23526
rect 35256 23462 35308 23468
rect 35268 21622 35296 23462
rect 35256 21616 35308 21622
rect 35256 21558 35308 21564
rect 35072 19508 35124 19514
rect 35072 19450 35124 19456
rect 34428 18896 34480 18902
rect 34428 18838 34480 18844
rect 35820 14414 35848 23666
rect 37188 23656 37240 23662
rect 37188 23598 37240 23604
rect 37200 16697 37228 23598
rect 37740 23520 37792 23526
rect 37740 23462 37792 23468
rect 37752 18426 37780 23462
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 38672 20913 38700 24006
rect 40052 23254 40080 24074
rect 41156 23730 41184 26302
rect 41510 26200 41566 27000
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43442 26330 43498 27000
rect 43442 26302 43668 26330
rect 43442 26200 43498 26302
rect 41524 24188 41552 26200
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 41604 24200 41656 24206
rect 41524 24160 41604 24188
rect 41604 24142 41656 24148
rect 43640 23798 43668 26302
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26330 45430 27000
rect 45374 26302 45508 26330
rect 45374 26200 45430 26302
rect 43628 23792 43680 23798
rect 43628 23734 43680 23740
rect 41144 23724 41196 23730
rect 44100 23712 44128 26200
rect 44744 24206 44772 26200
rect 45480 24290 45508 26302
rect 46018 26200 46074 27000
rect 46662 26200 46718 27000
rect 47306 26200 47362 27000
rect 47950 26200 48006 27000
rect 48594 26200 48650 27000
rect 45480 24262 45600 24290
rect 45572 24206 45600 24262
rect 46032 24206 46060 26200
rect 44732 24200 44784 24206
rect 44732 24142 44784 24148
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 46020 24200 46072 24206
rect 46020 24142 46072 24148
rect 45376 24064 45428 24070
rect 45376 24006 45428 24012
rect 46112 24064 46164 24070
rect 46112 24006 46164 24012
rect 46388 24064 46440 24070
rect 46388 24006 46440 24012
rect 44180 23724 44232 23730
rect 44100 23684 44180 23712
rect 41144 23666 41196 23672
rect 44180 23666 44232 23672
rect 41328 23520 41380 23526
rect 41328 23462 41380 23468
rect 40040 23248 40092 23254
rect 40040 23190 40092 23196
rect 40052 22710 40080 23190
rect 40040 22704 40092 22710
rect 40040 22646 40092 22652
rect 39672 22432 39724 22438
rect 39672 22374 39724 22380
rect 39684 22166 39712 22374
rect 39672 22160 39724 22166
rect 39672 22102 39724 22108
rect 38658 20904 38714 20913
rect 38658 20839 38714 20848
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 41340 19786 41368 23462
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 42800 22976 42852 22982
rect 42800 22918 42852 22924
rect 41328 19780 41380 19786
rect 41328 19722 41380 19728
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 37740 18420 37792 18426
rect 37740 18362 37792 18368
rect 42812 17610 42840 22918
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 45388 18902 45416 24006
rect 46124 23866 46152 24006
rect 46112 23860 46164 23866
rect 46112 23802 46164 23808
rect 45376 18896 45428 18902
rect 45376 18838 45428 18844
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 42800 17604 42852 17610
rect 42800 17546 42852 17552
rect 46400 17542 46428 24006
rect 46676 23730 46704 26200
rect 47320 24206 47348 26200
rect 47964 24206 47992 26200
rect 48318 24848 48374 24857
rect 48318 24783 48374 24792
rect 47308 24200 47360 24206
rect 47308 24142 47360 24148
rect 47952 24200 48004 24206
rect 47952 24142 48004 24148
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 48332 23730 48360 24783
rect 46664 23724 46716 23730
rect 46664 23666 46716 23672
rect 48320 23724 48372 23730
rect 48320 23666 48372 23672
rect 46940 23520 46992 23526
rect 46940 23462 46992 23468
rect 48504 23520 48556 23526
rect 48504 23462 48556 23468
rect 46952 22001 46980 23462
rect 48412 22976 48464 22982
rect 48412 22918 48464 22924
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 48424 22574 48452 22918
rect 48412 22568 48464 22574
rect 48412 22510 48464 22516
rect 46938 21992 46994 22001
rect 46938 21927 46994 21936
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 47860 21548 47912 21554
rect 47860 21490 47912 21496
rect 46388 17536 46440 17542
rect 46388 17478 46440 17484
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 37186 16688 37242 16697
rect 37186 16623 37242 16632
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 35808 14408 35860 14414
rect 35808 14350 35860 14356
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 47872 11082 47900 21490
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 48516 18698 48544 23462
rect 48608 23118 48636 26200
rect 48780 24064 48832 24070
rect 48780 24006 48832 24012
rect 48688 23520 48740 23526
rect 48688 23462 48740 23468
rect 48596 23112 48648 23118
rect 48596 23054 48648 23060
rect 48700 21457 48728 23462
rect 48686 21448 48742 21457
rect 48686 21383 48742 21392
rect 48504 18692 48556 18698
rect 48504 18634 48556 18640
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 48792 17241 48820 24006
rect 49054 23896 49110 23905
rect 49054 23831 49110 23840
rect 49068 23730 49096 23831
rect 49056 23724 49108 23730
rect 49056 23666 49108 23672
rect 49056 23112 49108 23118
rect 49056 23054 49108 23060
rect 49068 22953 49096 23054
rect 49054 22944 49110 22953
rect 49054 22879 49110 22888
rect 49056 22024 49108 22030
rect 49054 21992 49056 22001
rect 49108 21992 49110 22001
rect 49054 21927 49110 21936
rect 49240 21888 49292 21894
rect 49240 21830 49292 21836
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 49160 21049 49188 21422
rect 49146 21040 49202 21049
rect 49146 20975 49202 20984
rect 48778 17232 48834 17241
rect 48778 17167 48834 17176
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 49252 13870 49280 21830
rect 49240 13864 49292 13870
rect 49240 13806 49292 13812
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47860 11076 47912 11082
rect 47860 11018 47912 11024
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 34334 9480 34390 9489
rect 34334 9415 34390 9424
rect 31668 9376 31720 9382
rect 31668 9318 31720 9324
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 31392 5160 31444 5166
rect 31392 5102 31444 5108
rect 30392 3738 30420 5102
rect 33508 5092 33560 5098
rect 33508 5034 33560 5040
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 30380 3732 30432 3738
rect 30380 3674 30432 3680
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 33520 2650 33548 5034
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 41420 3732 41472 3738
rect 41420 3674 41472 3680
rect 38752 3460 38804 3466
rect 38752 3402 38804 3408
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 28908 2644 28960 2650
rect 28908 2586 28960 2592
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 27436 2508 27488 2514
rect 27436 2450 27488 2456
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 20088 1142 20208 1170
rect 20088 800 20116 1142
rect 22756 800 22784 2450
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 25424 800 25452 2382
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28092 870 28212 898
rect 28092 800 28120 870
rect 1504 734 1808 762
rect 4066 0 4122 800
rect 6734 0 6790 800
rect 9402 0 9458 800
rect 12070 0 12126 800
rect 14738 0 14794 800
rect 17406 0 17462 800
rect 20074 0 20130 800
rect 22742 0 22798 800
rect 25410 0 25466 800
rect 28078 0 28134 800
rect 28184 762 28212 870
rect 28368 762 28396 2382
rect 30760 800 30788 2382
rect 33428 800 33456 2382
rect 36096 800 36124 2382
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38764 800 38792 3402
rect 41432 800 41460 3674
rect 44088 3664 44140 3670
rect 44088 3606 44140 3612
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 44100 800 44128 3606
rect 46756 3596 46808 3602
rect 46756 3538 46808 3544
rect 46768 800 46796 3538
rect 49424 3528 49476 3534
rect 49424 3470 49476 3476
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49436 800 49464 3470
rect 28184 734 28396 762
rect 30746 0 30802 800
rect 33414 0 33470 800
rect 36082 0 36138 800
rect 38750 0 38806 800
rect 41418 0 41474 800
rect 44086 0 44142 800
rect 46754 0 46810 800
rect 49422 0 49478 800
<< via2 >>
rect 1490 24384 1546 24440
rect 938 10920 994 10976
rect 1306 20712 1362 20768
rect 1398 18672 1454 18728
rect 1766 19216 1822 19272
rect 1214 17040 1270 17096
rect 1306 16632 1362 16688
rect 2042 19896 2098 19952
rect 2042 18264 2098 18320
rect 1858 17584 1914 17640
rect 1306 16224 1362 16280
rect 1306 15816 1362 15872
rect 1306 15408 1362 15464
rect 1306 15000 1362 15056
rect 1306 14592 1362 14648
rect 1398 8880 1454 8936
rect 938 8472 994 8528
rect 1306 8064 1362 8120
rect 1582 13368 1638 13424
rect 1582 9696 1638 9752
rect 1858 14456 1914 14512
rect 1766 12844 1822 12880
rect 1766 12824 1768 12844
rect 1768 12824 1820 12844
rect 1820 12824 1822 12844
rect 1766 12552 1822 12608
rect 3330 25608 3386 25664
rect 3422 25200 3478 25256
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 3882 24792 3938 24848
rect 3422 23432 3478 23488
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2502 22752 2558 22808
rect 2686 21528 2742 21584
rect 2778 21120 2834 21176
rect 3606 22480 3662 22536
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 3422 22208 3478 22264
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2594 20440 2650 20496
rect 2502 17856 2558 17912
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2870 19488 2926 19544
rect 2778 19080 2834 19136
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2870 17720 2926 17776
rect 2778 17448 2834 17504
rect 3330 16904 3386 16960
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2778 14184 2834 14240
rect 2686 13776 2742 13832
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 3330 12960 3386 13016
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2778 12164 2834 12200
rect 2778 12144 2780 12164
rect 2780 12144 2832 12164
rect 2832 12144 2834 12164
rect 2870 12008 2926 12064
rect 2778 11212 2834 11248
rect 2778 11192 2780 11212
rect 2780 11192 2832 11212
rect 2832 11192 2834 11212
rect 3606 21664 3662 21720
rect 3974 23976 4030 24032
rect 3790 22072 3846 22128
rect 4802 24148 4804 24168
rect 4804 24148 4856 24168
rect 4856 24148 4858 24168
rect 4802 24112 4858 24148
rect 4066 23568 4122 23624
rect 4066 22072 4122 22128
rect 4158 20748 4160 20768
rect 4160 20748 4212 20768
rect 4212 20748 4214 20768
rect 4158 20712 4214 20748
rect 3882 20340 3884 20360
rect 3884 20340 3936 20360
rect 3936 20340 3938 20360
rect 3882 20304 3938 20340
rect 3882 17312 3938 17368
rect 3698 13932 3754 13968
rect 3698 13912 3700 13932
rect 3700 13912 3752 13932
rect 3752 13912 3754 13932
rect 3422 11736 3478 11792
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2870 10512 2926 10568
rect 2778 9288 2834 9344
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 3330 10104 3386 10160
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3514 11056 3570 11112
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 1766 7656 1822 7712
rect 4434 21936 4490 21992
rect 4066 17176 4122 17232
rect 4158 15816 4214 15872
rect 4342 16496 4398 16552
rect 4434 15272 4490 15328
rect 4986 23160 5042 23216
rect 4894 22888 4950 22944
rect 6642 23432 6698 23488
rect 4894 18672 4950 18728
rect 4710 15564 4766 15600
rect 4710 15544 4712 15564
rect 4712 15544 4764 15564
rect 4764 15544 4766 15564
rect 4894 15952 4950 16008
rect 4434 12280 4490 12336
rect 4710 12552 4766 12608
rect 4710 11328 4766 11384
rect 4158 9016 4214 9072
rect 5262 17312 5318 17368
rect 5354 17176 5410 17232
rect 5354 17076 5356 17096
rect 5356 17076 5408 17096
rect 5408 17076 5410 17096
rect 5354 17040 5410 17076
rect 5354 16632 5410 16688
rect 5078 15680 5134 15736
rect 5170 11056 5226 11112
rect 6366 21528 6422 21584
rect 6182 21256 6238 21312
rect 5630 18284 5686 18320
rect 5630 18264 5632 18284
rect 5632 18264 5684 18284
rect 5684 18264 5686 18284
rect 5814 18808 5870 18864
rect 5446 11756 5502 11792
rect 5446 11736 5448 11756
rect 5448 11736 5500 11756
rect 5500 11736 5502 11756
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 8114 23724 8170 23760
rect 8114 23704 8116 23724
rect 8116 23704 8168 23724
rect 8168 23704 8170 23724
rect 6826 23024 6882 23080
rect 6826 21392 6882 21448
rect 6642 19352 6698 19408
rect 7010 21972 7012 21992
rect 7012 21972 7064 21992
rect 7064 21972 7066 21992
rect 7010 21936 7066 21972
rect 6918 20576 6974 20632
rect 6918 20476 6920 20496
rect 6920 20476 6972 20496
rect 6972 20476 6974 20496
rect 6918 20440 6974 20476
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7286 20712 7342 20768
rect 7010 18672 7066 18728
rect 5998 9560 6054 9616
rect 6642 15428 6698 15464
rect 6642 15408 6644 15428
rect 6644 15408 6696 15428
rect 6696 15408 6698 15428
rect 6734 13640 6790 13696
rect 6366 9424 6422 9480
rect 2870 7248 2926 7304
rect 2778 6840 2834 6896
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 7102 16088 7158 16144
rect 7378 15564 7434 15600
rect 7378 15544 7380 15564
rect 7380 15544 7432 15564
rect 7432 15544 7434 15564
rect 7102 15408 7158 15464
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 9954 23568 10010 23624
rect 8298 18828 8354 18864
rect 8298 18808 8300 18828
rect 8300 18808 8352 18828
rect 8352 18808 8354 18828
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 8482 18264 8538 18320
rect 8022 17584 8078 17640
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 8206 16532 8208 16552
rect 8208 16532 8260 16552
rect 8260 16532 8262 16552
rect 8206 16496 8262 16532
rect 7562 15544 7618 15600
rect 7746 15408 7802 15464
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 8206 15680 8262 15736
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7746 15000 7802 15056
rect 7470 12280 7526 12336
rect 7286 11636 7288 11656
rect 7288 11636 7340 11656
rect 7340 11636 7342 11656
rect 7286 11600 7342 11636
rect 7102 11056 7158 11112
rect 7194 9832 7250 9888
rect 1214 6432 1270 6488
rect 938 6024 994 6080
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 938 5652 940 5672
rect 940 5652 992 5672
rect 992 5652 994 5672
rect 938 5616 994 5652
rect 938 5228 994 5264
rect 938 5208 940 5228
rect 940 5208 992 5228
rect 992 5208 994 5228
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 938 4800 994 4856
rect 1766 4392 1822 4448
rect 1306 3984 1362 4040
rect 938 3576 994 3632
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 1214 3168 1270 3224
rect 938 2760 994 2816
rect 938 2388 940 2408
rect 940 2388 992 2408
rect 992 2388 994 2408
rect 938 2352 994 2388
rect 2778 1944 2834 2000
rect 8482 17212 8484 17232
rect 8484 17212 8536 17232
rect 8536 17212 8538 17232
rect 8482 17176 8538 17212
rect 8390 15816 8446 15872
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 8298 13676 8300 13696
rect 8300 13676 8352 13696
rect 8352 13676 8354 13696
rect 8298 13640 8354 13676
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7746 11056 7802 11112
rect 7562 10648 7618 10704
rect 7470 8916 7472 8936
rect 7472 8916 7524 8936
rect 7524 8916 7526 8936
rect 7470 8880 7526 8916
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7930 9968 7986 10024
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 8850 10512 8906 10568
rect 9310 21292 9312 21312
rect 9312 21292 9364 21312
rect 9364 21292 9366 21312
rect 9310 21256 9366 21292
rect 9954 22636 10010 22672
rect 9954 22616 9956 22636
rect 9956 22616 10008 22636
rect 10008 22616 10010 22636
rect 9310 19624 9366 19680
rect 9402 19216 9458 19272
rect 9034 15136 9090 15192
rect 9218 15272 9274 15328
rect 9402 15544 9458 15600
rect 10046 17312 10102 17368
rect 9862 16904 9918 16960
rect 9770 16632 9826 16688
rect 9586 15136 9642 15192
rect 9770 15136 9826 15192
rect 9586 15000 9642 15056
rect 9218 12416 9274 12472
rect 9770 14048 9826 14104
rect 9402 12552 9458 12608
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 9126 9424 9182 9480
rect 9770 13368 9826 13424
rect 9402 9560 9458 9616
rect 10598 22092 10654 22128
rect 10598 22072 10600 22092
rect 10600 22072 10652 22092
rect 10652 22072 10654 22092
rect 10874 21392 10930 21448
rect 10782 20984 10838 21040
rect 10874 20712 10930 20768
rect 11150 24792 11206 24848
rect 11334 24656 11390 24712
rect 10414 18536 10470 18592
rect 10230 15580 10232 15600
rect 10232 15580 10284 15600
rect 10284 15580 10286 15600
rect 10230 15544 10286 15580
rect 10230 15444 10232 15464
rect 10232 15444 10284 15464
rect 10284 15444 10286 15464
rect 10230 15408 10286 15444
rect 10046 14184 10102 14240
rect 10874 18672 10930 18728
rect 10506 18400 10562 18456
rect 10598 16632 10654 16688
rect 10322 14592 10378 14648
rect 10322 14048 10378 14104
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 2870 1536 2926 1592
rect 10782 15136 10838 15192
rect 11978 22752 12034 22808
rect 11886 20440 11942 20496
rect 11426 19624 11482 19680
rect 11702 19216 11758 19272
rect 11610 17312 11666 17368
rect 11610 17040 11666 17096
rect 11150 15680 11206 15736
rect 11058 15136 11114 15192
rect 10782 12300 10838 12336
rect 10782 12280 10784 12300
rect 10784 12280 10836 12300
rect 10836 12280 10838 12300
rect 10782 11076 10838 11112
rect 11426 15408 11482 15464
rect 10782 11056 10784 11076
rect 10784 11056 10836 11076
rect 10836 11056 10838 11076
rect 10782 9596 10784 9616
rect 10784 9596 10836 9616
rect 10836 9596 10838 9616
rect 10782 9560 10838 9596
rect 11518 15036 11520 15056
rect 11520 15036 11572 15056
rect 11572 15036 11574 15056
rect 11518 15000 11574 15036
rect 11426 14864 11482 14920
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12530 24248 12586 24304
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12806 23160 12862 23216
rect 12530 22480 12586 22536
rect 12254 20460 12310 20496
rect 12254 20440 12256 20460
rect 12256 20440 12308 20460
rect 12308 20440 12310 20460
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12530 20324 12586 20360
rect 12530 20304 12532 20324
rect 12532 20304 12584 20324
rect 12584 20304 12586 20324
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12990 19760 13046 19816
rect 13542 21256 13598 21312
rect 12070 18128 12126 18184
rect 12070 17312 12126 17368
rect 12070 16088 12126 16144
rect 12438 18420 12494 18456
rect 12438 18400 12440 18420
rect 12440 18400 12492 18420
rect 12492 18400 12494 18420
rect 12346 17992 12402 18048
rect 12438 17448 12494 17504
rect 12254 15952 12310 16008
rect 11978 15020 12034 15056
rect 11978 15000 11980 15020
rect 11980 15000 12032 15020
rect 12032 15000 12034 15020
rect 10966 8200 11022 8256
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12714 18264 12770 18320
rect 12622 17992 12678 18048
rect 13358 18264 13414 18320
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13818 18808 13874 18864
rect 14830 24112 14886 24168
rect 13726 17720 13782 17776
rect 13726 17584 13782 17640
rect 13634 16904 13690 16960
rect 13450 16224 13506 16280
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12714 14184 12770 14240
rect 12714 13252 12770 13288
rect 12714 13232 12716 13252
rect 12716 13232 12768 13252
rect 12768 13232 12770 13252
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12622 12688 12678 12744
rect 12806 12688 12862 12744
rect 13450 14592 13506 14648
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12806 10104 12862 10160
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 13450 9988 13506 10024
rect 13450 9968 13452 9988
rect 13452 9968 13504 9988
rect 13504 9968 13506 9988
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 14370 20984 14426 21040
rect 15750 22752 15806 22808
rect 15014 19216 15070 19272
rect 15106 18264 15162 18320
rect 15290 17584 15346 17640
rect 15474 18400 15530 18456
rect 15014 17448 15070 17504
rect 14094 17040 14150 17096
rect 14186 16940 14188 16960
rect 14188 16940 14240 16960
rect 14240 16940 14242 16960
rect 14186 16904 14242 16940
rect 14186 16768 14242 16824
rect 14462 13640 14518 13696
rect 15106 15680 15162 15736
rect 15014 13252 15070 13288
rect 15014 13232 15016 13252
rect 15016 13232 15068 13252
rect 15068 13232 15070 13252
rect 15290 12008 15346 12064
rect 16578 23024 16634 23080
rect 15842 18536 15898 18592
rect 16118 17856 16174 17912
rect 15658 16768 15714 16824
rect 15658 15136 15714 15192
rect 16118 16496 16174 16552
rect 16302 14864 16358 14920
rect 16486 17992 16542 18048
rect 15290 9988 15346 10024
rect 15290 9968 15292 9988
rect 15292 9968 15344 9988
rect 15344 9968 15346 9988
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 16486 13232 16542 13288
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17406 21936 17462 21992
rect 17314 21256 17370 21312
rect 16946 20848 17002 20904
rect 16854 19352 16910 19408
rect 17130 17312 17186 17368
rect 16946 14320 17002 14376
rect 16578 10648 16634 10704
rect 16210 10104 16266 10160
rect 16118 9968 16174 10024
rect 17038 12008 17094 12064
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 19522 23840 19578 23896
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 18602 21664 18658 21720
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18418 20748 18420 20768
rect 18420 20748 18472 20768
rect 18472 20748 18474 20768
rect 18418 20712 18474 20748
rect 17866 19896 17922 19952
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17774 19080 17830 19136
rect 17498 18400 17554 18456
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18326 17992 18382 18048
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18602 19252 18604 19272
rect 18604 19252 18656 19272
rect 18656 19252 18658 19272
rect 18602 19216 18658 19252
rect 18602 18808 18658 18864
rect 18602 18400 18658 18456
rect 18602 17584 18658 17640
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17590 12008 17646 12064
rect 18970 19252 18972 19272
rect 18972 19252 19024 19272
rect 19024 19252 19026 19272
rect 18970 19216 19026 19252
rect 18970 19080 19026 19136
rect 18694 14592 18750 14648
rect 18602 12416 18658 12472
rect 19522 22228 19578 22264
rect 19522 22208 19524 22228
rect 19524 22208 19576 22228
rect 19576 22208 19578 22228
rect 19338 21836 19340 21856
rect 19340 21836 19392 21856
rect 19392 21836 19394 21856
rect 19338 21800 19394 21836
rect 19522 20576 19578 20632
rect 19522 19660 19524 19680
rect 19524 19660 19576 19680
rect 19576 19660 19578 19680
rect 19522 19624 19578 19660
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 19522 15952 19578 16008
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17866 9988 17922 10024
rect 17866 9968 17868 9988
rect 17868 9968 17920 9988
rect 17920 9968 17922 9988
rect 18418 9968 18474 10024
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 19062 12416 19118 12472
rect 19522 11056 19578 11112
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18970 9560 19026 9616
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 19890 23160 19946 23216
rect 19982 22228 20038 22264
rect 19982 22208 19984 22228
rect 19984 22208 20036 22228
rect 20036 22208 20038 22228
rect 20534 21800 20590 21856
rect 20074 21528 20130 21584
rect 20074 20712 20130 20768
rect 19890 17040 19946 17096
rect 19798 16496 19854 16552
rect 20350 17176 20406 17232
rect 20166 16632 20222 16688
rect 19982 13640 20038 13696
rect 20442 13368 20498 13424
rect 21270 18028 21272 18048
rect 21272 18028 21324 18048
rect 21324 18028 21326 18048
rect 21270 17992 21326 18028
rect 20994 17040 21050 17096
rect 20902 15816 20958 15872
rect 20902 14728 20958 14784
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22190 22208 22246 22264
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23202 21004 23258 21040
rect 23202 20984 23204 21004
rect 23204 20984 23256 21004
rect 23256 20984 23258 21004
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22650 19488 22706 19544
rect 22190 19352 22246 19408
rect 21730 17856 21786 17912
rect 21822 16496 21878 16552
rect 22190 17992 22246 18048
rect 22282 17720 22338 17776
rect 22282 17040 22338 17096
rect 20902 12824 20958 12880
rect 20442 12280 20498 12336
rect 22466 18808 22522 18864
rect 22466 18400 22522 18456
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22374 13504 22430 13560
rect 22650 15680 22706 15736
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 27158 24112 27214 24168
rect 23386 20984 23442 21040
rect 23386 20032 23442 20088
rect 23386 19624 23442 19680
rect 23662 21120 23718 21176
rect 23662 20748 23664 20768
rect 23664 20748 23716 20768
rect 23716 20748 23718 20768
rect 23662 20712 23718 20748
rect 23570 17584 23626 17640
rect 26238 23840 26294 23896
rect 28078 24656 28134 24712
rect 24950 21936 25006 21992
rect 25042 21800 25098 21856
rect 25042 21528 25098 21584
rect 25594 21412 25650 21448
rect 25594 21392 25596 21412
rect 25596 21392 25648 21412
rect 25648 21392 25650 21412
rect 25870 21664 25926 21720
rect 25594 20440 25650 20496
rect 25594 20168 25650 20224
rect 25226 20032 25282 20088
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23386 10512 23442 10568
rect 24858 18944 24914 19000
rect 24214 17176 24270 17232
rect 24490 17584 24546 17640
rect 25410 19216 25466 19272
rect 25134 16652 25190 16688
rect 25134 16632 25136 16652
rect 25136 16632 25188 16652
rect 25188 16632 25190 16652
rect 25226 16516 25282 16552
rect 25226 16496 25228 16516
rect 25228 16496 25280 16516
rect 25280 16496 25282 16516
rect 26238 19916 26294 19952
rect 26238 19896 26240 19916
rect 26240 19896 26292 19916
rect 26292 19896 26294 19916
rect 27526 22752 27582 22808
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 28262 23296 28318 23352
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27158 20712 27214 20768
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27894 21548 27950 21584
rect 27894 21528 27896 21548
rect 27896 21528 27948 21548
rect 27948 21528 27950 21548
rect 28814 23296 28870 23352
rect 25778 17176 25834 17232
rect 25134 14320 25190 14376
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 24858 8880 24914 8936
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 28538 20884 28540 20904
rect 28540 20884 28592 20904
rect 28592 20884 28594 20904
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27618 19488 27674 19544
rect 27434 18264 27490 18320
rect 28538 20848 28594 20884
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27618 18128 27674 18184
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27526 12144 27582 12200
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 28814 20712 28870 20768
rect 28998 20576 29054 20632
rect 29182 20440 29238 20496
rect 28998 20168 29054 20224
rect 29090 18808 29146 18864
rect 28814 17620 28816 17640
rect 28816 17620 28868 17640
rect 28868 17620 28870 17640
rect 28814 17584 28870 17620
rect 28722 16496 28778 16552
rect 28998 16088 29054 16144
rect 29550 20712 29606 20768
rect 29458 18944 29514 19000
rect 29826 19352 29882 19408
rect 29366 15544 29422 15600
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 30562 21120 30618 21176
rect 30286 20576 30342 20632
rect 31666 22072 31722 22128
rect 30286 17720 30342 17776
rect 29918 11192 29974 11248
rect 31298 9016 31354 9072
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 31942 23160 31998 23216
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 34610 24248 34666 24304
rect 32494 23568 32550 23624
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 33506 23024 33562 23080
rect 31482 15408 31538 15464
rect 32218 13912 32274 13968
rect 32310 13232 32366 13288
rect 32586 19760 32642 19816
rect 33230 22480 33286 22536
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32678 15000 32734 15056
rect 32402 11736 32458 11792
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 33506 20304 33562 20360
rect 33414 18672 33470 18728
rect 34242 22616 34298 22672
rect 34058 15952 34114 16008
rect 33322 13368 33378 13424
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 35162 24792 35218 24848
rect 35990 23740 35992 23760
rect 35992 23740 36044 23760
rect 36044 23740 36046 23760
rect 35990 23704 36046 23740
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 38658 20848 38714 20904
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 48318 24792 48374 24848
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 46938 21936 46994 21992
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 37186 16632 37242 16688
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 48686 21392 48742 21448
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 49054 23840 49110 23896
rect 49054 22888 49110 22944
rect 49054 21972 49056 21992
rect 49056 21972 49108 21992
rect 49108 21972 49110 21992
rect 49054 21936 49110 21972
rect 49146 20984 49202 21040
rect 48778 17176 48834 17232
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 34334 9424 34390 9480
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 0 25666 800 25696
rect 3325 25666 3391 25669
rect 0 25664 3391 25666
rect 0 25608 3330 25664
rect 3386 25608 3391 25664
rect 0 25606 3391 25608
rect 0 25576 800 25606
rect 3325 25603 3391 25606
rect 0 25258 800 25288
rect 3417 25258 3483 25261
rect 0 25256 3483 25258
rect 0 25200 3422 25256
rect 3478 25200 3483 25256
rect 0 25198 3483 25200
rect 0 25168 800 25198
rect 3417 25195 3483 25198
rect 0 24850 800 24880
rect 3877 24850 3943 24853
rect 0 24848 3943 24850
rect 0 24792 3882 24848
rect 3938 24792 3943 24848
rect 0 24790 3943 24792
rect 0 24760 800 24790
rect 3877 24787 3943 24790
rect 11145 24850 11211 24853
rect 35157 24850 35223 24853
rect 11145 24848 35223 24850
rect 11145 24792 11150 24848
rect 11206 24792 35162 24848
rect 35218 24792 35223 24848
rect 11145 24790 35223 24792
rect 11145 24787 11211 24790
rect 35157 24787 35223 24790
rect 48313 24850 48379 24853
rect 50200 24850 51000 24880
rect 48313 24848 51000 24850
rect 48313 24792 48318 24848
rect 48374 24792 51000 24848
rect 48313 24790 51000 24792
rect 48313 24787 48379 24790
rect 50200 24760 51000 24790
rect 11329 24714 11395 24717
rect 28073 24714 28139 24717
rect 11329 24712 28139 24714
rect 11329 24656 11334 24712
rect 11390 24656 28078 24712
rect 28134 24656 28139 24712
rect 11329 24654 28139 24656
rect 11329 24651 11395 24654
rect 28073 24651 28139 24654
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 1485 24442 1551 24445
rect 0 24440 1551 24442
rect 0 24384 1490 24440
rect 1546 24384 1551 24440
rect 0 24382 1551 24384
rect 0 24352 800 24382
rect 1485 24379 1551 24382
rect 12525 24306 12591 24309
rect 34605 24306 34671 24309
rect 12525 24304 34671 24306
rect 12525 24248 12530 24304
rect 12586 24248 34610 24304
rect 34666 24248 34671 24304
rect 12525 24246 34671 24248
rect 12525 24243 12591 24246
rect 34605 24243 34671 24246
rect 4797 24170 4863 24173
rect 9438 24170 9444 24172
rect 4797 24168 9444 24170
rect 4797 24112 4802 24168
rect 4858 24112 9444 24168
rect 4797 24110 9444 24112
rect 4797 24107 4863 24110
rect 9438 24108 9444 24110
rect 9508 24108 9514 24172
rect 14825 24170 14891 24173
rect 27153 24170 27219 24173
rect 14825 24168 27219 24170
rect 14825 24112 14830 24168
rect 14886 24112 27158 24168
rect 27214 24112 27219 24168
rect 14825 24110 27219 24112
rect 14825 24107 14891 24110
rect 27153 24107 27219 24110
rect 0 24034 800 24064
rect 3969 24034 4035 24037
rect 0 24032 4035 24034
rect 0 23976 3974 24032
rect 4030 23976 4035 24032
rect 0 23974 4035 23976
rect 0 23944 800 23974
rect 3969 23971 4035 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 19517 23898 19583 23901
rect 26233 23898 26299 23901
rect 19517 23896 26299 23898
rect 19517 23840 19522 23896
rect 19578 23840 26238 23896
rect 26294 23840 26299 23896
rect 19517 23838 26299 23840
rect 19517 23835 19583 23838
rect 26233 23835 26299 23838
rect 49049 23898 49115 23901
rect 50200 23898 51000 23928
rect 49049 23896 51000 23898
rect 49049 23840 49054 23896
rect 49110 23840 51000 23896
rect 49049 23838 51000 23840
rect 49049 23835 49115 23838
rect 50200 23808 51000 23838
rect 8109 23762 8175 23765
rect 35985 23762 36051 23765
rect 8109 23760 36051 23762
rect 8109 23704 8114 23760
rect 8170 23704 35990 23760
rect 36046 23704 36051 23760
rect 8109 23702 36051 23704
rect 8109 23699 8175 23702
rect 35985 23699 36051 23702
rect 0 23626 800 23656
rect 4061 23626 4127 23629
rect 0 23624 4127 23626
rect 0 23568 4066 23624
rect 4122 23568 4127 23624
rect 0 23566 4127 23568
rect 0 23536 800 23566
rect 4061 23563 4127 23566
rect 9949 23626 10015 23629
rect 32489 23626 32555 23629
rect 9949 23624 32555 23626
rect 9949 23568 9954 23624
rect 10010 23568 32494 23624
rect 32550 23568 32555 23624
rect 9949 23566 32555 23568
rect 9949 23563 10015 23566
rect 32489 23563 32555 23566
rect 3417 23490 3483 23493
rect 3918 23490 3924 23492
rect 3417 23488 3924 23490
rect 3417 23432 3422 23488
rect 3478 23432 3924 23488
rect 3417 23430 3924 23432
rect 3417 23427 3483 23430
rect 3918 23428 3924 23430
rect 3988 23428 3994 23492
rect 6637 23490 6703 23493
rect 11646 23490 11652 23492
rect 6637 23488 11652 23490
rect 6637 23432 6642 23488
rect 6698 23432 11652 23488
rect 6637 23430 11652 23432
rect 6637 23427 6703 23430
rect 11646 23428 11652 23430
rect 11716 23428 11722 23492
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 28257 23354 28323 23357
rect 28809 23354 28875 23357
rect 28257 23352 28875 23354
rect 28257 23296 28262 23352
rect 28318 23296 28814 23352
rect 28870 23296 28875 23352
rect 28257 23294 28875 23296
rect 28257 23291 28323 23294
rect 28809 23291 28875 23294
rect 0 23218 800 23248
rect 4981 23218 5047 23221
rect 0 23216 5047 23218
rect 0 23160 4986 23216
rect 5042 23160 5047 23216
rect 0 23158 5047 23160
rect 0 23128 800 23158
rect 4981 23155 5047 23158
rect 12801 23218 12867 23221
rect 19885 23218 19951 23221
rect 31937 23218 32003 23221
rect 12801 23216 18660 23218
rect 12801 23160 12806 23216
rect 12862 23160 18660 23216
rect 12801 23158 18660 23160
rect 12801 23155 12867 23158
rect 5390 23020 5396 23084
rect 5460 23082 5466 23084
rect 6821 23082 6887 23085
rect 5460 23080 6887 23082
rect 5460 23024 6826 23080
rect 6882 23024 6887 23080
rect 5460 23022 6887 23024
rect 5460 23020 5466 23022
rect 6821 23019 6887 23022
rect 16573 23082 16639 23085
rect 18600 23082 18660 23158
rect 19885 23216 32003 23218
rect 19885 23160 19890 23216
rect 19946 23160 31942 23216
rect 31998 23160 32003 23216
rect 19885 23158 32003 23160
rect 19885 23155 19951 23158
rect 31937 23155 32003 23158
rect 33501 23082 33567 23085
rect 16573 23080 18522 23082
rect 16573 23024 16578 23080
rect 16634 23024 18522 23080
rect 16573 23022 18522 23024
rect 18600 23080 33567 23082
rect 18600 23024 33506 23080
rect 33562 23024 33567 23080
rect 18600 23022 33567 23024
rect 16573 23019 16639 23022
rect 4889 22948 4955 22949
rect 4838 22946 4844 22948
rect 4798 22886 4844 22946
rect 4908 22944 4955 22948
rect 4950 22888 4955 22944
rect 4838 22884 4844 22886
rect 4908 22884 4955 22888
rect 18462 22946 18522 23022
rect 33501 23019 33567 23022
rect 49049 22946 49115 22949
rect 50200 22946 51000 22976
rect 18462 22886 22110 22946
rect 4889 22883 4955 22884
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 2497 22810 2563 22813
rect 0 22808 2563 22810
rect 0 22752 2502 22808
rect 2558 22752 2563 22808
rect 0 22750 2563 22752
rect 0 22720 800 22750
rect 2497 22747 2563 22750
rect 11973 22810 12039 22813
rect 15745 22810 15811 22813
rect 11973 22808 15811 22810
rect 11973 22752 11978 22808
rect 12034 22752 15750 22808
rect 15806 22752 15811 22808
rect 11973 22750 15811 22752
rect 22050 22810 22110 22886
rect 49049 22944 51000 22946
rect 49049 22888 49054 22944
rect 49110 22888 51000 22944
rect 49049 22886 51000 22888
rect 49049 22883 49115 22886
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 50200 22856 51000 22886
rect 47946 22815 48262 22816
rect 27521 22810 27587 22813
rect 22050 22808 27587 22810
rect 22050 22752 27526 22808
rect 27582 22752 27587 22808
rect 22050 22750 27587 22752
rect 11973 22747 12039 22750
rect 15745 22747 15811 22750
rect 27521 22747 27587 22750
rect 9949 22674 10015 22677
rect 34237 22674 34303 22677
rect 9949 22672 34303 22674
rect 9949 22616 9954 22672
rect 10010 22616 34242 22672
rect 34298 22616 34303 22672
rect 9949 22614 34303 22616
rect 9949 22611 10015 22614
rect 34237 22611 34303 22614
rect 3601 22538 3667 22541
rect 2270 22536 3667 22538
rect 2270 22480 3606 22536
rect 3662 22480 3667 22536
rect 2270 22478 3667 22480
rect 0 22402 800 22432
rect 2270 22402 2330 22478
rect 3601 22475 3667 22478
rect 12525 22538 12591 22541
rect 33225 22538 33291 22541
rect 12525 22536 33291 22538
rect 12525 22480 12530 22536
rect 12586 22480 33230 22536
rect 33286 22480 33291 22536
rect 12525 22478 33291 22480
rect 12525 22475 12591 22478
rect 33225 22475 33291 22478
rect 0 22342 2330 22402
rect 0 22312 800 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 3417 22266 3483 22269
rect 3550 22266 3556 22268
rect 3417 22264 3556 22266
rect 3417 22208 3422 22264
rect 3478 22208 3556 22264
rect 3417 22206 3556 22208
rect 3417 22203 3483 22206
rect 3550 22204 3556 22206
rect 3620 22204 3626 22268
rect 19517 22266 19583 22269
rect 19977 22266 20043 22269
rect 22185 22268 22251 22269
rect 22134 22266 22140 22268
rect 19517 22264 20043 22266
rect 19517 22208 19522 22264
rect 19578 22208 19982 22264
rect 20038 22208 20043 22264
rect 19517 22206 20043 22208
rect 22094 22206 22140 22266
rect 22204 22264 22251 22268
rect 22246 22208 22251 22264
rect 19517 22203 19583 22206
rect 19977 22203 20043 22206
rect 22134 22204 22140 22206
rect 22204 22204 22251 22208
rect 22185 22203 22251 22204
rect 3785 22130 3851 22133
rect 4061 22130 4127 22133
rect 3785 22128 4127 22130
rect 3785 22072 3790 22128
rect 3846 22072 4066 22128
rect 4122 22072 4127 22128
rect 3785 22070 4127 22072
rect 3785 22067 3851 22070
rect 4061 22067 4127 22070
rect 10593 22130 10659 22133
rect 31661 22130 31727 22133
rect 10593 22128 31727 22130
rect 10593 22072 10598 22128
rect 10654 22072 31666 22128
rect 31722 22072 31727 22128
rect 10593 22070 31727 22072
rect 10593 22067 10659 22070
rect 31661 22067 31727 22070
rect 0 21994 800 22024
rect 4429 21994 4495 21997
rect 7005 21996 7071 21997
rect 7005 21994 7052 21996
rect 0 21992 4495 21994
rect 0 21936 4434 21992
rect 4490 21936 4495 21992
rect 0 21934 4495 21936
rect 6960 21992 7052 21994
rect 6960 21936 7010 21992
rect 6960 21934 7052 21936
rect 0 21904 800 21934
rect 4429 21931 4495 21934
rect 7005 21932 7052 21934
rect 7116 21932 7122 21996
rect 17401 21994 17467 21997
rect 24945 21994 25011 21997
rect 46933 21994 46999 21997
rect 17401 21992 22110 21994
rect 17401 21936 17406 21992
rect 17462 21936 22110 21992
rect 17401 21934 22110 21936
rect 7005 21931 7071 21932
rect 17401 21931 17467 21934
rect 19333 21858 19399 21861
rect 20529 21858 20595 21861
rect 19333 21856 20595 21858
rect 19333 21800 19338 21856
rect 19394 21800 20534 21856
rect 20590 21800 20595 21856
rect 19333 21798 20595 21800
rect 22050 21858 22110 21934
rect 24945 21992 46999 21994
rect 24945 21936 24950 21992
rect 25006 21936 46938 21992
rect 46994 21936 46999 21992
rect 24945 21934 46999 21936
rect 24945 21931 25011 21934
rect 46933 21931 46999 21934
rect 49049 21994 49115 21997
rect 50200 21994 51000 22024
rect 49049 21992 51000 21994
rect 49049 21936 49054 21992
rect 49110 21936 51000 21992
rect 49049 21934 51000 21936
rect 49049 21931 49115 21934
rect 50200 21904 51000 21934
rect 25037 21858 25103 21861
rect 22050 21856 25103 21858
rect 22050 21800 25042 21856
rect 25098 21800 25103 21856
rect 22050 21798 25103 21800
rect 19333 21795 19399 21798
rect 20529 21795 20595 21798
rect 25037 21795 25103 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 3601 21722 3667 21725
rect 3734 21722 3740 21724
rect 3601 21720 3740 21722
rect 3601 21664 3606 21720
rect 3662 21664 3740 21720
rect 3601 21662 3740 21664
rect 3601 21659 3667 21662
rect 3734 21660 3740 21662
rect 3804 21660 3810 21724
rect 18597 21722 18663 21725
rect 25865 21722 25931 21725
rect 18597 21720 25931 21722
rect 18597 21664 18602 21720
rect 18658 21664 25870 21720
rect 25926 21664 25931 21720
rect 18597 21662 25931 21664
rect 18597 21659 18663 21662
rect 25865 21659 25931 21662
rect 0 21586 800 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 800 21526
rect 2681 21523 2747 21526
rect 6361 21586 6427 21589
rect 20069 21586 20135 21589
rect 6361 21584 20135 21586
rect 6361 21528 6366 21584
rect 6422 21528 20074 21584
rect 20130 21528 20135 21584
rect 6361 21526 20135 21528
rect 6361 21523 6427 21526
rect 20069 21523 20135 21526
rect 25037 21586 25103 21589
rect 27889 21586 27955 21589
rect 25037 21584 27955 21586
rect 25037 21528 25042 21584
rect 25098 21528 27894 21584
rect 27950 21528 27955 21584
rect 25037 21526 27955 21528
rect 25037 21523 25103 21526
rect 27889 21523 27955 21526
rect 6821 21450 6887 21453
rect 10869 21450 10935 21453
rect 6821 21448 10935 21450
rect 6821 21392 6826 21448
rect 6882 21392 10874 21448
rect 10930 21392 10935 21448
rect 6821 21390 10935 21392
rect 6821 21387 6887 21390
rect 10869 21387 10935 21390
rect 11646 21388 11652 21452
rect 11716 21450 11722 21452
rect 25589 21450 25655 21453
rect 11716 21448 25655 21450
rect 11716 21392 25594 21448
rect 25650 21392 25655 21448
rect 11716 21390 25655 21392
rect 11716 21388 11722 21390
rect 25589 21387 25655 21390
rect 27654 21388 27660 21452
rect 27724 21450 27730 21452
rect 48681 21450 48747 21453
rect 27724 21448 48747 21450
rect 27724 21392 48686 21448
rect 48742 21392 48747 21448
rect 27724 21390 48747 21392
rect 27724 21388 27730 21390
rect 48681 21387 48747 21390
rect 6177 21314 6243 21317
rect 9305 21314 9371 21317
rect 6177 21312 9371 21314
rect 6177 21256 6182 21312
rect 6238 21256 9310 21312
rect 9366 21256 9371 21312
rect 6177 21254 9371 21256
rect 6177 21251 6243 21254
rect 9305 21251 9371 21254
rect 13537 21314 13603 21317
rect 17309 21314 17375 21317
rect 13537 21312 17375 21314
rect 13537 21256 13542 21312
rect 13598 21256 17314 21312
rect 17370 21256 17375 21312
rect 13537 21254 17375 21256
rect 13537 21251 13603 21254
rect 17309 21251 17375 21254
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 23657 21178 23723 21181
rect 30557 21178 30623 21181
rect 23657 21176 30623 21178
rect 23657 21120 23662 21176
rect 23718 21120 30562 21176
rect 30618 21120 30623 21176
rect 23657 21118 30623 21120
rect 23657 21115 23723 21118
rect 30557 21115 30623 21118
rect 10777 21044 10843 21045
rect 10726 20980 10732 21044
rect 10796 21042 10843 21044
rect 14365 21042 14431 21045
rect 23197 21042 23263 21045
rect 10796 21040 10888 21042
rect 10838 20984 10888 21040
rect 10796 20982 10888 20984
rect 14365 21040 23263 21042
rect 14365 20984 14370 21040
rect 14426 20984 23202 21040
rect 23258 20984 23263 21040
rect 14365 20982 23263 20984
rect 10796 20980 10843 20982
rect 10777 20979 10843 20980
rect 14365 20979 14431 20982
rect 23197 20979 23263 20982
rect 23381 21042 23447 21045
rect 49141 21042 49207 21045
rect 50200 21042 51000 21072
rect 23381 21040 35910 21042
rect 23381 20984 23386 21040
rect 23442 20984 35910 21040
rect 23381 20982 35910 20984
rect 23381 20979 23447 20982
rect 16941 20906 17007 20909
rect 28533 20906 28599 20909
rect 16941 20904 28599 20906
rect 16941 20848 16946 20904
rect 17002 20848 28538 20904
rect 28594 20848 28599 20904
rect 16941 20846 28599 20848
rect 35850 20906 35910 20982
rect 49141 21040 51000 21042
rect 49141 20984 49146 21040
rect 49202 20984 51000 21040
rect 49141 20982 51000 20984
rect 49141 20979 49207 20982
rect 50200 20952 51000 20982
rect 38653 20906 38719 20909
rect 35850 20904 38719 20906
rect 35850 20848 38658 20904
rect 38714 20848 38719 20904
rect 35850 20846 38719 20848
rect 16941 20843 17007 20846
rect 28533 20843 28599 20846
rect 38653 20843 38719 20846
rect 0 20770 800 20800
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 800 20710
rect 1301 20707 1367 20710
rect 4153 20770 4219 20773
rect 4286 20770 4292 20772
rect 4153 20768 4292 20770
rect 4153 20712 4158 20768
rect 4214 20712 4292 20768
rect 4153 20710 4292 20712
rect 4153 20707 4219 20710
rect 4286 20708 4292 20710
rect 4356 20708 4362 20772
rect 7281 20770 7347 20773
rect 10869 20772 10935 20773
rect 7414 20770 7420 20772
rect 7281 20768 7420 20770
rect 7281 20712 7286 20768
rect 7342 20712 7420 20768
rect 7281 20710 7420 20712
rect 7281 20707 7347 20710
rect 7414 20708 7420 20710
rect 7484 20708 7490 20772
rect 10869 20770 10916 20772
rect 10824 20768 10916 20770
rect 10824 20712 10874 20768
rect 10824 20710 10916 20712
rect 10869 20708 10916 20710
rect 10980 20708 10986 20772
rect 18413 20770 18479 20773
rect 20069 20770 20135 20773
rect 18413 20768 20135 20770
rect 18413 20712 18418 20768
rect 18474 20712 20074 20768
rect 20130 20712 20135 20768
rect 18413 20710 20135 20712
rect 10869 20707 10935 20708
rect 18413 20707 18479 20710
rect 20069 20707 20135 20710
rect 23657 20770 23723 20773
rect 27153 20770 27219 20773
rect 23657 20768 27219 20770
rect 23657 20712 23662 20768
rect 23718 20712 27158 20768
rect 27214 20712 27219 20768
rect 23657 20710 27219 20712
rect 23657 20707 23723 20710
rect 27153 20707 27219 20710
rect 28809 20770 28875 20773
rect 29545 20770 29611 20773
rect 28809 20768 29611 20770
rect 28809 20712 28814 20768
rect 28870 20712 29550 20768
rect 29606 20712 29611 20768
rect 28809 20710 29611 20712
rect 28809 20707 28875 20710
rect 29545 20707 29611 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 6913 20634 6979 20637
rect 2730 20632 6979 20634
rect 2730 20576 6918 20632
rect 6974 20576 6979 20632
rect 2730 20574 6979 20576
rect 2589 20498 2655 20501
rect 2730 20498 2790 20574
rect 6913 20571 6979 20574
rect 19517 20634 19583 20637
rect 28993 20634 29059 20637
rect 30281 20634 30347 20637
rect 19517 20632 26802 20634
rect 19517 20576 19522 20632
rect 19578 20576 26802 20632
rect 19517 20574 26802 20576
rect 19517 20571 19583 20574
rect 2589 20496 2790 20498
rect 2589 20440 2594 20496
rect 2650 20440 2790 20496
rect 2589 20438 2790 20440
rect 6913 20498 6979 20501
rect 11881 20498 11947 20501
rect 6913 20496 11947 20498
rect 6913 20440 6918 20496
rect 6974 20440 11886 20496
rect 11942 20440 11947 20496
rect 6913 20438 11947 20440
rect 2589 20435 2655 20438
rect 6913 20435 6979 20438
rect 11881 20435 11947 20438
rect 12249 20498 12315 20501
rect 25589 20498 25655 20501
rect 12249 20496 25655 20498
rect 12249 20440 12254 20496
rect 12310 20440 25594 20496
rect 25650 20440 25655 20496
rect 12249 20438 25655 20440
rect 26742 20498 26802 20574
rect 28993 20632 30347 20634
rect 28993 20576 28998 20632
rect 29054 20576 30286 20632
rect 30342 20576 30347 20632
rect 28993 20574 30347 20576
rect 28993 20571 29059 20574
rect 30281 20571 30347 20574
rect 29177 20498 29243 20501
rect 26742 20496 29243 20498
rect 26742 20440 29182 20496
rect 29238 20440 29243 20496
rect 26742 20438 29243 20440
rect 12249 20435 12315 20438
rect 25589 20435 25655 20438
rect 29177 20435 29243 20438
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 12525 20362 12591 20365
rect 33501 20362 33567 20365
rect 12525 20360 33567 20362
rect 12525 20304 12530 20360
rect 12586 20304 33506 20360
rect 33562 20304 33567 20360
rect 12525 20302 33567 20304
rect 12525 20299 12591 20302
rect 33501 20299 33567 20302
rect 25589 20226 25655 20229
rect 28993 20226 29059 20229
rect 25589 20224 29059 20226
rect 25589 20168 25594 20224
rect 25650 20168 28998 20224
rect 29054 20168 29059 20224
rect 25589 20166 29059 20168
rect 25589 20163 25655 20166
rect 28993 20163 29059 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 23381 20090 23447 20093
rect 25221 20090 25287 20093
rect 23381 20088 25287 20090
rect 23381 20032 23386 20088
rect 23442 20032 25226 20088
rect 25282 20032 25287 20088
rect 23381 20030 25287 20032
rect 23381 20027 23447 20030
rect 25221 20027 25287 20030
rect 0 19954 800 19984
rect 2037 19954 2103 19957
rect 0 19952 2103 19954
rect 0 19896 2042 19952
rect 2098 19896 2103 19952
rect 0 19894 2103 19896
rect 0 19864 800 19894
rect 2037 19891 2103 19894
rect 17861 19954 17927 19957
rect 26233 19954 26299 19957
rect 17861 19952 26299 19954
rect 17861 19896 17866 19952
rect 17922 19896 26238 19952
rect 26294 19896 26299 19952
rect 17861 19894 26299 19896
rect 17861 19891 17927 19894
rect 26233 19891 26299 19894
rect 12985 19818 13051 19821
rect 32581 19818 32647 19821
rect 12985 19816 32647 19818
rect 12985 19760 12990 19816
rect 13046 19760 32586 19816
rect 32642 19760 32647 19816
rect 12985 19758 32647 19760
rect 12985 19755 13051 19758
rect 32581 19755 32647 19758
rect 9305 19682 9371 19685
rect 11094 19682 11100 19684
rect 9305 19680 11100 19682
rect 9305 19624 9310 19680
rect 9366 19624 11100 19680
rect 9305 19622 11100 19624
rect 9305 19619 9371 19622
rect 11094 19620 11100 19622
rect 11164 19682 11170 19684
rect 11421 19682 11487 19685
rect 11164 19680 11487 19682
rect 11164 19624 11426 19680
rect 11482 19624 11487 19680
rect 11164 19622 11487 19624
rect 11164 19620 11170 19622
rect 11421 19619 11487 19622
rect 19517 19682 19583 19685
rect 23381 19682 23447 19685
rect 19517 19680 23447 19682
rect 19517 19624 19522 19680
rect 19578 19624 23386 19680
rect 23442 19624 23447 19680
rect 19517 19622 23447 19624
rect 19517 19619 19583 19622
rect 23381 19619 23447 19622
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 2865 19546 2931 19549
rect 22645 19546 22711 19549
rect 27613 19546 27679 19549
rect 0 19544 2931 19546
rect 0 19488 2870 19544
rect 2926 19488 2931 19544
rect 0 19486 2931 19488
rect 0 19456 800 19486
rect 2865 19483 2931 19486
rect 22050 19486 22570 19546
rect 6126 19348 6132 19412
rect 6196 19410 6202 19412
rect 6637 19410 6703 19413
rect 6196 19408 6703 19410
rect 6196 19352 6642 19408
rect 6698 19352 6703 19408
rect 6196 19350 6703 19352
rect 6196 19348 6202 19350
rect 6637 19347 6703 19350
rect 16849 19410 16915 19413
rect 22050 19410 22110 19486
rect 16849 19408 22110 19410
rect 16849 19352 16854 19408
rect 16910 19352 22110 19408
rect 16849 19350 22110 19352
rect 22185 19410 22251 19413
rect 22318 19410 22324 19412
rect 22185 19408 22324 19410
rect 22185 19352 22190 19408
rect 22246 19352 22324 19408
rect 22185 19350 22324 19352
rect 16849 19347 16915 19350
rect 22185 19347 22251 19350
rect 22318 19348 22324 19350
rect 22388 19348 22394 19412
rect 22510 19410 22570 19486
rect 22645 19544 27679 19546
rect 22645 19488 22650 19544
rect 22706 19488 27618 19544
rect 27674 19488 27679 19544
rect 22645 19486 27679 19488
rect 22645 19483 22711 19486
rect 27613 19483 27679 19486
rect 29821 19410 29887 19413
rect 22510 19408 29887 19410
rect 22510 19352 29826 19408
rect 29882 19352 29887 19408
rect 22510 19350 29887 19352
rect 29821 19347 29887 19350
rect 1761 19274 1827 19277
rect 9397 19274 9463 19277
rect 1761 19272 9463 19274
rect 1761 19216 1766 19272
rect 1822 19216 9402 19272
rect 9458 19216 9463 19272
rect 1761 19214 9463 19216
rect 1761 19211 1827 19214
rect 9397 19211 9463 19214
rect 11697 19274 11763 19277
rect 15009 19274 15075 19277
rect 11697 19272 15075 19274
rect 11697 19216 11702 19272
rect 11758 19216 15014 19272
rect 15070 19216 15075 19272
rect 11697 19214 15075 19216
rect 11697 19211 11763 19214
rect 15009 19211 15075 19214
rect 18597 19274 18663 19277
rect 18965 19274 19031 19277
rect 18597 19272 19031 19274
rect 18597 19216 18602 19272
rect 18658 19216 18970 19272
rect 19026 19216 19031 19272
rect 18597 19214 19031 19216
rect 18597 19211 18663 19214
rect 18965 19211 19031 19214
rect 25405 19274 25471 19277
rect 27654 19274 27660 19276
rect 25405 19272 27660 19274
rect 25405 19216 25410 19272
rect 25466 19216 27660 19272
rect 25405 19214 27660 19216
rect 25405 19211 25471 19214
rect 27654 19212 27660 19214
rect 27724 19212 27730 19276
rect 0 19138 800 19168
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 800 19078
rect 2773 19075 2839 19078
rect 17769 19138 17835 19141
rect 18965 19138 19031 19141
rect 17769 19136 19031 19138
rect 17769 19080 17774 19136
rect 17830 19080 18970 19136
rect 19026 19080 19031 19136
rect 17769 19078 19031 19080
rect 17769 19075 17835 19078
rect 18965 19075 19031 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 24853 19002 24919 19005
rect 29453 19002 29519 19005
rect 24853 19000 29519 19002
rect 24853 18944 24858 19000
rect 24914 18944 29458 19000
rect 29514 18944 29519 19000
rect 24853 18942 29519 18944
rect 24853 18939 24919 18942
rect 29453 18939 29519 18942
rect 5809 18866 5875 18869
rect 8293 18866 8359 18869
rect 5809 18864 8359 18866
rect 5809 18808 5814 18864
rect 5870 18808 8298 18864
rect 8354 18808 8359 18864
rect 5809 18806 8359 18808
rect 5809 18803 5875 18806
rect 8293 18803 8359 18806
rect 13813 18866 13879 18869
rect 18597 18866 18663 18869
rect 13813 18864 18663 18866
rect 13813 18808 13818 18864
rect 13874 18808 18602 18864
rect 18658 18808 18663 18864
rect 13813 18806 18663 18808
rect 13813 18803 13879 18806
rect 18597 18803 18663 18806
rect 22461 18866 22527 18869
rect 29085 18866 29151 18869
rect 22461 18864 29151 18866
rect 22461 18808 22466 18864
rect 22522 18808 29090 18864
rect 29146 18808 29151 18864
rect 22461 18806 29151 18808
rect 22461 18803 22527 18806
rect 29085 18803 29151 18806
rect 0 18730 800 18760
rect 1393 18730 1459 18733
rect 0 18728 1459 18730
rect 0 18672 1398 18728
rect 1454 18672 1459 18728
rect 0 18670 1459 18672
rect 0 18640 800 18670
rect 1393 18667 1459 18670
rect 4889 18730 4955 18733
rect 7005 18730 7071 18733
rect 4889 18728 7071 18730
rect 4889 18672 4894 18728
rect 4950 18672 7010 18728
rect 7066 18672 7071 18728
rect 4889 18670 7071 18672
rect 4889 18667 4955 18670
rect 7005 18667 7071 18670
rect 10869 18730 10935 18733
rect 33409 18730 33475 18733
rect 10869 18728 33475 18730
rect 10869 18672 10874 18728
rect 10930 18672 33414 18728
rect 33470 18672 33475 18728
rect 10869 18670 33475 18672
rect 10869 18667 10935 18670
rect 33409 18667 33475 18670
rect 10409 18594 10475 18597
rect 15837 18594 15903 18597
rect 10409 18592 15903 18594
rect 10409 18536 10414 18592
rect 10470 18536 15842 18592
rect 15898 18536 15903 18592
rect 10409 18534 15903 18536
rect 10409 18531 10475 18534
rect 15837 18531 15903 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 47946 18463 48262 18464
rect 10501 18458 10567 18461
rect 12433 18458 12499 18461
rect 10501 18456 12499 18458
rect 10501 18400 10506 18456
rect 10562 18400 12438 18456
rect 12494 18400 12499 18456
rect 10501 18398 12499 18400
rect 10501 18395 10567 18398
rect 12433 18395 12499 18398
rect 15469 18458 15535 18461
rect 17493 18458 17559 18461
rect 15469 18456 17559 18458
rect 15469 18400 15474 18456
rect 15530 18400 17498 18456
rect 17554 18400 17559 18456
rect 15469 18398 17559 18400
rect 15469 18395 15535 18398
rect 17493 18395 17559 18398
rect 18597 18458 18663 18461
rect 22461 18458 22527 18461
rect 18597 18456 22527 18458
rect 18597 18400 18602 18456
rect 18658 18400 22466 18456
rect 22522 18400 22527 18456
rect 18597 18398 22527 18400
rect 18597 18395 18663 18398
rect 22461 18395 22527 18398
rect 0 18322 800 18352
rect 2037 18322 2103 18325
rect 0 18320 2103 18322
rect 0 18264 2042 18320
rect 2098 18264 2103 18320
rect 0 18262 2103 18264
rect 0 18232 800 18262
rect 2037 18259 2103 18262
rect 5625 18322 5691 18325
rect 8477 18322 8543 18325
rect 5625 18320 8543 18322
rect 5625 18264 5630 18320
rect 5686 18264 8482 18320
rect 8538 18264 8543 18320
rect 5625 18262 8543 18264
rect 5625 18259 5691 18262
rect 8477 18259 8543 18262
rect 12709 18322 12775 18325
rect 13353 18322 13419 18325
rect 12709 18320 13419 18322
rect 12709 18264 12714 18320
rect 12770 18264 13358 18320
rect 13414 18264 13419 18320
rect 12709 18262 13419 18264
rect 12709 18259 12775 18262
rect 13353 18259 13419 18262
rect 15101 18322 15167 18325
rect 27429 18322 27495 18325
rect 15101 18320 27495 18322
rect 15101 18264 15106 18320
rect 15162 18264 27434 18320
rect 27490 18264 27495 18320
rect 15101 18262 27495 18264
rect 15101 18259 15167 18262
rect 27429 18259 27495 18262
rect 12065 18186 12131 18189
rect 27613 18186 27679 18189
rect 12065 18184 27679 18186
rect 12065 18128 12070 18184
rect 12126 18128 27618 18184
rect 27674 18128 27679 18184
rect 12065 18126 27679 18128
rect 12065 18123 12131 18126
rect 27613 18123 27679 18126
rect 12341 18050 12407 18053
rect 12617 18050 12683 18053
rect 12341 18048 12683 18050
rect 12341 17992 12346 18048
rect 12402 17992 12622 18048
rect 12678 17992 12683 18048
rect 12341 17990 12683 17992
rect 12341 17987 12407 17990
rect 12617 17987 12683 17990
rect 16481 18050 16547 18053
rect 18321 18050 18387 18053
rect 16481 18048 18387 18050
rect 16481 17992 16486 18048
rect 16542 17992 18326 18048
rect 18382 17992 18387 18048
rect 16481 17990 18387 17992
rect 16481 17987 16547 17990
rect 18321 17987 18387 17990
rect 21265 18050 21331 18053
rect 22185 18050 22251 18053
rect 21265 18048 22251 18050
rect 21265 17992 21270 18048
rect 21326 17992 22190 18048
rect 22246 17992 22251 18048
rect 21265 17990 22251 17992
rect 21265 17987 21331 17990
rect 22185 17987 22251 17990
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 2497 17914 2563 17917
rect 0 17912 2563 17914
rect 0 17856 2502 17912
rect 2558 17856 2563 17912
rect 0 17854 2563 17856
rect 0 17824 800 17854
rect 2497 17851 2563 17854
rect 16113 17914 16179 17917
rect 21725 17914 21791 17917
rect 16113 17912 21791 17914
rect 16113 17856 16118 17912
rect 16174 17856 21730 17912
rect 21786 17856 21791 17912
rect 16113 17854 21791 17856
rect 16113 17851 16179 17854
rect 21725 17851 21791 17854
rect 2865 17778 2931 17781
rect 13721 17778 13787 17781
rect 2865 17776 13787 17778
rect 2865 17720 2870 17776
rect 2926 17720 13726 17776
rect 13782 17720 13787 17776
rect 2865 17718 13787 17720
rect 2865 17715 2931 17718
rect 13721 17715 13787 17718
rect 22277 17778 22343 17781
rect 30281 17778 30347 17781
rect 22277 17776 30347 17778
rect 22277 17720 22282 17776
rect 22338 17720 30286 17776
rect 30342 17720 30347 17776
rect 22277 17718 30347 17720
rect 22277 17715 22343 17718
rect 30281 17715 30347 17718
rect 1853 17642 1919 17645
rect 8017 17642 8083 17645
rect 1853 17640 8083 17642
rect 1853 17584 1858 17640
rect 1914 17584 8022 17640
rect 8078 17584 8083 17640
rect 1853 17582 8083 17584
rect 1853 17579 1919 17582
rect 8017 17579 8083 17582
rect 13721 17642 13787 17645
rect 15285 17642 15351 17645
rect 13721 17640 15351 17642
rect 13721 17584 13726 17640
rect 13782 17584 15290 17640
rect 15346 17584 15351 17640
rect 13721 17582 15351 17584
rect 13721 17579 13787 17582
rect 15285 17579 15351 17582
rect 18597 17642 18663 17645
rect 23565 17642 23631 17645
rect 24485 17642 24551 17645
rect 28809 17642 28875 17645
rect 18597 17640 28875 17642
rect 18597 17584 18602 17640
rect 18658 17584 23570 17640
rect 23626 17584 24490 17640
rect 24546 17584 28814 17640
rect 28870 17584 28875 17640
rect 18597 17582 28875 17584
rect 18597 17579 18663 17582
rect 23565 17579 23631 17582
rect 24485 17579 24551 17582
rect 28809 17579 28875 17582
rect 0 17506 800 17536
rect 2773 17506 2839 17509
rect 0 17504 2839 17506
rect 0 17448 2778 17504
rect 2834 17448 2839 17504
rect 0 17446 2839 17448
rect 0 17416 800 17446
rect 2773 17443 2839 17446
rect 12433 17506 12499 17509
rect 15009 17506 15075 17509
rect 12433 17504 15075 17506
rect 12433 17448 12438 17504
rect 12494 17448 15014 17504
rect 15070 17448 15075 17504
rect 12433 17446 15075 17448
rect 12433 17443 12499 17446
rect 15009 17443 15075 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 3877 17370 3943 17373
rect 5257 17370 5323 17373
rect 3877 17368 5323 17370
rect 3877 17312 3882 17368
rect 3938 17312 5262 17368
rect 5318 17312 5323 17368
rect 3877 17310 5323 17312
rect 3877 17307 3943 17310
rect 5257 17307 5323 17310
rect 10041 17370 10107 17373
rect 11605 17370 11671 17373
rect 10041 17368 11671 17370
rect 10041 17312 10046 17368
rect 10102 17312 11610 17368
rect 11666 17312 11671 17368
rect 10041 17310 11671 17312
rect 10041 17307 10107 17310
rect 11605 17307 11671 17310
rect 12065 17370 12131 17373
rect 17125 17370 17191 17373
rect 12065 17368 17191 17370
rect 12065 17312 12070 17368
rect 12126 17312 17130 17368
rect 17186 17312 17191 17368
rect 12065 17310 17191 17312
rect 12065 17307 12131 17310
rect 17125 17307 17191 17310
rect 4061 17234 4127 17237
rect 5349 17234 5415 17237
rect 4061 17232 5415 17234
rect 4061 17176 4066 17232
rect 4122 17176 5354 17232
rect 5410 17176 5415 17232
rect 4061 17174 5415 17176
rect 4061 17171 4127 17174
rect 5349 17171 5415 17174
rect 8477 17234 8543 17237
rect 20345 17234 20411 17237
rect 24209 17234 24275 17237
rect 8477 17232 24275 17234
rect 8477 17176 8482 17232
rect 8538 17176 20350 17232
rect 20406 17176 24214 17232
rect 24270 17176 24275 17232
rect 8477 17174 24275 17176
rect 8477 17171 8543 17174
rect 20345 17171 20411 17174
rect 24209 17171 24275 17174
rect 25773 17234 25839 17237
rect 48773 17234 48839 17237
rect 25773 17232 48839 17234
rect 25773 17176 25778 17232
rect 25834 17176 48778 17232
rect 48834 17176 48839 17232
rect 25773 17174 48839 17176
rect 25773 17171 25839 17174
rect 48773 17171 48839 17174
rect 0 17098 800 17128
rect 1209 17098 1275 17101
rect 0 17096 1275 17098
rect 0 17040 1214 17096
rect 1270 17040 1275 17096
rect 0 17038 1275 17040
rect 0 17008 800 17038
rect 1209 17035 1275 17038
rect 3734 17036 3740 17100
rect 3804 17098 3810 17100
rect 5349 17098 5415 17101
rect 11605 17098 11671 17101
rect 3804 17096 11671 17098
rect 3804 17040 5354 17096
rect 5410 17040 11610 17096
rect 11666 17040 11671 17096
rect 3804 17038 11671 17040
rect 3804 17036 3810 17038
rect 5349 17035 5415 17038
rect 11605 17035 11671 17038
rect 14089 17098 14155 17101
rect 19885 17098 19951 17101
rect 14089 17096 19951 17098
rect 14089 17040 14094 17096
rect 14150 17040 19890 17096
rect 19946 17040 19951 17096
rect 14089 17038 19951 17040
rect 14089 17035 14155 17038
rect 19885 17035 19951 17038
rect 20989 17098 21055 17101
rect 22277 17098 22343 17101
rect 20989 17096 22343 17098
rect 20989 17040 20994 17096
rect 21050 17040 22282 17096
rect 22338 17040 22343 17096
rect 20989 17038 22343 17040
rect 20989 17035 21055 17038
rect 22277 17035 22343 17038
rect 3325 16962 3391 16965
rect 9857 16962 9923 16965
rect 3325 16960 9923 16962
rect 3325 16904 3330 16960
rect 3386 16904 9862 16960
rect 9918 16904 9923 16960
rect 3325 16902 9923 16904
rect 3325 16899 3391 16902
rect 9857 16899 9923 16902
rect 13629 16962 13695 16965
rect 14181 16962 14247 16965
rect 13629 16960 14247 16962
rect 13629 16904 13634 16960
rect 13690 16904 14186 16960
rect 14242 16904 14247 16960
rect 13629 16902 14247 16904
rect 13629 16899 13695 16902
rect 14181 16899 14247 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 14181 16826 14247 16829
rect 15653 16826 15719 16829
rect 14181 16824 15719 16826
rect 14181 16768 14186 16824
rect 14242 16768 15658 16824
rect 15714 16768 15719 16824
rect 14181 16766 15719 16768
rect 14181 16763 14247 16766
rect 15653 16763 15719 16766
rect 0 16690 800 16720
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 800 16630
rect 1301 16627 1367 16630
rect 5349 16690 5415 16693
rect 9765 16690 9831 16693
rect 10593 16690 10659 16693
rect 20161 16690 20227 16693
rect 5349 16688 20227 16690
rect 5349 16632 5354 16688
rect 5410 16632 9770 16688
rect 9826 16632 10598 16688
rect 10654 16632 20166 16688
rect 20222 16632 20227 16688
rect 5349 16630 20227 16632
rect 5349 16627 5415 16630
rect 9765 16627 9831 16630
rect 10593 16627 10659 16630
rect 20161 16627 20227 16630
rect 25129 16690 25195 16693
rect 37181 16690 37247 16693
rect 25129 16688 37247 16690
rect 25129 16632 25134 16688
rect 25190 16632 37186 16688
rect 37242 16632 37247 16688
rect 25129 16630 37247 16632
rect 25129 16627 25195 16630
rect 37181 16627 37247 16630
rect 3918 16492 3924 16556
rect 3988 16554 3994 16556
rect 4337 16554 4403 16557
rect 3988 16552 4403 16554
rect 3988 16496 4342 16552
rect 4398 16496 4403 16552
rect 3988 16494 4403 16496
rect 3988 16492 3994 16494
rect 4337 16491 4403 16494
rect 8201 16554 8267 16557
rect 16113 16554 16179 16557
rect 19793 16554 19859 16557
rect 8201 16552 16179 16554
rect 8201 16496 8206 16552
rect 8262 16496 16118 16552
rect 16174 16496 16179 16552
rect 8201 16494 16179 16496
rect 8201 16491 8267 16494
rect 16113 16491 16179 16494
rect 17726 16552 19859 16554
rect 17726 16496 19798 16552
rect 19854 16496 19859 16552
rect 17726 16494 19859 16496
rect 17726 16418 17786 16494
rect 19793 16491 19859 16494
rect 21817 16554 21883 16557
rect 25221 16554 25287 16557
rect 28717 16554 28783 16557
rect 21817 16552 28783 16554
rect 21817 16496 21822 16552
rect 21878 16496 25226 16552
rect 25282 16496 28722 16552
rect 28778 16496 28783 16552
rect 21817 16494 28783 16496
rect 21817 16491 21883 16494
rect 25221 16491 25287 16494
rect 28717 16491 28783 16494
rect 11470 16358 17786 16418
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 7097 16146 7163 16149
rect 11470 16146 11530 16358
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 13445 16282 13511 16285
rect 7097 16144 11530 16146
rect 7097 16088 7102 16144
rect 7158 16088 11530 16144
rect 7097 16086 11530 16088
rect 11654 16280 13511 16282
rect 11654 16224 13450 16280
rect 13506 16224 13511 16280
rect 11654 16222 13511 16224
rect 7097 16083 7163 16086
rect 4889 16010 4955 16013
rect 11654 16010 11714 16222
rect 13445 16219 13511 16222
rect 12065 16146 12131 16149
rect 28993 16146 29059 16149
rect 12065 16144 29059 16146
rect 12065 16088 12070 16144
rect 12126 16088 28998 16144
rect 29054 16088 29059 16144
rect 12065 16086 29059 16088
rect 12065 16083 12131 16086
rect 28993 16083 29059 16086
rect 4889 16008 11714 16010
rect 4889 15952 4894 16008
rect 4950 15952 11714 16008
rect 4889 15950 11714 15952
rect 12249 16010 12315 16013
rect 19517 16010 19583 16013
rect 34053 16010 34119 16013
rect 12249 16008 16682 16010
rect 12249 15952 12254 16008
rect 12310 15952 16682 16008
rect 12249 15950 16682 15952
rect 4889 15947 4955 15950
rect 12249 15947 12315 15950
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 4153 15874 4219 15877
rect 8385 15874 8451 15877
rect 4153 15872 8451 15874
rect 4153 15816 4158 15872
rect 4214 15816 8390 15872
rect 8446 15816 8451 15872
rect 4153 15814 8451 15816
rect 16622 15874 16682 15950
rect 19517 16008 34119 16010
rect 19517 15952 19522 16008
rect 19578 15952 34058 16008
rect 34114 15952 34119 16008
rect 19517 15950 34119 15952
rect 19517 15947 19583 15950
rect 34053 15947 34119 15950
rect 20897 15874 20963 15877
rect 16622 15872 20963 15874
rect 16622 15816 20902 15872
rect 20958 15816 20963 15872
rect 16622 15814 20963 15816
rect 4153 15811 4219 15814
rect 8385 15811 8451 15814
rect 20897 15811 20963 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 5073 15738 5139 15741
rect 8201 15738 8267 15741
rect 11145 15740 11211 15741
rect 5073 15736 8267 15738
rect 5073 15680 5078 15736
rect 5134 15680 8206 15736
rect 8262 15680 8267 15736
rect 5073 15678 8267 15680
rect 5073 15675 5139 15678
rect 8201 15675 8267 15678
rect 11094 15676 11100 15740
rect 11164 15738 11211 15740
rect 15101 15738 15167 15741
rect 22645 15738 22711 15741
rect 11164 15736 11256 15738
rect 11206 15680 11256 15736
rect 11164 15678 11256 15680
rect 15101 15736 22711 15738
rect 15101 15680 15106 15736
rect 15162 15680 22650 15736
rect 22706 15680 22711 15736
rect 15101 15678 22711 15680
rect 11164 15676 11211 15678
rect 11145 15675 11211 15676
rect 15101 15675 15167 15678
rect 22645 15675 22711 15678
rect 4705 15602 4771 15605
rect 7373 15602 7439 15605
rect 4705 15600 7439 15602
rect 4705 15544 4710 15600
rect 4766 15544 7378 15600
rect 7434 15544 7439 15600
rect 4705 15542 7439 15544
rect 4705 15539 4771 15542
rect 7373 15539 7439 15542
rect 7557 15602 7623 15605
rect 9397 15602 9463 15605
rect 7557 15600 9463 15602
rect 7557 15544 7562 15600
rect 7618 15544 9402 15600
rect 9458 15544 9463 15600
rect 7557 15542 9463 15544
rect 7557 15539 7623 15542
rect 9397 15539 9463 15542
rect 10225 15602 10291 15605
rect 29361 15602 29427 15605
rect 10225 15600 29427 15602
rect 10225 15544 10230 15600
rect 10286 15544 29366 15600
rect 29422 15544 29427 15600
rect 10225 15542 29427 15544
rect 10225 15539 10291 15542
rect 29361 15539 29427 15542
rect 0 15466 800 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 800 15406
rect 1301 15403 1367 15406
rect 6637 15466 6703 15469
rect 7097 15466 7163 15469
rect 6637 15464 7163 15466
rect 6637 15408 6642 15464
rect 6698 15408 7102 15464
rect 7158 15408 7163 15464
rect 6637 15406 7163 15408
rect 6637 15403 6703 15406
rect 7097 15403 7163 15406
rect 7741 15466 7807 15469
rect 9990 15466 9996 15468
rect 7741 15464 9996 15466
rect 7741 15408 7746 15464
rect 7802 15408 9996 15464
rect 7741 15406 9996 15408
rect 7741 15403 7807 15406
rect 9990 15404 9996 15406
rect 10060 15404 10066 15468
rect 10225 15466 10291 15469
rect 11421 15466 11487 15469
rect 31477 15466 31543 15469
rect 10225 15464 11487 15466
rect 10225 15408 10230 15464
rect 10286 15408 11426 15464
rect 11482 15408 11487 15464
rect 10225 15406 11487 15408
rect 10225 15403 10291 15406
rect 11421 15403 11487 15406
rect 12390 15464 31543 15466
rect 12390 15408 31482 15464
rect 31538 15408 31543 15464
rect 12390 15406 31543 15408
rect 3550 15268 3556 15332
rect 3620 15330 3626 15332
rect 4429 15330 4495 15333
rect 3620 15328 4495 15330
rect 3620 15272 4434 15328
rect 4490 15272 4495 15328
rect 3620 15270 4495 15272
rect 3620 15268 3626 15270
rect 4429 15267 4495 15270
rect 9213 15330 9279 15333
rect 12390 15330 12450 15406
rect 31477 15403 31543 15406
rect 9213 15328 12450 15330
rect 9213 15272 9218 15328
rect 9274 15272 12450 15328
rect 9213 15270 12450 15272
rect 9213 15267 9279 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 9029 15194 9095 15197
rect 9581 15194 9647 15197
rect 9029 15192 9647 15194
rect 9029 15136 9034 15192
rect 9090 15136 9586 15192
rect 9642 15136 9647 15192
rect 9029 15134 9647 15136
rect 9029 15131 9095 15134
rect 9581 15131 9647 15134
rect 9765 15192 9831 15197
rect 9765 15136 9770 15192
rect 9826 15136 9831 15192
rect 9765 15131 9831 15136
rect 10777 15194 10843 15197
rect 10910 15194 10916 15196
rect 10777 15192 10916 15194
rect 10777 15136 10782 15192
rect 10838 15136 10916 15192
rect 10777 15134 10916 15136
rect 10777 15131 10843 15134
rect 10910 15132 10916 15134
rect 10980 15132 10986 15196
rect 11053 15194 11119 15197
rect 15653 15194 15719 15197
rect 11053 15192 15719 15194
rect 11053 15136 11058 15192
rect 11114 15136 15658 15192
rect 15714 15136 15719 15192
rect 11053 15134 15719 15136
rect 11053 15131 11119 15134
rect 15653 15131 15719 15134
rect 0 15058 800 15088
rect 1301 15058 1367 15061
rect 0 15056 1367 15058
rect 0 15000 1306 15056
rect 1362 15000 1367 15056
rect 0 14998 1367 15000
rect 0 14968 800 14998
rect 1301 14995 1367 14998
rect 7741 15058 7807 15061
rect 9581 15058 9647 15061
rect 7741 15056 9647 15058
rect 7741 15000 7746 15056
rect 7802 15000 9586 15056
rect 9642 15000 9647 15056
rect 7741 14998 9647 15000
rect 9768 15058 9828 15131
rect 11513 15058 11579 15061
rect 9768 15056 11579 15058
rect 9768 15000 11518 15056
rect 11574 15000 11579 15056
rect 9768 14998 11579 15000
rect 7741 14995 7807 14998
rect 9581 14995 9647 14998
rect 11513 14995 11579 14998
rect 11973 15058 12039 15061
rect 32673 15058 32739 15061
rect 11973 15056 32739 15058
rect 11973 15000 11978 15056
rect 12034 15000 32678 15056
rect 32734 15000 32739 15056
rect 11973 14998 32739 15000
rect 11973 14995 12039 14998
rect 32673 14995 32739 14998
rect 7598 14860 7604 14924
rect 7668 14922 7674 14924
rect 11421 14922 11487 14925
rect 16297 14922 16363 14925
rect 7668 14920 16363 14922
rect 7668 14864 11426 14920
rect 11482 14864 16302 14920
rect 16358 14864 16363 14920
rect 7668 14862 16363 14864
rect 7668 14860 7674 14862
rect 11421 14859 11487 14862
rect 16297 14859 16363 14862
rect 20897 14786 20963 14789
rect 22318 14786 22324 14788
rect 20897 14784 22324 14786
rect 20897 14728 20902 14784
rect 20958 14728 22324 14784
rect 20897 14726 22324 14728
rect 20897 14723 20963 14726
rect 22318 14724 22324 14726
rect 22388 14724 22394 14788
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 1301 14650 1367 14653
rect 10317 14650 10383 14653
rect 0 14648 1367 14650
rect 0 14592 1306 14648
rect 1362 14592 1367 14648
rect 0 14590 1367 14592
rect 0 14560 800 14590
rect 1301 14587 1367 14590
rect 10182 14648 10383 14650
rect 10182 14592 10322 14648
rect 10378 14592 10383 14648
rect 10182 14590 10383 14592
rect 1853 14514 1919 14517
rect 10182 14514 10242 14590
rect 10317 14587 10383 14590
rect 13445 14650 13511 14653
rect 18689 14650 18755 14653
rect 13445 14648 18755 14650
rect 13445 14592 13450 14648
rect 13506 14592 18694 14648
rect 18750 14592 18755 14648
rect 13445 14590 18755 14592
rect 13445 14587 13511 14590
rect 18689 14587 18755 14590
rect 1853 14512 10242 14514
rect 1853 14456 1858 14512
rect 1914 14456 10242 14512
rect 1853 14454 10242 14456
rect 1853 14451 1919 14454
rect 9990 14316 9996 14380
rect 10060 14378 10066 14380
rect 16941 14378 17007 14381
rect 25129 14378 25195 14381
rect 10060 14376 25195 14378
rect 10060 14320 16946 14376
rect 17002 14320 25134 14376
rect 25190 14320 25195 14376
rect 10060 14318 25195 14320
rect 10060 14316 10066 14318
rect 16941 14315 17007 14318
rect 25129 14315 25195 14318
rect 0 14242 800 14272
rect 2773 14242 2839 14245
rect 0 14240 2839 14242
rect 0 14184 2778 14240
rect 2834 14184 2839 14240
rect 0 14182 2839 14184
rect 0 14152 800 14182
rect 2773 14179 2839 14182
rect 10041 14242 10107 14245
rect 12709 14242 12775 14245
rect 10041 14240 12775 14242
rect 10041 14184 10046 14240
rect 10102 14184 12714 14240
rect 12770 14184 12775 14240
rect 10041 14182 12775 14184
rect 10041 14179 10107 14182
rect 12709 14179 12775 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 9765 14106 9831 14109
rect 10317 14106 10383 14109
rect 9765 14104 10383 14106
rect 9765 14048 9770 14104
rect 9826 14048 10322 14104
rect 10378 14048 10383 14104
rect 9765 14046 10383 14048
rect 9765 14043 9831 14046
rect 10317 14043 10383 14046
rect 3693 13970 3759 13973
rect 32213 13970 32279 13973
rect 3693 13968 32279 13970
rect 3693 13912 3698 13968
rect 3754 13912 32218 13968
rect 32274 13912 32279 13968
rect 3693 13910 32279 13912
rect 3693 13907 3759 13910
rect 32213 13907 32279 13910
rect 0 13834 800 13864
rect 2681 13834 2747 13837
rect 0 13832 2747 13834
rect 0 13776 2686 13832
rect 2742 13776 2747 13832
rect 0 13774 2747 13776
rect 0 13744 800 13774
rect 2681 13771 2747 13774
rect 6729 13698 6795 13701
rect 8293 13698 8359 13701
rect 6729 13696 8359 13698
rect 6729 13640 6734 13696
rect 6790 13640 8298 13696
rect 8354 13640 8359 13696
rect 6729 13638 8359 13640
rect 6729 13635 6795 13638
rect 8293 13635 8359 13638
rect 14457 13698 14523 13701
rect 19977 13698 20043 13701
rect 14457 13696 20043 13698
rect 14457 13640 14462 13696
rect 14518 13640 19982 13696
rect 20038 13640 20043 13696
rect 14457 13638 20043 13640
rect 14457 13635 14523 13638
rect 19977 13635 20043 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 22369 13562 22435 13565
rect 19290 13560 22435 13562
rect 19290 13504 22374 13560
rect 22430 13504 22435 13560
rect 19290 13502 22435 13504
rect 0 13426 800 13456
rect 1577 13426 1643 13429
rect 0 13424 1643 13426
rect 0 13368 1582 13424
rect 1638 13368 1643 13424
rect 0 13366 1643 13368
rect 0 13336 800 13366
rect 1577 13363 1643 13366
rect 9765 13426 9831 13429
rect 19290 13426 19350 13502
rect 22369 13499 22435 13502
rect 9765 13424 19350 13426
rect 9765 13368 9770 13424
rect 9826 13368 19350 13424
rect 9765 13366 19350 13368
rect 20437 13426 20503 13429
rect 33317 13426 33383 13429
rect 20437 13424 33383 13426
rect 20437 13368 20442 13424
rect 20498 13368 33322 13424
rect 33378 13368 33383 13424
rect 20437 13366 33383 13368
rect 9765 13363 9831 13366
rect 20437 13363 20503 13366
rect 33317 13363 33383 13366
rect 12709 13290 12775 13293
rect 15009 13290 15075 13293
rect 12709 13288 15075 13290
rect 12709 13232 12714 13288
rect 12770 13232 15014 13288
rect 15070 13232 15075 13288
rect 12709 13230 15075 13232
rect 12709 13227 12775 13230
rect 15009 13227 15075 13230
rect 16481 13290 16547 13293
rect 32305 13290 32371 13293
rect 16481 13288 32371 13290
rect 16481 13232 16486 13288
rect 16542 13232 32310 13288
rect 32366 13232 32371 13288
rect 16481 13230 32371 13232
rect 16481 13227 16547 13230
rect 32305 13227 32371 13230
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 3325 13018 3391 13021
rect 0 13016 3391 13018
rect 0 12960 3330 13016
rect 3386 12960 3391 13016
rect 0 12958 3391 12960
rect 0 12928 800 12958
rect 3325 12955 3391 12958
rect 1761 12882 1827 12885
rect 20897 12882 20963 12885
rect 1761 12880 20963 12882
rect 1761 12824 1766 12880
rect 1822 12824 20902 12880
rect 20958 12824 20963 12880
rect 1761 12822 20963 12824
rect 1761 12819 1827 12822
rect 20897 12819 20963 12822
rect 12617 12746 12683 12749
rect 12801 12746 12867 12749
rect 12617 12744 12867 12746
rect 12617 12688 12622 12744
rect 12678 12688 12806 12744
rect 12862 12688 12867 12744
rect 12617 12686 12867 12688
rect 12617 12683 12683 12686
rect 12801 12683 12867 12686
rect 0 12610 800 12640
rect 1761 12610 1827 12613
rect 0 12608 1827 12610
rect 0 12552 1766 12608
rect 1822 12552 1827 12608
rect 0 12550 1827 12552
rect 0 12520 800 12550
rect 1761 12547 1827 12550
rect 4705 12610 4771 12613
rect 9397 12610 9463 12613
rect 4705 12608 9463 12610
rect 4705 12552 4710 12608
rect 4766 12552 9402 12608
rect 9458 12552 9463 12608
rect 4705 12550 9463 12552
rect 4705 12547 4771 12550
rect 9397 12547 9463 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 9213 12474 9279 12477
rect 4478 12472 9279 12474
rect 4478 12416 9218 12472
rect 9274 12416 9279 12472
rect 4478 12414 9279 12416
rect 4478 12341 4538 12414
rect 9213 12411 9279 12414
rect 18597 12474 18663 12477
rect 19057 12474 19123 12477
rect 18597 12472 19123 12474
rect 18597 12416 18602 12472
rect 18658 12416 19062 12472
rect 19118 12416 19123 12472
rect 18597 12414 19123 12416
rect 18597 12411 18663 12414
rect 19057 12411 19123 12414
rect 4429 12336 4538 12341
rect 4429 12280 4434 12336
rect 4490 12280 4538 12336
rect 4429 12278 4538 12280
rect 7465 12338 7531 12341
rect 7598 12338 7604 12340
rect 7465 12336 7604 12338
rect 7465 12280 7470 12336
rect 7526 12280 7604 12336
rect 7465 12278 7604 12280
rect 4429 12275 4495 12278
rect 7465 12275 7531 12278
rect 7598 12276 7604 12278
rect 7668 12276 7674 12340
rect 10777 12338 10843 12341
rect 20437 12338 20503 12341
rect 10777 12336 20503 12338
rect 10777 12280 10782 12336
rect 10838 12280 20442 12336
rect 20498 12280 20503 12336
rect 10777 12278 20503 12280
rect 10777 12275 10843 12278
rect 20437 12275 20503 12278
rect 0 12202 800 12232
rect 2773 12202 2839 12205
rect 27521 12202 27587 12205
rect 0 12142 1594 12202
rect 0 12112 800 12142
rect 1534 12066 1594 12142
rect 2773 12200 27587 12202
rect 2773 12144 2778 12200
rect 2834 12144 27526 12200
rect 27582 12144 27587 12200
rect 2773 12142 27587 12144
rect 2773 12139 2839 12142
rect 27521 12139 27587 12142
rect 2865 12066 2931 12069
rect 1534 12064 2931 12066
rect 1534 12008 2870 12064
rect 2926 12008 2931 12064
rect 1534 12006 2931 12008
rect 2865 12003 2931 12006
rect 15285 12066 15351 12069
rect 17033 12066 17099 12069
rect 17585 12066 17651 12069
rect 15285 12064 17651 12066
rect 15285 12008 15290 12064
rect 15346 12008 17038 12064
rect 17094 12008 17590 12064
rect 17646 12008 17651 12064
rect 15285 12006 17651 12008
rect 15285 12003 15351 12006
rect 17033 12003 17099 12006
rect 17585 12003 17651 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 0 11794 800 11824
rect 3417 11794 3483 11797
rect 0 11792 3483 11794
rect 0 11736 3422 11792
rect 3478 11736 3483 11792
rect 0 11734 3483 11736
rect 0 11704 800 11734
rect 3417 11731 3483 11734
rect 5441 11794 5507 11797
rect 32397 11794 32463 11797
rect 5441 11792 32463 11794
rect 5441 11736 5446 11792
rect 5502 11736 32402 11792
rect 32458 11736 32463 11792
rect 5441 11734 32463 11736
rect 5441 11731 5507 11734
rect 32397 11731 32463 11734
rect 7281 11658 7347 11661
rect 22134 11658 22140 11660
rect 7281 11656 22140 11658
rect 7281 11600 7286 11656
rect 7342 11600 22140 11656
rect 7281 11598 22140 11600
rect 7281 11595 7347 11598
rect 22134 11596 22140 11598
rect 22204 11596 22210 11660
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 4705 11386 4771 11389
rect 5390 11386 5396 11388
rect 0 11326 1594 11386
rect 0 11296 800 11326
rect 1534 11114 1594 11326
rect 4705 11384 5396 11386
rect 4705 11328 4710 11384
rect 4766 11328 5396 11384
rect 4705 11326 5396 11328
rect 4705 11323 4771 11326
rect 5390 11324 5396 11326
rect 5460 11324 5466 11388
rect 2773 11250 2839 11253
rect 29913 11250 29979 11253
rect 2773 11248 29979 11250
rect 2773 11192 2778 11248
rect 2834 11192 29918 11248
rect 29974 11192 29979 11248
rect 2773 11190 29979 11192
rect 2773 11187 2839 11190
rect 29913 11187 29979 11190
rect 3509 11114 3575 11117
rect 1534 11112 3575 11114
rect 1534 11056 3514 11112
rect 3570 11056 3575 11112
rect 1534 11054 3575 11056
rect 3509 11051 3575 11054
rect 4838 11052 4844 11116
rect 4908 11114 4914 11116
rect 5165 11114 5231 11117
rect 7097 11116 7163 11117
rect 7046 11114 7052 11116
rect 4908 11112 5231 11114
rect 4908 11056 5170 11112
rect 5226 11056 5231 11112
rect 4908 11054 5231 11056
rect 7006 11054 7052 11114
rect 7116 11112 7163 11116
rect 7158 11056 7163 11112
rect 4908 11052 4914 11054
rect 5165 11051 5231 11054
rect 7046 11052 7052 11054
rect 7116 11052 7163 11056
rect 7414 11052 7420 11116
rect 7484 11114 7490 11116
rect 7741 11114 7807 11117
rect 7484 11112 7807 11114
rect 7484 11056 7746 11112
rect 7802 11056 7807 11112
rect 7484 11054 7807 11056
rect 7484 11052 7490 11054
rect 7097 11051 7163 11052
rect 7741 11051 7807 11054
rect 10777 11114 10843 11117
rect 19517 11114 19583 11117
rect 10777 11112 19583 11114
rect 10777 11056 10782 11112
rect 10838 11056 19522 11112
rect 19578 11056 19583 11112
rect 10777 11054 19583 11056
rect 10777 11051 10843 11054
rect 19517 11051 19583 11054
rect 0 10978 800 11008
rect 933 10978 999 10981
rect 0 10976 999 10978
rect 0 10920 938 10976
rect 994 10920 999 10976
rect 0 10918 999 10920
rect 0 10888 800 10918
rect 933 10915 999 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 7557 10706 7623 10709
rect 16573 10706 16639 10709
rect 7557 10704 16639 10706
rect 7557 10648 7562 10704
rect 7618 10648 16578 10704
rect 16634 10648 16639 10704
rect 7557 10646 16639 10648
rect 7557 10643 7623 10646
rect 16573 10643 16639 10646
rect 0 10570 800 10600
rect 2865 10570 2931 10573
rect 0 10568 2931 10570
rect 0 10512 2870 10568
rect 2926 10512 2931 10568
rect 0 10510 2931 10512
rect 0 10480 800 10510
rect 2865 10507 2931 10510
rect 8845 10570 8911 10573
rect 23381 10570 23447 10573
rect 8845 10568 23447 10570
rect 8845 10512 8850 10568
rect 8906 10512 23386 10568
rect 23442 10512 23447 10568
rect 8845 10510 23447 10512
rect 8845 10507 8911 10510
rect 23381 10507 23447 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 42946 10303 43262 10304
rect 0 10162 800 10192
rect 3325 10162 3391 10165
rect 0 10160 3391 10162
rect 0 10104 3330 10160
rect 3386 10104 3391 10160
rect 0 10102 3391 10104
rect 0 10072 800 10102
rect 3325 10099 3391 10102
rect 12801 10162 12867 10165
rect 16205 10162 16271 10165
rect 12801 10160 16271 10162
rect 12801 10104 12806 10160
rect 12862 10104 16210 10160
rect 16266 10104 16271 10160
rect 12801 10102 16271 10104
rect 12801 10099 12867 10102
rect 16205 10099 16271 10102
rect 7925 10026 7991 10029
rect 7790 10024 7991 10026
rect 7790 9968 7930 10024
rect 7986 9968 7991 10024
rect 7790 9966 7991 9968
rect 7189 9890 7255 9893
rect 7790 9890 7850 9966
rect 7925 9963 7991 9966
rect 13445 10026 13511 10029
rect 15285 10026 15351 10029
rect 16113 10026 16179 10029
rect 17861 10026 17927 10029
rect 18413 10026 18479 10029
rect 13445 10024 18479 10026
rect 13445 9968 13450 10024
rect 13506 9968 15290 10024
rect 15346 9968 16118 10024
rect 16174 9968 17866 10024
rect 17922 9968 18418 10024
rect 18474 9968 18479 10024
rect 13445 9966 18479 9968
rect 13445 9963 13511 9966
rect 15285 9963 15351 9966
rect 16113 9963 16179 9966
rect 17861 9963 17927 9966
rect 18413 9963 18479 9966
rect 7189 9888 7850 9890
rect 7189 9832 7194 9888
rect 7250 9832 7850 9888
rect 7189 9830 7850 9832
rect 7189 9827 7255 9830
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 1577 9754 1643 9757
rect 0 9752 1643 9754
rect 0 9696 1582 9752
rect 1638 9696 1643 9752
rect 0 9694 1643 9696
rect 0 9664 800 9694
rect 1577 9691 1643 9694
rect 5993 9618 6059 9621
rect 9397 9620 9463 9621
rect 6126 9618 6132 9620
rect 5993 9616 6132 9618
rect 5993 9560 5998 9616
rect 6054 9560 6132 9616
rect 5993 9558 6132 9560
rect 5993 9555 6059 9558
rect 6126 9556 6132 9558
rect 6196 9556 6202 9620
rect 9397 9616 9444 9620
rect 9508 9618 9514 9620
rect 10777 9618 10843 9621
rect 18965 9618 19031 9621
rect 9397 9560 9402 9616
rect 9397 9556 9444 9560
rect 9508 9558 9554 9618
rect 10777 9616 19031 9618
rect 10777 9560 10782 9616
rect 10838 9560 18970 9616
rect 19026 9560 19031 9616
rect 10777 9558 19031 9560
rect 9508 9556 9514 9558
rect 9397 9555 9463 9556
rect 10777 9555 10843 9558
rect 18965 9555 19031 9558
rect 4286 9420 4292 9484
rect 4356 9482 4362 9484
rect 6361 9482 6427 9485
rect 4356 9480 6427 9482
rect 4356 9424 6366 9480
rect 6422 9424 6427 9480
rect 4356 9422 6427 9424
rect 4356 9420 4362 9422
rect 6361 9419 6427 9422
rect 9121 9482 9187 9485
rect 34329 9482 34395 9485
rect 9121 9480 34395 9482
rect 9121 9424 9126 9480
rect 9182 9424 34334 9480
rect 34390 9424 34395 9480
rect 9121 9422 34395 9424
rect 9121 9419 9187 9422
rect 34329 9419 34395 9422
rect 0 9346 800 9376
rect 2773 9346 2839 9349
rect 0 9344 2839 9346
rect 0 9288 2778 9344
rect 2834 9288 2839 9344
rect 0 9286 2839 9288
rect 0 9256 800 9286
rect 2773 9283 2839 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 4153 9074 4219 9077
rect 31293 9074 31359 9077
rect 4153 9072 31359 9074
rect 4153 9016 4158 9072
rect 4214 9016 31298 9072
rect 31354 9016 31359 9072
rect 4153 9014 31359 9016
rect 4153 9011 4219 9014
rect 31293 9011 31359 9014
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 7465 8938 7531 8941
rect 24853 8938 24919 8941
rect 7465 8936 24919 8938
rect 7465 8880 7470 8936
rect 7526 8880 24858 8936
rect 24914 8880 24919 8936
rect 7465 8878 24919 8880
rect 7465 8875 7531 8878
rect 24853 8875 24919 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 0 8530 800 8560
rect 933 8530 999 8533
rect 0 8528 999 8530
rect 0 8472 938 8528
rect 994 8472 999 8528
rect 0 8470 999 8472
rect 0 8440 800 8470
rect 933 8467 999 8470
rect 10726 8196 10732 8260
rect 10796 8258 10802 8260
rect 10961 8258 11027 8261
rect 10796 8256 11027 8258
rect 10796 8200 10966 8256
rect 11022 8200 11027 8256
rect 10796 8198 11027 8200
rect 10796 8196 10802 8198
rect 10961 8195 11027 8198
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 1301 8122 1367 8125
rect 0 8120 1367 8122
rect 0 8064 1306 8120
rect 1362 8064 1367 8120
rect 0 8062 1367 8064
rect 0 8032 800 8062
rect 1301 8059 1367 8062
rect 0 7714 800 7744
rect 1761 7714 1827 7717
rect 0 7712 1827 7714
rect 0 7656 1766 7712
rect 1822 7656 1827 7712
rect 0 7654 1827 7656
rect 0 7624 800 7654
rect 1761 7651 1827 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 0 7306 800 7336
rect 2865 7306 2931 7309
rect 0 7304 2931 7306
rect 0 7248 2870 7304
rect 2926 7248 2931 7304
rect 0 7246 2931 7248
rect 0 7216 800 7246
rect 2865 7243 2931 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 0 6898 800 6928
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6808 800 6838
rect 2773 6835 2839 6838
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1209 6490 1275 6493
rect 0 6488 1275 6490
rect 0 6432 1214 6488
rect 1270 6432 1275 6488
rect 0 6430 1275 6432
rect 0 6400 800 6430
rect 1209 6427 1275 6430
rect 0 6082 800 6112
rect 933 6082 999 6085
rect 0 6080 999 6082
rect 0 6024 938 6080
rect 994 6024 999 6080
rect 0 6022 999 6024
rect 0 5992 800 6022
rect 933 6019 999 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 0 5674 800 5704
rect 933 5674 999 5677
rect 0 5672 999 5674
rect 0 5616 938 5672
rect 994 5616 999 5672
rect 0 5614 999 5616
rect 0 5584 800 5614
rect 933 5611 999 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 933 5266 999 5269
rect 0 5264 999 5266
rect 0 5208 938 5264
rect 994 5208 999 5264
rect 0 5206 999 5208
rect 0 5176 800 5206
rect 933 5203 999 5206
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 0 4450 800 4480
rect 1761 4450 1827 4453
rect 0 4448 1827 4450
rect 0 4392 1766 4448
rect 1822 4392 1827 4448
rect 0 4390 1827 4392
rect 0 4360 800 4390
rect 1761 4387 1827 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 0 4042 800 4072
rect 1301 4042 1367 4045
rect 0 4040 1367 4042
rect 0 3984 1306 4040
rect 1362 3984 1367 4040
rect 0 3982 1367 3984
rect 0 3952 800 3982
rect 1301 3979 1367 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 933 3634 999 3637
rect 0 3632 999 3634
rect 0 3576 938 3632
rect 994 3576 999 3632
rect 0 3574 999 3576
rect 0 3544 800 3574
rect 933 3571 999 3574
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 1209 3226 1275 3229
rect 0 3224 1275 3226
rect 0 3168 1214 3224
rect 1270 3168 1275 3224
rect 0 3166 1275 3168
rect 0 3136 800 3166
rect 1209 3163 1275 3166
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 0 2410 800 2440
rect 933 2410 999 2413
rect 0 2408 999 2410
rect 0 2352 938 2408
rect 994 2352 999 2408
rect 0 2350 999 2352
rect 0 2320 800 2350
rect 933 2347 999 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 2773 2002 2839 2005
rect 0 2000 2839 2002
rect 0 1944 2778 2000
rect 2834 1944 2839 2000
rect 0 1942 2839 1944
rect 0 1912 800 1942
rect 2773 1939 2839 1942
rect 0 1594 800 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 800 1534
rect 2865 1531 2931 1534
<< via3 >>
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 9444 24108 9508 24172
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 3924 23428 3988 23492
rect 11652 23428 11716 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 5396 23020 5460 23084
rect 4844 22944 4908 22948
rect 4844 22888 4894 22944
rect 4894 22888 4908 22944
rect 4844 22884 4908 22888
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 3556 22204 3620 22268
rect 22140 22264 22204 22268
rect 22140 22208 22190 22264
rect 22190 22208 22204 22264
rect 22140 22204 22204 22208
rect 7052 21992 7116 21996
rect 7052 21936 7066 21992
rect 7066 21936 7116 21992
rect 7052 21932 7116 21936
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 3740 21660 3804 21724
rect 11652 21388 11716 21452
rect 27660 21388 27724 21452
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 10732 21040 10796 21044
rect 10732 20984 10782 21040
rect 10782 20984 10796 21040
rect 10732 20980 10796 20984
rect 4292 20708 4356 20772
rect 7420 20708 7484 20772
rect 10916 20768 10980 20772
rect 10916 20712 10930 20768
rect 10930 20712 10980 20768
rect 10916 20708 10980 20712
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 11100 19620 11164 19684
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 6132 19348 6196 19412
rect 22324 19348 22388 19412
rect 27660 19212 27724 19276
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 3740 17036 3804 17100
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 3924 16492 3988 16556
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 11100 15736 11164 15740
rect 11100 15680 11150 15736
rect 11150 15680 11164 15736
rect 11100 15676 11164 15680
rect 9996 15404 10060 15468
rect 3556 15268 3620 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 10916 15132 10980 15196
rect 7604 14860 7668 14924
rect 22324 14724 22388 14788
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 9996 14316 10060 14380
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 7604 12276 7668 12340
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 22140 11596 22204 11660
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 5396 11324 5460 11388
rect 4844 11052 4908 11116
rect 7052 11112 7116 11116
rect 7052 11056 7102 11112
rect 7102 11056 7116 11112
rect 7052 11052 7116 11056
rect 7420 11052 7484 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 6132 9556 6196 9620
rect 9444 9616 9508 9620
rect 9444 9560 9458 9616
rect 9458 9560 9508 9616
rect 9444 9556 9508 9560
rect 4292 9420 4356 9484
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 10732 8196 10796 8260
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 7944 23968 8264 24528
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 9443 24172 9509 24173
rect 9443 24108 9444 24172
rect 9508 24108 9509 24172
rect 9443 24107 9509 24108
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 3923 23492 3989 23493
rect 3923 23428 3924 23492
rect 3988 23428 3989 23492
rect 3923 23427 3989 23428
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 3555 22268 3621 22269
rect 3555 22204 3556 22268
rect 3620 22204 3621 22268
rect 3555 22203 3621 22204
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 3558 15333 3618 22203
rect 3739 21724 3805 21725
rect 3739 21660 3740 21724
rect 3804 21660 3805 21724
rect 3739 21659 3805 21660
rect 3742 17101 3802 21659
rect 3739 17100 3805 17101
rect 3739 17036 3740 17100
rect 3804 17036 3805 17100
rect 3739 17035 3805 17036
rect 3926 16557 3986 23427
rect 5395 23084 5461 23085
rect 5395 23020 5396 23084
rect 5460 23020 5461 23084
rect 5395 23019 5461 23020
rect 4843 22948 4909 22949
rect 4843 22884 4844 22948
rect 4908 22884 4909 22948
rect 4843 22883 4909 22884
rect 4291 20772 4357 20773
rect 4291 20708 4292 20772
rect 4356 20708 4357 20772
rect 4291 20707 4357 20708
rect 3923 16556 3989 16557
rect 3923 16492 3924 16556
rect 3988 16492 3989 16556
rect 3923 16491 3989 16492
rect 3555 15332 3621 15333
rect 3555 15268 3556 15332
rect 3620 15268 3621 15332
rect 3555 15267 3621 15268
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 4294 9485 4354 20707
rect 4846 11117 4906 22883
rect 5398 11389 5458 23019
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7051 21996 7117 21997
rect 7051 21932 7052 21996
rect 7116 21932 7117 21996
rect 7051 21931 7117 21932
rect 6131 19412 6197 19413
rect 6131 19348 6132 19412
rect 6196 19348 6197 19412
rect 6131 19347 6197 19348
rect 5395 11388 5461 11389
rect 5395 11324 5396 11388
rect 5460 11324 5461 11388
rect 5395 11323 5461 11324
rect 4843 11116 4909 11117
rect 4843 11052 4844 11116
rect 4908 11052 4909 11116
rect 4843 11051 4909 11052
rect 6134 9621 6194 19347
rect 7054 11117 7114 21931
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7419 20772 7485 20773
rect 7419 20708 7420 20772
rect 7484 20708 7485 20772
rect 7419 20707 7485 20708
rect 7422 11117 7482 20707
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7603 14924 7669 14925
rect 7603 14860 7604 14924
rect 7668 14860 7669 14924
rect 7603 14859 7669 14860
rect 7606 12341 7666 14859
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7603 12340 7669 12341
rect 7603 12276 7604 12340
rect 7668 12276 7669 12340
rect 7603 12275 7669 12276
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7051 11116 7117 11117
rect 7051 11052 7052 11116
rect 7116 11052 7117 11116
rect 7051 11051 7117 11052
rect 7419 11116 7485 11117
rect 7419 11052 7420 11116
rect 7484 11052 7485 11116
rect 7419 11051 7485 11052
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 6131 9620 6197 9621
rect 6131 9556 6132 9620
rect 6196 9556 6197 9620
rect 6131 9555 6197 9556
rect 4291 9484 4357 9485
rect 4291 9420 4292 9484
rect 4356 9420 4357 9484
rect 4291 9419 4357 9420
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 8736 8264 9760
rect 9446 9621 9506 24107
rect 11651 23492 11717 23493
rect 11651 23428 11652 23492
rect 11716 23428 11717 23492
rect 11651 23427 11717 23428
rect 11654 21453 11714 23427
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 11651 21452 11717 21453
rect 11651 21388 11652 21452
rect 11716 21388 11717 21452
rect 11651 21387 11717 21388
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 10731 21044 10797 21045
rect 10731 20980 10732 21044
rect 10796 20980 10797 21044
rect 10731 20979 10797 20980
rect 9995 15468 10061 15469
rect 9995 15404 9996 15468
rect 10060 15404 10061 15468
rect 9995 15403 10061 15404
rect 9998 14381 10058 15403
rect 9995 14380 10061 14381
rect 9995 14316 9996 14380
rect 10060 14316 10061 14380
rect 9995 14315 10061 14316
rect 9443 9620 9509 9621
rect 9443 9556 9444 9620
rect 9508 9556 9509 9620
rect 9443 9555 9509 9556
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 10734 8261 10794 20979
rect 10915 20772 10981 20773
rect 10915 20708 10916 20772
rect 10980 20708 10981 20772
rect 10915 20707 10981 20708
rect 10918 15197 10978 20707
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 11099 19684 11165 19685
rect 11099 19620 11100 19684
rect 11164 19620 11165 19684
rect 11099 19619 11165 19620
rect 11102 15741 11162 19619
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 11099 15740 11165 15741
rect 11099 15676 11100 15740
rect 11164 15676 11165 15740
rect 11099 15675 11165 15676
rect 10915 15196 10981 15197
rect 10915 15132 10916 15196
rect 10980 15132 10981 15196
rect 10915 15131 10981 15132
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 10731 8260 10797 8261
rect 10731 8196 10732 8260
rect 10796 8196 10797 8260
rect 10731 8195 10797 8196
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22139 22268 22205 22269
rect 22139 22204 22140 22268
rect 22204 22204 22205 22268
rect 22139 22203 22205 22204
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 22142 11661 22202 22203
rect 22944 21248 23264 22272
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27659 21452 27725 21453
rect 27659 21388 27660 21452
rect 27724 21388 27725 21452
rect 27659 21387 27725 21388
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22323 19412 22389 19413
rect 22323 19348 22324 19412
rect 22388 19348 22389 19412
rect 22323 19347 22389 19348
rect 22326 14789 22386 19347
rect 22944 19072 23264 20096
rect 27662 19277 27722 21387
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27659 19276 27725 19277
rect 27659 19212 27660 19276
rect 27724 19212 27725 19276
rect 27659 19211 27725 19212
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22323 14788 22389 14789
rect 22323 14724 22324 14788
rect 22388 14724 22389 14788
rect 22323 14723 22389 14724
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22139 11660 22205 11661
rect 22139 11596 22140 11660
rect 22204 11596 22205 11660
rect 22139 11595 22205 11596
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _096_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1676037725
transform 1 0 19504 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _099_
timestamp 1676037725
transform 1 0 13248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _100_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _101_
timestamp 1676037725
transform 1 0 6532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1676037725
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1676037725
transform 1 0 4140 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1676037725
transform 1 0 9200 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 6716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1676037725
transform 1 0 12144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1676037725
transform 1 0 6072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 4140 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 5796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 20976 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 3128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1676037725
transform 1 0 4508 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 3312 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1676037725
transform 1 0 2760 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _132_
timestamp 1676037725
transform 1 0 7452 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _133_
timestamp 1676037725
transform 1 0 9108 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _134_
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 3680 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 35696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 34040 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 34960 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 33304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 33028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 32292 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 34224 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 32568 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 32292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _147_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _149_
timestamp 1676037725
transform 1 0 28244 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _150_
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _152_
timestamp 1676037725
transform 1 0 3956 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _154_
timestamp 1676037725
transform 1 0 18400 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 11408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1676037725
transform 1 0 14996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1676037725
transform 1 0 20332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 14996 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 17020 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 13248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 22172 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 10304 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 4784 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 9292 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 4968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 5336 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 2576 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 7912 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 33948 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 10488 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 7820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 15364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 20148 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 22724 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 30912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 30912 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 23092 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 24472 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 20148 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 21620 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 2852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 5244 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1676037725
transform 1 0 9568 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1676037725
transform 1 0 16376 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1676037725
transform 1 0 22724 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1676037725
transform 1 0 22632 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9292 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6808 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7360 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4140 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 4140 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 4784 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 5336 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 5244 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 7360 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8188 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8464 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6992 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 5520 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10120 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9200 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__190 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9568 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 10396 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13616 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 4048 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 3404 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 9200 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 4048 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6348 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 6900 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__191
timestamp 1676037725
transform 1 0 5152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 5244 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 3956 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 3956 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5152 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7360 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 3956 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14260 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__192
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 8096 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10212 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 6992 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12788 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7820 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10856 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6624 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9384 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 15272 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__193
timestamp 1676037725
transform 1 0 9384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7636 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10580 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28612 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8832 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 26864 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22724 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 25760 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 23000 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22172 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27508 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17112 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9568 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 14352 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 14996 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 13892 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 19504 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 19136 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 23092 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 19688 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 21344 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 25024 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 25300 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1676037725
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1676037725
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1676037725
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 1676037725
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1676037725
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1676037725
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_268
timestamp 1676037725
transform 1 0 25760 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_297
timestamp 1676037725
transform 1 0 28428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_326
timestamp 1676037725
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1676037725
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1676037725
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1676037725
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1676037725
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1676037725
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1676037725
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1676037725
transform 1 0 48668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_22
timestamp 1676037725
transform 1 0 3128 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_34
timestamp 1676037725
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_104
timestamp 1676037725
transform 1 0 10672 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_128
timestamp 1676037725
transform 1 0 12880 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1676037725
transform 1 0 13616 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_142
timestamp 1676037725
transform 1 0 14168 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1676037725
transform 1 0 15272 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1676037725
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_174
timestamp 1676037725
transform 1 0 17112 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_182
timestamp 1676037725
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_188
timestamp 1676037725
transform 1 0 18400 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_200
timestamp 1676037725
transform 1 0 19504 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_208
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_212
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1676037725
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1676037725
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_8
timestamp 1676037725
transform 1 0 1840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp 1676037725
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_116
timestamp 1676037725
transform 1 0 11776 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_128
timestamp 1676037725
transform 1 0 12880 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1676037725
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_22
timestamp 1676037725
transform 1 0 3128 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_34
timestamp 1676037725
transform 1 0 4232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_46
timestamp 1676037725
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1676037725
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_154
timestamp 1676037725
transform 1 0 15272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_205
timestamp 1676037725
transform 1 0 19964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_217
timestamp 1676037725
transform 1 0 21068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_229
timestamp 1676037725
transform 1 0 22172 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1676037725
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1676037725
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_258
timestamp 1676037725
transform 1 0 24840 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_266
timestamp 1676037725
transform 1 0 25576 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1676037725
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1676037725
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_177
timestamp 1676037725
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_186
timestamp 1676037725
transform 1 0 18216 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_198
timestamp 1676037725
transform 1 0 19320 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_210
timestamp 1676037725
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_231
timestamp 1676037725
transform 1 0 22356 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_238
timestamp 1676037725
transform 1 0 23000 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_250
timestamp 1676037725
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_262
timestamp 1676037725
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1676037725
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_320
timestamp 1676037725
transform 1 0 30544 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1676037725
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_173
timestamp 1676037725
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_276
timestamp 1676037725
transform 1 0 26496 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_234
timestamp 1676037725
transform 1 0 22632 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_246
timestamp 1676037725
transform 1 0 23736 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_258
timestamp 1676037725
transform 1 0 24840 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_270
timestamp 1676037725
transform 1 0 25944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1676037725
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1676037725
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1676037725
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_237
timestamp 1676037725
transform 1 0 22908 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_244
timestamp 1676037725
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1676037725
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_89
timestamp 1676037725
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_101
timestamp 1676037725
transform 1 0 10396 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1676037725
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_120
timestamp 1676037725
transform 1 0 12144 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1676037725
transform 1 0 13248 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_139
timestamp 1676037725
transform 1 0 13892 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_151
timestamp 1676037725
transform 1 0 14996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1676037725
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1676037725
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1676037725
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_8
timestamp 1676037725
transform 1 0 1840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_22
timestamp 1676037725
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_75
timestamp 1676037725
transform 1 0 8004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1676037725
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1676037725
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1676037725
transform 1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_120
timestamp 1676037725
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_127
timestamp 1676037725
transform 1 0 12788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1676037725
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_157
timestamp 1676037725
transform 1 0 15548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_169
timestamp 1676037725
transform 1 0 16652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_181
timestamp 1676037725
transform 1 0 17756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1676037725
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp 1676037725
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_8
timestamp 1676037725
transform 1 0 1840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_22
timestamp 1676037725
transform 1 0 3128 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_34
timestamp 1676037725
transform 1 0 4232 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_46
timestamp 1676037725
transform 1 0 5336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_50
timestamp 1676037725
transform 1 0 5704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1676037725
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_63
timestamp 1676037725
transform 1 0 6900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1676037725
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1676037725
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_100
timestamp 1676037725
transform 1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1676037725
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_126
timestamp 1676037725
transform 1 0 12696 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1676037725
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1676037725
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_159
timestamp 1676037725
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_174
timestamp 1676037725
transform 1 0 17112 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_186
timestamp 1676037725
transform 1 0 18216 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_198
timestamp 1676037725
transform 1 0 19320 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_210
timestamp 1676037725
transform 1 0 20424 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1676037725
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1676037725
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1676037725
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1676037725
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1676037725
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_34
timestamp 1676037725
transform 1 0 4232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_47
timestamp 1676037725
transform 1 0 5428 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_51
timestamp 1676037725
transform 1 0 5796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1676037725
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1676037725
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1676037725
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_123
timestamp 1676037725
transform 1 0 12420 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_130
timestamp 1676037725
transform 1 0 13064 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1676037725
transform 1 0 13432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_160
timestamp 1676037725
transform 1 0 15824 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_182
timestamp 1676037725
transform 1 0 17848 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1676037725
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1676037725
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_19
timestamp 1676037725
transform 1 0 2852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_25
timestamp 1676037725
transform 1 0 3404 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_29
timestamp 1676037725
transform 1 0 3772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_36
timestamp 1676037725
transform 1 0 4416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_42
timestamp 1676037725
transform 1 0 4968 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_47
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1676037725
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1676037725
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_135
timestamp 1676037725
transform 1 0 13524 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1676037725
transform 1 0 14260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1676037725
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_191
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_204
timestamp 1676037725
transform 1 0 19872 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_216
timestamp 1676037725
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_294
timestamp 1676037725
transform 1 0 28152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_306
timestamp 1676037725
transform 1 0 29256 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_318
timestamp 1676037725
transform 1 0 30360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_330
timestamp 1676037725
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1676037725
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1676037725
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1676037725
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_47
timestamp 1676037725
transform 1 0 5428 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_54
timestamp 1676037725
transform 1 0 6072 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1676037725
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_89
timestamp 1676037725
transform 1 0 9292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1676037725
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_106
timestamp 1676037725
transform 1 0 10856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1676037725
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1676037725
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1676037725
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_166
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1676037725
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_225
timestamp 1676037725
transform 1 0 21804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_237
timestamp 1676037725
transform 1 0 22908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1676037725
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1676037725
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1676037725
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1676037725
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1676037725
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1676037725
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1676037725
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1676037725
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1676037725
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1676037725
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_20
timestamp 1676037725
transform 1 0 2944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_32
timestamp 1676037725
transform 1 0 4048 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_40
timestamp 1676037725
transform 1 0 4784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_44
timestamp 1676037725
transform 1 0 5152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_64
timestamp 1676037725
transform 1 0 6992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_91
timestamp 1676037725
transform 1 0 9476 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_99
timestamp 1676037725
transform 1 0 10212 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1676037725
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_139
timestamp 1676037725
transform 1 0 13892 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_143
timestamp 1676037725
transform 1 0 14260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1676037725
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1676037725
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1676037725
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1676037725
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1676037725
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1676037725
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1676037725
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1676037725
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1676037725
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1676037725
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1676037725
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1676037725
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1676037725
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_517
timestamp 1676037725
transform 1 0 48668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_12
timestamp 1676037725
transform 1 0 2208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_34
timestamp 1676037725
transform 1 0 4232 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_60
timestamp 1676037725
transform 1 0 6624 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_69
timestamp 1676037725
transform 1 0 7452 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1676037725
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_96
timestamp 1676037725
transform 1 0 9936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_168
timestamp 1676037725
transform 1 0 16560 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_211
timestamp 1676037725
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_235
timestamp 1676037725
transform 1 0 22724 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1676037725
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1676037725
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1676037725
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_334
timestamp 1676037725
transform 1 0 31832 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_346
timestamp 1676037725
transform 1 0 32936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1676037725
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1676037725
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1676037725
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1676037725
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1676037725
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1676037725
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1676037725
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1676037725
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1676037725
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_10
timestamp 1676037725
transform 1 0 2024 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_21
timestamp 1676037725
transform 1 0 3036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1676037725
transform 1 0 3772 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_40
timestamp 1676037725
transform 1 0 4784 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1676037725
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1676037725
transform 1 0 6808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1676037725
transform 1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1676037725
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_117
timestamp 1676037725
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_151
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_194
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_251
timestamp 1676037725
transform 1 0 24196 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_263
timestamp 1676037725
transform 1 0 25300 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1676037725
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1676037725
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1676037725
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1676037725
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1676037725
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1676037725
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1676037725
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1676037725
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_517
timestamp 1676037725
transform 1 0 48668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_19
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1676037725
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_45
timestamp 1676037725
transform 1 0 5244 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 1676037725
transform 1 0 7452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1676037725
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_155
timestamp 1676037725
transform 1 0 15364 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1676037725
transform 1 0 16100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_185
timestamp 1676037725
transform 1 0 18124 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1676037725
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_205
timestamp 1676037725
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1676037725
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1676037725
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1676037725
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1676037725
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1676037725
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1676037725
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1676037725
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1676037725
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1676037725
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1676037725
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1676037725
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1676037725
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1676037725
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1676037725
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1676037725
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1676037725
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_21
timestamp 1676037725
transform 1 0 3036 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1676037725
transform 1 0 3680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_41
timestamp 1676037725
transform 1 0 4876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1676037725
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_63
timestamp 1676037725
transform 1 0 6900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_73
timestamp 1676037725
transform 1 0 7820 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_100
timestamp 1676037725
transform 1 0 10304 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_106
timestamp 1676037725
transform 1 0 10856 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_117
timestamp 1676037725
transform 1 0 11868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_121
timestamp 1676037725
transform 1 0 12236 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1676037725
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1676037725
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1676037725
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_174
timestamp 1676037725
transform 1 0 17112 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1676037725
transform 1 0 17848 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_192
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_207
timestamp 1676037725
transform 1 0 20148 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_258
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_270
timestamp 1676037725
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1676037725
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1676037725
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1676037725
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1676037725
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1676037725
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1676037725
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1676037725
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1676037725
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1676037725
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1676037725
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1676037725
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1676037725
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1676037725
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1676037725
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1676037725
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_95
timestamp 1676037725
transform 1 0 9844 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_108
timestamp 1676037725
transform 1 0 11040 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1676037725
transform 1 0 16744 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_202
timestamp 1676037725
transform 1 0 19688 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_208
timestamp 1676037725
transform 1 0 20240 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_229
timestamp 1676037725
transform 1 0 22172 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_235
timestamp 1676037725
transform 1 0 22724 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1676037725
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_266
timestamp 1676037725
transform 1 0 25576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_278
timestamp 1676037725
transform 1 0 26680 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_290
timestamp 1676037725
transform 1 0 27784 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1676037725
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1676037725
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1676037725
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1676037725
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1676037725
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1676037725
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1676037725
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1676037725
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1676037725
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1676037725
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1676037725
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1676037725
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1676037725
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_35
timestamp 1676037725
transform 1 0 4324 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_43
timestamp 1676037725
transform 1 0 5060 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1676037725
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1676037725
transform 1 0 7728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_85
timestamp 1676037725
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_117
timestamp 1676037725
transform 1 0 11868 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1676037725
transform 1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_140
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1676037725
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1676037725
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_206
timestamp 1676037725
transform 1 0 20056 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_216
timestamp 1676037725
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1676037725
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1676037725
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1676037725
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1676037725
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1676037725
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1676037725
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1676037725
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1676037725
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1676037725
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1676037725
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1676037725
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1676037725
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1676037725
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1676037725
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1676037725
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1676037725
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1676037725
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1676037725
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_40
timestamp 1676037725
transform 1 0 4784 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_44
timestamp 1676037725
transform 1 0 5152 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1676037725
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_72
timestamp 1676037725
transform 1 0 7728 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_89
timestamp 1676037725
transform 1 0 9292 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1676037725
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_112
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_222
timestamp 1676037725
transform 1 0 21528 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_264
timestamp 1676037725
transform 1 0 25392 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1676037725
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1676037725
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1676037725
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1676037725
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1676037725
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1676037725
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1676037725
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1676037725
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1676037725
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1676037725
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1676037725
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1676037725
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1676037725
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1676037725
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1676037725
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1676037725
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1676037725
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1676037725
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_25
timestamp 1676037725
transform 1 0 3404 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_29
timestamp 1676037725
transform 1 0 3772 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1676037725
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_63
timestamp 1676037725
transform 1 0 6900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_67
timestamp 1676037725
transform 1 0 7268 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_77
timestamp 1676037725
transform 1 0 8188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1676037725
transform 1 0 8832 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_97
timestamp 1676037725
transform 1 0 10028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_138
timestamp 1676037725
transform 1 0 13800 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1676037725
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_194
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_198
timestamp 1676037725
transform 1 0 19320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_208
timestamp 1676037725
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_247
timestamp 1676037725
transform 1 0 23828 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_255
timestamp 1676037725
transform 1 0 24564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1676037725
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1676037725
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1676037725
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1676037725
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1676037725
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1676037725
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1676037725
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1676037725
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1676037725
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1676037725
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1676037725
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1676037725
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_517
timestamp 1676037725
transform 1 0 48668 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp 1676037725
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_66
timestamp 1676037725
transform 1 0 7176 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_72
timestamp 1676037725
transform 1 0 7728 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_91
timestamp 1676037725
transform 1 0 9476 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1676037725
transform 1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1676037725
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_128
timestamp 1676037725
transform 1 0 12880 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_134
timestamp 1676037725
transform 1 0 13432 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_147
timestamp 1676037725
transform 1 0 14628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_157
timestamp 1676037725
transform 1 0 15548 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_170
timestamp 1676037725
transform 1 0 16744 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1676037725
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_226
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1676037725
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_271
timestamp 1676037725
transform 1 0 26036 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_283
timestamp 1676037725
transform 1 0 27140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_295
timestamp 1676037725
transform 1 0 28244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1676037725
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1676037725
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1676037725
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1676037725
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1676037725
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1676037725
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1676037725
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1676037725
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1676037725
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_41
timestamp 1676037725
transform 1 0 4876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_63
timestamp 1676037725
transform 1 0 6900 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_76
timestamp 1676037725
transform 1 0 8096 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_101
timestamp 1676037725
transform 1 0 10396 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_139
timestamp 1676037725
transform 1 0 13892 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_154
timestamp 1676037725
transform 1 0 15272 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_162
timestamp 1676037725
transform 1 0 16008 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1676037725
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_203
timestamp 1676037725
transform 1 0 19780 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_209
timestamp 1676037725
transform 1 0 20332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_231
timestamp 1676037725
transform 1 0 22356 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_250
timestamp 1676037725
transform 1 0 24104 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1676037725
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1676037725
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1676037725
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1676037725
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1676037725
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1676037725
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1676037725
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1676037725
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1676037725
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1676037725
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_517
timestamp 1676037725
transform 1 0 48668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1676037725
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_55
timestamp 1676037725
transform 1 0 6164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_59
timestamp 1676037725
transform 1 0 6532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1676037725
transform 1 0 7452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1676037725
transform 1 0 9476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_107
timestamp 1676037725
transform 1 0 10948 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_115
timestamp 1676037725
transform 1 0 11684 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_147
timestamp 1676037725
transform 1 0 14628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_160
timestamp 1676037725
transform 1 0 15824 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_168
timestamp 1676037725
transform 1 0 16560 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1676037725
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_179
timestamp 1676037725
transform 1 0 17572 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_186
timestamp 1676037725
transform 1 0 18216 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1676037725
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_222
timestamp 1676037725
transform 1 0 21528 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1676037725
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1676037725
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1676037725
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_299
timestamp 1676037725
transform 1 0 28612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1676037725
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1676037725
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1676037725
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1676037725
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1676037725
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1676037725
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1676037725
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1676037725
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1676037725
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1676037725
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1676037725
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1676037725
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_21
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1676037725
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_61
timestamp 1676037725
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1676037725
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1676037725
transform 1 0 12420 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_133
timestamp 1676037725
transform 1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_152
timestamp 1676037725
transform 1 0 15088 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_180
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1676037725
transform 1 0 18032 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_205
timestamp 1676037725
transform 1 0 19964 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_235
timestamp 1676037725
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_250
timestamp 1676037725
transform 1 0 24104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_256
timestamp 1676037725
transform 1 0 24656 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1676037725
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_287
timestamp 1676037725
transform 1 0 27508 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_311
timestamp 1676037725
transform 1 0 29716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_323
timestamp 1676037725
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1676037725
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1676037725
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1676037725
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1676037725
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1676037725
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1676037725
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1676037725
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1676037725
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1676037725
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1676037725
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1676037725
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_37
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1676037725
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1676037725
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_102
timestamp 1676037725
transform 1 0 10488 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_112
timestamp 1676037725
transform 1 0 11408 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_147
timestamp 1676037725
transform 1 0 14628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_154
timestamp 1676037725
transform 1 0 15272 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_161
timestamp 1676037725
transform 1 0 15916 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_185
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_202
timestamp 1676037725
transform 1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_206
timestamp 1676037725
transform 1 0 20056 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_212
timestamp 1676037725
transform 1 0 20608 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_222
timestamp 1676037725
transform 1 0 21528 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_257
timestamp 1676037725
transform 1 0 24748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_298
timestamp 1676037725
transform 1 0 28520 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1676037725
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_320
timestamp 1676037725
transform 1 0 30544 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_326
timestamp 1676037725
transform 1 0 31096 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_338
timestamp 1676037725
transform 1 0 32200 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_350
timestamp 1676037725
transform 1 0 33304 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1676037725
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1676037725
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1676037725
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1676037725
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1676037725
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1676037725
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1676037725
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1676037725
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1676037725
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1676037725
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1676037725
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_41
timestamp 1676037725
transform 1 0 4876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1676037725
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_75
timestamp 1676037725
transform 1 0 8004 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_92
timestamp 1676037725
transform 1 0 9568 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_100
timestamp 1676037725
transform 1 0 10304 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_128
timestamp 1676037725
transform 1 0 12880 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_134
timestamp 1676037725
transform 1 0 13432 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_148
timestamp 1676037725
transform 1 0 14720 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1676037725
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_178
timestamp 1676037725
transform 1 0 17480 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_186
timestamp 1676037725
transform 1 0 18216 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_198
timestamp 1676037725
transform 1 0 19320 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_211
timestamp 1676037725
transform 1 0 20516 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1676037725
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_274
timestamp 1676037725
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_286
timestamp 1676037725
transform 1 0 27416 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_292
timestamp 1676037725
transform 1 0 27968 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1676037725
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_326
timestamp 1676037725
transform 1 0 31096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1676037725
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1676037725
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1676037725
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1676037725
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1676037725
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1676037725
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1676037725
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1676037725
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1676037725
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_517
timestamp 1676037725
transform 1 0 48668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_36
timestamp 1676037725
transform 1 0 4416 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_60
timestamp 1676037725
transform 1 0 6624 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_96
timestamp 1676037725
transform 1 0 9936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_102
timestamp 1676037725
transform 1 0 10488 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_115
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_128
timestamp 1676037725
transform 1 0 12880 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1676037725
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_148
timestamp 1676037725
transform 1 0 14720 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_172
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 1676037725
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1676037725
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_201
timestamp 1676037725
transform 1 0 19596 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1676037725
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_217
timestamp 1676037725
transform 1 0 21068 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_238
timestamp 1676037725
transform 1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1676037725
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1676037725
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_258
timestamp 1676037725
transform 1 0 24840 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1676037725
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_297
timestamp 1676037725
transform 1 0 28428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1676037725
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_320
timestamp 1676037725
transform 1 0 30544 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_326
timestamp 1676037725
transform 1 0 31096 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_338
timestamp 1676037725
transform 1 0 32200 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_350
timestamp 1676037725
transform 1 0 33304 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1676037725
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1676037725
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1676037725
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1676037725
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1676037725
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1676037725
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1676037725
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1676037725
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1676037725
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1676037725
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1676037725
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_63
timestamp 1676037725
transform 1 0 6900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_84
timestamp 1676037725
transform 1 0 8832 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1676037725
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_135
timestamp 1676037725
transform 1 0 13524 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_150
timestamp 1676037725
transform 1 0 14904 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1676037725
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_184
timestamp 1676037725
transform 1 0 18032 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_194
timestamp 1676037725
transform 1 0 18952 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_231
timestamp 1676037725
transform 1 0 22356 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_241
timestamp 1676037725
transform 1 0 23276 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_254
timestamp 1676037725
transform 1 0 24472 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_271
timestamp 1676037725
transform 1 0 26036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_287
timestamp 1676037725
transform 1 0 27508 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_291
timestamp 1676037725
transform 1 0 27876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_295
timestamp 1676037725
transform 1 0 28244 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_316
timestamp 1676037725
transform 1 0 30176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1676037725
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1676037725
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1676037725
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1676037725
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1676037725
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1676037725
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1676037725
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1676037725
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_517
timestamp 1676037725
transform 1 0 48668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1676037725
transform 1 0 6348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_92
timestamp 1676037725
transform 1 0 9568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_116
timestamp 1676037725
transform 1 0 11776 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_124
timestamp 1676037725
transform 1 0 12512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_128
timestamp 1676037725
transform 1 0 12880 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 1676037725
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_166
timestamp 1676037725
transform 1 0 16376 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1676037725
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_204
timestamp 1676037725
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_228
timestamp 1676037725
transform 1 0 22080 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_237
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_295
timestamp 1676037725
transform 1 0 28244 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_321
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_334
timestamp 1676037725
transform 1 0 31832 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_346
timestamp 1676037725
transform 1 0 32936 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_358
timestamp 1676037725
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1676037725
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1676037725
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1676037725
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1676037725
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1676037725
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1676037725
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1676037725
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1676037725
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1676037725
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1676037725
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_99
timestamp 1676037725
transform 1 0 10212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1676037725
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_123
timestamp 1676037725
transform 1 0 12420 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_133
timestamp 1676037725
transform 1 0 13340 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1676037725
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_194
timestamp 1676037725
transform 1 0 18952 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_231
timestamp 1676037725
transform 1 0 22356 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_248
timestamp 1676037725
transform 1 0 23920 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_272
timestamp 1676037725
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1676037725
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 1676037725
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1676037725
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1676037725
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1676037725
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1676037725
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1676037725
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1676037725
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1676037725
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1676037725
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1676037725
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_517
timestamp 1676037725
transform 1 0 48668 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1676037725
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_42
timestamp 1676037725
transform 1 0 4968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_68
timestamp 1676037725
transform 1 0 7360 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1676037725
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_103
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_114
timestamp 1676037725
transform 1 0 11592 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_134
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_162
timestamp 1676037725
transform 1 0 16008 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_168
timestamp 1676037725
transform 1 0 16560 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1676037725
transform 1 0 17756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_219
timestamp 1676037725
transform 1 0 21252 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_231
timestamp 1676037725
transform 1 0 22356 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1676037725
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_291
timestamp 1676037725
transform 1 0 27876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_321
timestamp 1676037725
transform 1 0 30636 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_335
timestamp 1676037725
transform 1 0 31924 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_343
timestamp 1676037725
transform 1 0 32660 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_355
timestamp 1676037725
transform 1 0 33764 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1676037725
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1676037725
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1676037725
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1676037725
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1676037725
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1676037725
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1676037725
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1676037725
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1676037725
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_85
timestamp 1676037725
transform 1 0 8924 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_91
timestamp 1676037725
transform 1 0 9476 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_104
timestamp 1676037725
transform 1 0 10672 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_126
timestamp 1676037725
transform 1 0 12696 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_147
timestamp 1676037725
transform 1 0 14628 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_211
timestamp 1676037725
transform 1 0 20516 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1676037725
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1676037725
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_293
timestamp 1676037725
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_317
timestamp 1676037725
transform 1 0 30268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_330
timestamp 1676037725
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_343
timestamp 1676037725
transform 1 0 32660 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_350
timestamp 1676037725
transform 1 0 33304 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_362
timestamp 1676037725
transform 1 0 34408 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_374
timestamp 1676037725
transform 1 0 35512 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_386
timestamp 1676037725
transform 1 0 36616 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1676037725
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1676037725
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1676037725
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1676037725
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1676037725
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1676037725
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_47
timestamp 1676037725
transform 1 0 5428 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_58
timestamp 1676037725
transform 1 0 6440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_78
timestamp 1676037725
transform 1 0 8280 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_98
timestamp 1676037725
transform 1 0 10120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_120
timestamp 1676037725
transform 1 0 12144 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_147
timestamp 1676037725
transform 1 0 14628 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_169
timestamp 1676037725
transform 1 0 16652 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_173
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_203
timestamp 1676037725
transform 1 0 19780 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_225
timestamp 1676037725
transform 1 0 21804 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 1676037725
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1676037725
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_295
timestamp 1676037725
transform 1 0 28244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 1676037725
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_324
timestamp 1676037725
transform 1 0 30912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_332
timestamp 1676037725
transform 1 0 31648 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_340
timestamp 1676037725
transform 1 0 32384 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_352
timestamp 1676037725
transform 1 0 33488 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1676037725
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1676037725
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1676037725
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1676037725
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1676037725
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1676037725
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_513
timestamp 1676037725
transform 1 0 48300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1676037725
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_70
timestamp 1676037725
transform 1 0 7544 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_92
timestamp 1676037725
transform 1 0 9568 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_119
timestamp 1676037725
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_143
timestamp 1676037725
transform 1 0 14260 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1676037725
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_231
timestamp 1676037725
transform 1 0 22356 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_235
timestamp 1676037725
transform 1 0 22724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1676037725
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_272
timestamp 1676037725
transform 1 0 26128 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_292
timestamp 1676037725
transform 1 0 27968 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_316
timestamp 1676037725
transform 1 0 30176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1676037725
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1676037725
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_343
timestamp 1676037725
transform 1 0 32660 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_351
timestamp 1676037725
transform 1 0 33396 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_366
timestamp 1676037725
transform 1 0 34776 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_378
timestamp 1676037725
transform 1 0 35880 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1676037725
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_399
timestamp 1676037725
transform 1 0 37812 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_420
timestamp 1676037725
transform 1 0 39744 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_432
timestamp 1676037725
transform 1 0 40848 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_444
timestamp 1676037725
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1676037725
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1676037725
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_63
timestamp 1676037725
transform 1 0 6900 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_108
timestamp 1676037725
transform 1 0 11040 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1676037725
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_147
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1676037725
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1676037725
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1676037725
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_277
timestamp 1676037725
transform 1 0 26588 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_305
timestamp 1676037725
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_331
timestamp 1676037725
transform 1 0 31556 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_338
timestamp 1676037725
transform 1 0 32200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_346
timestamp 1676037725
transform 1 0 32936 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_354
timestamp 1676037725
transform 1 0 33672 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1676037725
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1676037725
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1676037725
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1676037725
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1676037725
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1676037725
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1676037725
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1676037725
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_513
timestamp 1676037725
transform 1 0 48300 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_517
timestamp 1676037725
transform 1 0 48668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_9
timestamp 1676037725
transform 1 0 1932 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1676037725
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_63
timestamp 1676037725
transform 1 0 6900 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1676037725
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1676037725
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1676037725
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_212
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1676037725
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1676037725
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1676037725
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_303
timestamp 1676037725
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_310
timestamp 1676037725
transform 1 0 29624 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_324
timestamp 1676037725
transform 1 0 30912 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_331
timestamp 1676037725
transform 1 0 31556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_342
timestamp 1676037725
transform 1 0 32568 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_349
timestamp 1676037725
transform 1 0 33212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_356
timestamp 1676037725
transform 1 0 33856 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_364
timestamp 1676037725
transform 1 0 34592 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_372
timestamp 1676037725
transform 1 0 35328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_380
timestamp 1676037725
transform 1 0 36064 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_387
timestamp 1676037725
transform 1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1676037725
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_397
timestamp 1676037725
transform 1 0 37628 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_401
timestamp 1676037725
transform 1 0 37996 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_413
timestamp 1676037725
transform 1 0 39100 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_425
timestamp 1676037725
transform 1 0 40204 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_440
timestamp 1676037725
transform 1 0 41584 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_465
timestamp 1676037725
transform 1 0 43884 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_485
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_493
timestamp 1676037725
transform 1 0 46460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1676037725
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_517
timestamp 1676037725
transform 1 0 48668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_525
timestamp 1676037725
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1676037725
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1676037725
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1676037725
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1676037725
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1676037725
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_299
timestamp 1676037725
transform 1 0 28612 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1676037725
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_327
timestamp 1676037725
transform 1 0 31188 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_331
timestamp 1676037725
transform 1 0 31556 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_335
timestamp 1676037725
transform 1 0 31924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1676037725
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_342
timestamp 1676037725
transform 1 0 32568 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_348
timestamp 1676037725
transform 1 0 33120 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_353
timestamp 1676037725
transform 1 0 33580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1676037725
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_371
timestamp 1676037725
transform 1 0 35236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_379
timestamp 1676037725
transform 1 0 35972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_386
timestamp 1676037725
transform 1 0 36616 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1676037725
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_398
timestamp 1676037725
transform 1 0 37720 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_404
timestamp 1676037725
transform 1 0 38272 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_409
timestamp 1676037725
transform 1 0 38732 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_417
timestamp 1676037725
transform 1 0 39468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_433
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_440
timestamp 1676037725
transform 1 0 41584 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1676037725
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_471
timestamp 1676037725
transform 1 0 44436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1676037725
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_483
timestamp 1676037725
transform 1 0 45540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_491
timestamp 1676037725
transform 1 0 46276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_499
timestamp 1676037725
transform 1 0 47012 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1676037725
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1676037725
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_511
timestamp 1676037725
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_519
timestamp 1676037725
transform 1 0 48852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 48392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1676037725
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 3128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 2852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1676037725
transform 1 0 32292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1676037725
transform 1 0 29992 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 31280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 32936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 33580 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1676037725
transform 1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1676037725
transform 1 0 33948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 34868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 28612 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 35604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 36340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 36432 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 37444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 37720 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1676037725
transform 1 0 38364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1676037725
transform 1 0 39100 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 40020 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 41308 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1676037725
transform 1 0 41308 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1676037725
transform 1 0 7268 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1676037725
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 28980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 28336 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 29348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1676037725
transform 1 0 31280 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 33488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1676037725
transform 1 0 36064 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  input68
timestamp 1676037725
transform 1 0 42596 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1676037725
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 46644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1676037725
transform 1 0 46736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1676037725
transform 1 0 47748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1676037725
transform 1 0 48484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 44252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 49036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 49036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1676037725
transform 1 0 49036 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1676037725
transform 1 0 48300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 3404 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 3404 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 3404 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 3956 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 6992 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 6532 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 3404 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 9200 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 10672 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 11960 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 12328 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 17204 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 15272 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 14904 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 16928 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 5428 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 6808 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 8096 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 9476 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 12144 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18676 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21160 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18768 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20056 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24288 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25852 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26036 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25760 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27324 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28428 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28336 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 26680 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24748 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37904 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27876 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 24840 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24840 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22356 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20884 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19688 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23000 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17480 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16008 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14720 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14628 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12052 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11224 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11500 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12052 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9936 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8372 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 4784 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7084 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9200 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11408 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12420 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12788 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15088 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18124 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31004 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27784 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_1.mux_l1_in_1__194
timestamp 1676037725
transform 1 0 27232 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17112 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_3.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 18584 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31280 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_5.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16928 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10672 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_7.mux_l1_in_1__162
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14352 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_9.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9384 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25760 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_11.mux_l2_in_0__195
timestamp 1676037725
transform 1 0 31924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 1748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14352 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_13.mux_l2_in_0__196
timestamp 1676037725
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28336 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_15.mux_l2_in_0__197
timestamp 1676037725
transform 1 0 18584 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25760 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_17.mux_l2_in_0__198
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_19.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 21252 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_29.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 22632 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22448 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9568 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27232 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_31.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23092 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_33.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 22448 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30544 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_35.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 24196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30084 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_45.mux_l2_in_0__157
timestamp 1676037725
transform 1 0 27968 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25576 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30636 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_47.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 26404 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30544 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l2_in_0_
timestamp 1676037725
transform 1 0 27600 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_49.mux_l2_in_0__159
timestamp 1676037725
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17296 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_51.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 21252 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_0.mux_l2_in_1__164
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 20700 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23644 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23368 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25760 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_2.mux_l2_in_1__170
timestamp 1676037725
transform 1 0 15456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 13064 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19044 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23184 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22172 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17940 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11868 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_4.mux_l2_in_1__181
timestamp 1676037725
transform 1 0 13156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17940 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 13800 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_6.mux_l2_in_1__188
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19412 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24656 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_8.mux_l2_in_1__189
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20148 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23368 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_10.mux_l2_in_1__165
timestamp 1676037725
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14996 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_12.mux_l1_in_1__166
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_14.mux_l1_in_1__167
timestamp 1676037725
transform 1 0 10672 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_1_
timestamp 1676037725
transform 1 0 9844 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_1_
timestamp 1676037725
transform 1 0 11592 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_16.mux_l1_in_1__168
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10212 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21896 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13156 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_18.mux_l1_in_1__169
timestamp 1676037725
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15916 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_20.mux_l2_in_0__171
timestamp 1676037725
transform 1 0 16652 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14720 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_22.mux_l2_in_0__172
timestamp 1676037725
transform 1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14352 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_24.mux_l2_in_0__173
timestamp 1676037725
transform 1 0 15640 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14444 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3404 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10304 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_26.mux_l2_in_0__174
timestamp 1676037725
transform 1 0 13432 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10488 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10304 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10304 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_28.mux_l2_in_0__175
timestamp 1676037725
transform 1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5152 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12052 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_30.mux_l2_in_0__176
timestamp 1676037725
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12052 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_32.mux_l2_in_0__177
timestamp 1676037725
transform 1 0 12512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27600 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10856 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_34.mux_l2_in_0__178
timestamp 1676037725
transform 1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 33028 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12052 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_36.mux_l2_in_0__179
timestamp 1676037725
transform 1 0 4140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 7268 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 4140 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_38.mux_l2_in_0__180
timestamp 1676037725
transform 1 0 5520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 8004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 6716 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_40.mux_l2_in_0__182
timestamp 1676037725
transform 1 0 1932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_42.mux_l2_in_0__183
timestamp 1676037725
transform 1 0 34500 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9292 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17848 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_44.mux_l1_in_1__184
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 34132 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_46.mux_l1_in_1__185
timestamp 1676037725
transform 1 0 7176 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32568 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19688 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_1_
timestamp 1676037725
transform 1 0 11776 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_48.mux_l1_in_1__186
timestamp 1676037725
transform 1 0 3496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15088 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_50.mux_l1_in_1__187
timestamp 1676037725
transform 1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31004 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 66 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 67 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 68 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 69 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 70 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 71 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 72 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 73 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 74 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 75 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 76 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 77 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 78 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 79 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 80 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 81 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 82 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 83 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 84 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 85 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 86 nsew signal input
flabel metal2 s 40866 26200 40922 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 87 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 88 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 89 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 90 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 91 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 92 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 93 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 94 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 95 nsew signal input
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 96 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 97 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 98 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 99 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 100 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 101 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 102 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 103 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 104 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 105 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 106 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 107 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 108 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 109 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 110 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 111 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 112 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 113 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 114 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 115 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 116 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 117 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 41510 26200 41566 27000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 140 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 reset_top_in
port 141 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 test_enable_top_in
port 142 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 143 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 144 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 145 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 146 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 147 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 148 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 149 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 150 nsew signal input
flabel metal3 s 50200 21904 51000 22024 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 151 nsew signal input
flabel metal3 s 50200 22856 51000 22976 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 152 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 50200 24760 51000 24880 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 154 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 155 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 156 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 158 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal1 17020 5202 17020 5202 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 15594 6222 15594 6222 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 15548 5746 15548 5746 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 12650 7888 12650 7888 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal2 21298 16864 21298 16864 0 cbx_8__0_.cbx_8__0_.ccff_head
rlabel metal1 9154 9894 9154 9894 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 12650 13804 12650 13804 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 8970 14450 8970 14450 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 10028 9350 10028 9350 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 5704 12138 5704 12138 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal1 4186 22542 4186 22542 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 6900 9622 6900 9622 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 5842 13804 5842 13804 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 7682 12682 7682 12682 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal1 5704 21454 5704 21454 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal2 12650 16592 12650 16592 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 8372 13430 8372 13430 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal2 5934 17476 5934 17476 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 7590 17102 7590 17102 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 9384 19482 9384 19482 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal1 8418 14382 8418 14382 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9752 7514 9752 7514 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 13846 8194 13846 8194 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 8234 14416 8234 14416 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 7866 15742 7866 15742 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9522 14994 9522 14994 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11546 14042 11546 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8096 11186 8096 11186 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8326 11118 8326 11118 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9706 7378 9706 7378 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10028 7514 10028 7514 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10580 8942 10580 8942 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 4324 12410 4324 12410 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 4830 10778 4830 10778 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 12098 7412 12098 7412 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 4462 14093 4462 14093 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6808 15402 6808 15402 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 6854 15334 6854 15334 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 7406 9452 7406 9452 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 4922 12954 4922 12954 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6026 14042 6026 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 6946 10098 6946 10098 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 5474 10642 5474 10642 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 4968 14042 4968 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 4462 18428 4462 18428 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 7406 13056 7406 13056 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 12558 12070 12558 12070 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 4048 14586 4048 14586 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6302 13906 6302 13906 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7314 14416 7314 14416 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8326 12308 8326 12308 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8648 14042 8648 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6946 14008 6946 14008 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9292 12410 9292 12410 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 13662 15045 13662 15045 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 7544 12954 7544 12954 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 7314 17952 7314 17952 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10212 17782 10212 17782 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 4784 19142 4784 19142 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 7222 18802 7222 18802 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6210 16626 6210 16626 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7452 15674 7452 15674 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10396 14382 10396 14382 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 6992 17306 6992 17306 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6670 16456 6670 16456 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9890 14552 9890 14552 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 13754 17561 13754 17561 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 6302 19482 6302 19482 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 17434 4284 17434 4284 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 23362 4590 23362 4590 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal2 20562 4012 20562 4012 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal2 28842 4964 28842 4964 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 22494 6834 22494 6834 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 22557 5202 22557 5202 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 18124 3026 18124 3026 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal2 27094 5474 27094 5474 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 23644 6970 23644 6970 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel via1 22143 5202 22143 5202 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 17066 4284 17066 4284 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal2 25990 4760 25990 4760 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 22527 6290 22527 6290 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 15226 6052 15226 6052 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal2 24794 5916 24794 5916 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 1426 823 1426 823 0 ccff_head
rlabel metal2 48622 24694 48622 24694 0 ccff_head_1
rlabel metal2 49174 21233 49174 21233 0 ccff_tail
rlabel metal2 2254 22314 2254 22314 0 ccff_tail_0
rlabel metal3 1786 1564 1786 1564 0 chanx_left_in[0]
rlabel metal3 820 5644 820 5644 0 chanx_left_in[10]
rlabel metal3 820 6052 820 6052 0 chanx_left_in[11]
rlabel metal3 958 6460 958 6460 0 chanx_left_in[12]
rlabel metal2 2806 7123 2806 7123 0 chanx_left_in[13]
rlabel metal2 2898 7021 2898 7021 0 chanx_left_in[14]
rlabel metal3 1234 7684 1234 7684 0 chanx_left_in[15]
rlabel metal3 1004 8092 1004 8092 0 chanx_left_in[16]
rlabel metal3 820 8500 820 8500 0 chanx_left_in[17]
rlabel metal3 1050 8908 1050 8908 0 chanx_left_in[18]
rlabel metal2 2806 8585 2806 8585 0 chanx_left_in[19]
rlabel metal3 1740 1972 1740 1972 0 chanx_left_in[1]
rlabel metal3 1142 9724 1142 9724 0 chanx_left_in[20]
rlabel metal2 3358 9537 3358 9537 0 chanx_left_in[21]
rlabel metal2 2898 9503 2898 9503 0 chanx_left_in[22]
rlabel metal3 820 10948 820 10948 0 chanx_left_in[23]
rlabel metal3 1119 11356 1119 11356 0 chanx_left_in[24]
rlabel metal2 3450 10659 3450 10659 0 chanx_left_in[25]
rlabel metal3 1119 12172 1119 12172 0 chanx_left_in[26]
rlabel metal3 1234 12580 1234 12580 0 chanx_left_in[27]
rlabel metal1 1794 8534 1794 8534 0 chanx_left_in[28]
rlabel metal3 1142 13396 1142 13396 0 chanx_left_in[29]
rlabel metal3 820 2380 820 2380 0 chanx_left_in[2]
rlabel metal3 820 2788 820 2788 0 chanx_left_in[3]
rlabel metal3 958 3196 958 3196 0 chanx_left_in[4]
rlabel metal3 820 3604 820 3604 0 chanx_left_in[5]
rlabel metal3 1004 4012 1004 4012 0 chanx_left_in[6]
rlabel metal3 1234 4420 1234 4420 0 chanx_left_in[7]
rlabel metal3 820 4828 820 4828 0 chanx_left_in[8]
rlabel metal3 820 5236 820 5236 0 chanx_left_in[9]
rlabel metal3 1694 13804 1694 13804 0 chanx_left_out[0]
rlabel metal3 1602 17884 1602 17884 0 chanx_left_out[10]
rlabel metal3 1372 18292 1372 18292 0 chanx_left_out[11]
rlabel metal3 1050 18700 1050 18700 0 chanx_left_out[12]
rlabel metal2 2806 19737 2806 19737 0 chanx_left_out[13]
rlabel metal2 2898 20179 2898 20179 0 chanx_left_out[14]
rlabel metal3 1372 19924 1372 19924 0 chanx_left_out[15]
rlabel via2 3910 20349 3910 20349 0 chanx_left_out[16]
rlabel metal3 1004 20740 1004 20740 0 chanx_left_out[17]
rlabel metal2 2852 21148 2852 21148 0 chanx_left_out[18]
rlabel metal3 1694 21556 1694 21556 0 chanx_left_out[19]
rlabel metal2 2806 13787 2806 13787 0 chanx_left_out[1]
rlabel metal3 2568 21964 2568 21964 0 chanx_left_out[20]
rlabel metal3 1487 22372 1487 22372 0 chanx_left_out[21]
rlabel metal3 1602 22780 1602 22780 0 chanx_left_out[22]
rlabel metal1 9016 20978 9016 20978 0 chanx_left_out[23]
rlabel metal1 3864 17102 3864 17102 0 chanx_left_out[24]
rlabel metal1 4462 16490 4462 16490 0 chanx_left_out[25]
rlabel metal1 4738 18802 4738 18802 0 chanx_left_out[26]
rlabel metal2 3910 23885 3910 23885 0 chanx_left_out[27]
rlabel metal3 4163 16524 4163 16524 0 chanx_left_out[28]
rlabel metal1 9384 19414 9384 19414 0 chanx_left_out[29]
rlabel metal3 1004 14620 1004 14620 0 chanx_left_out[2]
rlabel metal3 1004 15028 1004 15028 0 chanx_left_out[3]
rlabel metal3 1004 15436 1004 15436 0 chanx_left_out[4]
rlabel metal3 1004 15844 1004 15844 0 chanx_left_out[5]
rlabel metal3 1004 16252 1004 16252 0 chanx_left_out[6]
rlabel metal3 1004 16660 1004 16660 0 chanx_left_out[7]
rlabel metal3 958 17068 958 17068 0 chanx_left_out[8]
rlabel metal2 2806 17833 2806 17833 0 chanx_left_out[9]
rlabel via3 22195 22236 22195 22236 0 chany_top_in[0]
rlabel metal1 32522 24140 32522 24140 0 chany_top_in[10]
rlabel metal1 29670 24242 29670 24242 0 chany_top_in[11]
rlabel metal2 30038 25007 30038 25007 0 chany_top_in[12]
rlabel metal1 31050 24174 31050 24174 0 chany_top_in[13]
rlabel metal1 33166 23664 33166 23664 0 chany_top_in[14]
rlabel metal1 32200 23698 32200 23698 0 chany_top_in[15]
rlabel metal1 33810 23732 33810 23732 0 chany_top_in[16]
rlabel metal2 33350 24701 33350 24701 0 chany_top_in[17]
rlabel metal1 33948 24174 33948 24174 0 chany_top_in[18]
rlabel metal1 34776 24174 34776 24174 0 chany_top_in[19]
rlabel metal2 26174 22593 26174 22593 0 chany_top_in[1]
rlabel metal1 35420 24174 35420 24174 0 chany_top_in[20]
rlabel metal1 36248 24174 36248 24174 0 chany_top_in[21]
rlabel metal2 36662 25007 36662 25007 0 chany_top_in[22]
rlabel metal1 37490 24174 37490 24174 0 chany_top_in[23]
rlabel metal1 37812 23698 37812 23698 0 chany_top_in[24]
rlabel metal2 38502 25245 38502 25245 0 chany_top_in[25]
rlabel metal2 39238 25245 39238 25245 0 chany_top_in[26]
rlabel metal2 40066 24531 40066 24531 0 chany_top_in[27]
rlabel metal1 41078 24174 41078 24174 0 chany_top_in[28]
rlabel metal1 41354 23698 41354 23698 0 chany_top_in[29]
rlabel metal2 23506 25510 23506 25510 0 chany_top_in[2]
rlabel metal1 18722 24208 18722 24208 0 chany_top_in[3]
rlabel metal2 24794 24796 24794 24796 0 chany_top_in[4]
rlabel metal1 24748 24174 24748 24174 0 chany_top_in[5]
rlabel metal2 26082 25544 26082 25544 0 chany_top_in[6]
rlabel metal1 27646 24174 27646 24174 0 chany_top_in[7]
rlabel metal1 29578 23766 29578 23766 0 chany_top_in[8]
rlabel metal1 30820 23698 30820 23698 0 chany_top_in[9]
rlabel metal1 3542 23222 3542 23222 0 chany_top_out[0]
rlabel metal1 8786 24242 8786 24242 0 chany_top_out[10]
rlabel metal1 9430 23766 9430 23766 0 chany_top_out[11]
rlabel metal2 10718 24497 10718 24497 0 chany_top_out[12]
rlabel metal1 11454 21998 11454 21998 0 chany_top_out[13]
rlabel metal2 12650 21828 12650 21828 0 chany_top_out[14]
rlabel metal2 12466 25041 12466 25041 0 chany_top_out[15]
rlabel metal2 13301 26316 13301 26316 0 chany_top_out[16]
rlabel metal2 13846 25306 13846 25306 0 chany_top_out[17]
rlabel metal1 13938 24242 13938 24242 0 chany_top_out[18]
rlabel metal1 15410 22134 15410 22134 0 chany_top_out[19]
rlabel metal1 3404 24242 3404 24242 0 chany_top_out[1]
rlabel metal1 15042 23766 15042 23766 0 chany_top_out[20]
rlabel metal2 16146 24497 16146 24497 0 chany_top_out[21]
rlabel metal1 17388 21454 17388 21454 0 chany_top_out[22]
rlabel metal1 16974 23154 16974 23154 0 chany_top_out[23]
rlabel metal1 17250 23630 17250 23630 0 chany_top_out[24]
rlabel metal1 16192 24106 16192 24106 0 chany_top_out[25]
rlabel metal1 18768 23766 18768 23766 0 chany_top_out[26]
rlabel metal1 20562 22066 20562 22066 0 chany_top_out[27]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[28]
rlabel metal1 22494 24310 22494 24310 0 chany_top_out[29]
rlabel metal1 4048 23766 4048 23766 0 chany_top_out[2]
rlabel metal2 5106 24429 5106 24429 0 chany_top_out[3]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[4]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[5]
rlabel metal1 7107 22066 7107 22066 0 chany_top_out[6]
rlabel metal1 6624 24242 6624 24242 0 chany_top_out[7]
rlabel metal2 7866 24735 7866 24735 0 chany_top_out[8]
rlabel metal2 8694 24422 8694 24422 0 chany_top_out[9]
rlabel metal2 19734 17000 19734 17000 0 clknet_0_prog_clk
rlabel metal1 8004 9486 8004 9486 0 clknet_4_0_0_prog_clk
rlabel metal1 22310 11662 22310 11662 0 clknet_4_10_0_prog_clk
rlabel metal2 21942 16388 21942 16388 0 clknet_4_11_0_prog_clk
rlabel metal2 19734 19040 19734 19040 0 clknet_4_12_0_prog_clk
rlabel metal1 18860 23630 18860 23630 0 clknet_4_13_0_prog_clk
rlabel metal1 28106 18292 28106 18292 0 clknet_4_14_0_prog_clk
rlabel metal1 23138 22474 23138 22474 0 clknet_4_15_0_prog_clk
rlabel metal1 8234 12852 8234 12852 0 clknet_4_1_0_prog_clk
rlabel metal1 14950 11186 14950 11186 0 clknet_4_2_0_prog_clk
rlabel metal1 15088 13362 15088 13362 0 clknet_4_3_0_prog_clk
rlabel metal1 5198 20910 5198 20910 0 clknet_4_4_0_prog_clk
rlabel metal1 9614 17714 9614 17714 0 clknet_4_5_0_prog_clk
rlabel metal2 14582 19652 14582 19652 0 clknet_4_6_0_prog_clk
rlabel metal2 13754 19890 13754 19890 0 clknet_4_7_0_prog_clk
rlabel metal2 16882 7616 16882 7616 0 clknet_4_8_0_prog_clk
rlabel metal1 20056 12750 20056 12750 0 clknet_4_9_0_prog_clk
rlabel metal2 4094 1622 4094 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 6762 1622 6762 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 9430 1622 9430 1622 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 12098 1622 12098 1622 0 gfpga_pad_io_soc_dir[3]
rlabel metal2 25438 1588 25438 1588 0 gfpga_pad_io_soc_in[0]
rlabel metal2 28106 823 28106 823 0 gfpga_pad_io_soc_in[1]
rlabel metal2 30774 1588 30774 1588 0 gfpga_pad_io_soc_in[2]
rlabel metal2 33442 1588 33442 1588 0 gfpga_pad_io_soc_in[3]
rlabel metal2 14766 1622 14766 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 17434 1622 17434 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 20102 959 20102 959 0 gfpga_pad_io_soc_out[2]
rlabel metal2 22770 1622 22770 1622 0 gfpga_pad_io_soc_out[3]
rlabel metal2 36110 1588 36110 1588 0 isol_n
rlabel metal1 5474 2278 5474 2278 0 net1
rlabel metal1 12673 17170 12673 17170 0 net10
rlabel metal1 4600 16558 4600 16558 0 net100
rlabel metal1 14306 18802 14306 18802 0 net101
rlabel metal1 6486 18258 6486 18258 0 net102
rlabel metal1 4646 16082 4646 16082 0 net103
rlabel metal1 7774 16150 7774 16150 0 net104
rlabel metal2 13754 17799 13754 17799 0 net105
rlabel metal1 10902 18224 10902 18224 0 net106
rlabel metal2 2530 13362 2530 13362 0 net107
rlabel metal1 2277 16082 2277 16082 0 net108
rlabel metal1 4002 16592 4002 16592 0 net109
rlabel metal2 1886 11747 1886 11747 0 net11
rlabel metal2 3358 17884 3358 17884 0 net110
rlabel metal2 1794 18445 1794 18445 0 net111
rlabel metal1 1886 18258 1886 18258 0 net112
rlabel metal1 2990 14926 2990 14926 0 net113
rlabel metal2 4738 11033 4738 11033 0 net114
rlabel via2 36018 23749 36018 23749 0 net115
rlabel metal2 34270 22797 34270 22797 0 net116
rlabel metal2 35190 24327 35190 24327 0 net117
rlabel metal2 33534 23001 33534 23001 0 net118
rlabel metal2 32522 23171 32522 23171 0 net119
rlabel metal2 7636 12852 7636 12852 0 net12
rlabel metal2 33258 22457 33258 22457 0 net120
rlabel metal2 32062 23392 32062 23392 0 net121
rlabel metal2 34638 24021 34638 24021 0 net122
rlabel metal2 32798 22576 32798 22576 0 net123
rlabel metal1 2346 24174 2346 24174 0 net124
rlabel metal2 31786 24531 31786 24531 0 net125
rlabel metal3 24817 22780 24817 22780 0 net126
rlabel metal1 16928 21522 16928 21522 0 net127
rlabel metal1 16238 23086 16238 23086 0 net128
rlabel metal3 18400 19108 18400 19108 0 net129
rlabel metal1 2254 7752 2254 7752 0 net13
rlabel metal1 14950 24208 14950 24208 0 net130
rlabel metal2 12650 23001 12650 23001 0 net131
rlabel metal2 19090 22202 19090 22202 0 net132
rlabel metal1 19274 18258 19274 18258 0 net133
rlabel metal1 22126 24242 22126 24242 0 net134
rlabel metal2 1150 16898 1150 16898 0 net135
rlabel metal1 4140 22474 4140 22474 0 net136
rlabel metal1 4370 14382 4370 14382 0 net137
rlabel metal2 4048 16388 4048 16388 0 net138
rlabel via2 7038 21981 7038 21981 0 net139
rlabel metal1 2944 3162 2944 3162 0 net14
rlabel via3 9453 9588 9453 9588 0 net140
rlabel metal3 7383 20740 7383 20740 0 net141
rlabel metal3 4600 17340 4600 17340 0 net142
rlabel metal1 4370 2380 4370 2380 0 net143
rlabel metal1 7682 2414 7682 2414 0 net144
rlabel metal1 9706 2414 9706 2414 0 net145
rlabel metal1 12466 2414 12466 2414 0 net146
rlabel metal2 15042 3162 15042 3162 0 net147
rlabel metal1 17204 2822 17204 2822 0 net148
rlabel metal1 19136 2822 19136 2822 0 net149
rlabel metal1 5888 17238 5888 17238 0 net15
rlabel metal1 22356 2414 22356 2414 0 net150
rlabel metal1 21942 21522 21942 21522 0 net151
rlabel metal1 22724 19482 22724 19482 0 net152
rlabel metal2 18814 18292 18814 18292 0 net153
rlabel metal1 23184 20570 23184 20570 0 net154
rlabel metal1 23184 22678 23184 22678 0 net155
rlabel metal1 24564 23698 24564 23698 0 net156
rlabel metal1 26358 21658 26358 21658 0 net157
rlabel metal1 26496 19278 26496 19278 0 net158
rlabel metal1 27554 18258 27554 18258 0 net159
rlabel metal1 5750 15402 5750 15402 0 net16
rlabel metal2 17342 20927 17342 20927 0 net160
rlabel metal1 21298 17306 21298 17306 0 net161
rlabel metal1 24242 18938 24242 18938 0 net162
rlabel metal2 15042 20553 15042 20553 0 net163
rlabel metal2 21114 16932 21114 16932 0 net164
rlabel metal1 14214 8942 14214 8942 0 net165
rlabel metal1 16284 12614 16284 12614 0 net166
rlabel metal2 10258 8058 10258 8058 0 net167
rlabel metal1 11500 7378 11500 7378 0 net168
rlabel metal2 12834 13362 12834 13362 0 net169
rlabel metal2 1610 17307 1610 17307 0 net17
rlabel metal1 15686 8500 15686 8500 0 net170
rlabel metal2 16882 16966 16882 16966 0 net171
rlabel metal2 15410 16524 15410 16524 0 net172
rlabel metal2 14858 16592 14858 16592 0 net173
rlabel metal1 13248 10234 13248 10234 0 net174
rlabel metal2 9614 9350 9614 9350 0 net175
rlabel metal2 11178 12716 11178 12716 0 net176
rlabel metal1 12926 18122 12926 18122 0 net177
rlabel metal2 13202 18394 13202 18394 0 net178
rlabel via2 9338 21301 9338 21301 0 net179
rlabel metal1 2070 10098 2070 10098 0 net18
rlabel metal1 5198 21046 5198 21046 0 net180
rlabel metal2 13386 8262 13386 8262 0 net181
rlabel metal1 2392 11322 2392 11322 0 net182
rlabel metal1 32844 22474 32844 22474 0 net183
rlabel metal2 6992 15028 6992 15028 0 net184
rlabel metal1 7590 11322 7590 11322 0 net185
rlabel metal1 5474 14790 5474 14790 0 net186
rlabel metal1 12926 12648 12926 12648 0 net187
rlabel metal2 17066 11084 17066 11084 0 net188
rlabel metal1 17020 8466 17020 8466 0 net189
rlabel metal2 13478 16439 13478 16439 0 net19
rlabel metal1 9798 10030 9798 10030 0 net190
rlabel metal1 5520 9554 5520 9554 0 net191
rlabel metal1 9154 14926 9154 14926 0 net192
rlabel metal3 14950 16796 14950 16796 0 net193
rlabel metal2 28198 16762 28198 16762 0 net194
rlabel metal2 32154 24310 32154 24310 0 net195
rlabel metal1 14398 20774 14398 20774 0 net196
rlabel metal1 18676 16082 18676 16082 0 net197
rlabel metal1 22034 18292 22034 18292 0 net198
rlabel metal2 48438 22746 48438 22746 0 net2
rlabel metal2 3772 14076 3772 14076 0 net20
rlabel metal1 6118 16082 6118 16082 0 net21
rlabel metal1 1886 8058 1886 8058 0 net22
rlabel metal2 2070 11356 2070 11356 0 net23
rlabel metal2 20194 16371 20194 16371 0 net24
rlabel metal1 1886 2550 1886 2550 0 net25
rlabel metal1 1886 3060 1886 3060 0 net26
rlabel metal2 14766 9180 14766 9180 0 net27
rlabel metal1 13386 8568 13386 8568 0 net28
rlabel metal1 6624 3978 6624 3978 0 net29
rlabel metal1 13570 8364 13570 8364 0 net3
rlabel metal2 12098 6222 12098 6222 0 net30
rlabel metal1 6762 4590 6762 4590 0 net31
rlabel metal2 7406 7123 7406 7123 0 net32
rlabel metal1 15870 13974 15870 13974 0 net33
rlabel metal1 22310 23188 22310 23188 0 net34
rlabel metal2 28106 24497 28106 24497 0 net35
rlabel metal1 11730 20434 11730 20434 0 net36
rlabel metal1 29072 23766 29072 23766 0 net37
rlabel metal2 31786 22508 31786 22508 0 net38
rlabel metal2 27646 23018 27646 23018 0 net39
rlabel metal1 6256 5678 6256 5678 0 net4
rlabel metal2 31050 23120 31050 23120 0 net40
rlabel metal2 33442 24820 33442 24820 0 net41
rlabel metal2 34178 24786 34178 24786 0 net42
rlabel metal2 34546 24888 34546 24888 0 net43
rlabel metal1 28658 21896 28658 21896 0 net44
rlabel metal2 35926 24684 35926 24684 0 net45
rlabel metal1 32522 22032 32522 22032 0 net46
rlabel metal2 35282 22542 35282 22542 0 net47
rlabel metal1 37490 24072 37490 24072 0 net48
rlabel metal2 37766 20944 37766 20944 0 net49
rlabel metal1 6808 6222 6808 6222 0 net5
rlabel metal2 38686 24548 38686 24548 0 net50
rlabel metal2 39330 24718 39330 24718 0 net51
rlabel metal1 39330 24208 39330 24208 0 net52
rlabel metal2 38686 22457 38686 22457 0 net53
rlabel metal2 41354 21624 41354 21624 0 net54
rlabel metal2 18814 24412 18814 24412 0 net55
rlabel metal1 15686 21012 15686 21012 0 net56
rlabel metal1 19504 23290 19504 23290 0 net57
rlabel metal1 23874 24072 23874 24072 0 net58
rlabel metal1 27002 23120 27002 23120 0 net59
rlabel metal1 2507 6630 2507 6630 0 net6
rlabel metal1 27002 22950 27002 22950 0 net60
rlabel metal1 25990 22746 25990 22746 0 net61
rlabel metal1 30958 23494 30958 23494 0 net62
rlabel metal2 25530 4114 25530 4114 0 net63
rlabel metal1 28014 2618 28014 2618 0 net64
rlabel metal1 29900 2618 29900 2618 0 net65
rlabel metal2 33534 3842 33534 3842 0 net66
rlabel metal1 25254 6766 25254 6766 0 net67
rlabel metal1 39751 22678 39751 22678 0 net68
rlabel metal2 45402 21454 45402 21454 0 net69
rlabel metal2 8418 8296 8418 8296 0 net7
rlabel metal2 34454 21284 34454 21284 0 net70
rlabel metal2 28428 23460 28428 23460 0 net71
rlabel metal2 46966 22729 46966 22729 0 net72
rlabel metal2 46414 20774 46414 20774 0 net73
rlabel metal2 48806 20621 48806 20621 0 net74
rlabel metal1 39859 23562 39859 23562 0 net75
rlabel metal2 37214 20145 37214 20145 0 net76
rlabel metal2 49266 17850 49266 17850 0 net77
rlabel metal2 42826 20264 42826 20264 0 net78
rlabel metal2 48714 22457 48714 22457 0 net79
rlabel metal1 7774 15470 7774 15470 0 net8
rlabel metal2 48530 21080 48530 21080 0 net80
rlabel metal1 47932 21522 47932 21522 0 net81
rlabel metal2 7268 20468 7268 20468 0 net82
rlabel via2 1794 12835 1794 12835 0 net83
rlabel metal1 1794 18768 1794 18768 0 net84
rlabel metal1 1794 19380 1794 19380 0 net85
rlabel metal2 1794 20740 1794 20740 0 net86
rlabel metal1 1840 20434 1840 20434 0 net87
rlabel metal2 4370 19380 4370 19380 0 net88
rlabel metal2 2346 19380 2346 19380 0 net89
rlabel metal1 1656 6630 1656 6630 0 net9
rlabel metal1 3634 20468 3634 20468 0 net90
rlabel metal1 2024 21998 2024 21998 0 net91
rlabel metal2 1702 22950 1702 22950 0 net92
rlabel metal2 1794 22882 1794 22882 0 net93
rlabel metal2 19918 18377 19918 18377 0 net94
rlabel metal2 2346 22780 2346 22780 0 net95
rlabel metal1 4508 19346 4508 19346 0 net96
rlabel metal1 6716 22202 6716 22202 0 net97
rlabel metal2 14950 21726 14950 21726 0 net98
rlabel metal2 3450 14756 3450 14756 0 net99
rlabel metal2 38778 2098 38778 2098 0 prog_clk
rlabel metal1 42136 24174 42136 24174 0 prog_reset_top_in
rlabel metal1 19412 17102 19412 17102 0 sb_8__0_.mem_left_track_1.ccff_head
rlabel metal2 25346 19244 25346 19244 0 sb_8__0_.mem_left_track_1.ccff_tail
rlabel metal1 30038 16626 30038 16626 0 sb_8__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 18078 21862 18078 21862 0 sb_8__0_.mem_left_track_11.ccff_head
rlabel metal1 16376 23018 16376 23018 0 sb_8__0_.mem_left_track_11.ccff_tail
rlabel metal1 22218 24820 22218 24820 0 sb_8__0_.mem_left_track_11.mem_out\[0\]
rlabel metal2 20010 21461 20010 21461 0 sb_8__0_.mem_left_track_13.ccff_tail
rlabel metal2 25898 24514 25898 24514 0 sb_8__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 18860 20366 18860 20366 0 sb_8__0_.mem_left_track_15.ccff_tail
rlabel metal2 25162 22950 25162 22950 0 sb_8__0_.mem_left_track_15.mem_out\[0\]
rlabel via1 23414 22525 23414 22525 0 sb_8__0_.mem_left_track_17.ccff_tail
rlabel metal2 23782 23358 23782 23358 0 sb_8__0_.mem_left_track_17.mem_out\[0\]
rlabel metal1 23920 21454 23920 21454 0 sb_8__0_.mem_left_track_19.ccff_tail
rlabel metal1 24426 22406 24426 22406 0 sb_8__0_.mem_left_track_19.mem_out\[0\]
rlabel metal2 26174 19482 26174 19482 0 sb_8__0_.mem_left_track_29.ccff_tail
rlabel metal1 26910 20298 26910 20298 0 sb_8__0_.mem_left_track_29.mem_out\[0\]
rlabel metal1 17940 19890 17940 19890 0 sb_8__0_.mem_left_track_3.ccff_tail
rlabel metal1 19918 19278 19918 19278 0 sb_8__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 26036 21930 26036 21930 0 sb_8__0_.mem_left_track_31.ccff_tail
rlabel metal1 27738 20026 27738 20026 0 sb_8__0_.mem_left_track_31.mem_out\[0\]
rlabel metal1 24702 22134 24702 22134 0 sb_8__0_.mem_left_track_33.ccff_tail
rlabel metal2 25898 23460 25898 23460 0 sb_8__0_.mem_left_track_33.mem_out\[0\]
rlabel metal2 25254 24480 25254 24480 0 sb_8__0_.mem_left_track_35.ccff_tail
rlabel metal1 28842 23494 28842 23494 0 sb_8__0_.mem_left_track_35.mem_out\[0\]
rlabel metal1 29578 22406 29578 22406 0 sb_8__0_.mem_left_track_45.ccff_tail
rlabel metal1 31142 22134 31142 22134 0 sb_8__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 28566 19278 28566 19278 0 sb_8__0_.mem_left_track_47.ccff_tail
rlabel metal2 30222 20842 30222 20842 0 sb_8__0_.mem_left_track_47.mem_out\[0\]
rlabel metal1 27876 18802 27876 18802 0 sb_8__0_.mem_left_track_49.ccff_tail
rlabel metal2 30130 18666 30130 18666 0 sb_8__0_.mem_left_track_49.mem_out\[0\]
rlabel metal2 20562 20060 20562 20060 0 sb_8__0_.mem_left_track_5.ccff_tail
rlabel metal1 20516 21386 20516 21386 0 sb_8__0_.mem_left_track_5.mem_out\[0\]
rlabel metal2 30866 17884 30866 17884 0 sb_8__0_.mem_left_track_51.mem_out\[0\]
rlabel metal2 20010 19652 20010 19652 0 sb_8__0_.mem_left_track_7.ccff_tail
rlabel metal1 21804 19958 21804 19958 0 sb_8__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 17480 21930 17480 21930 0 sb_8__0_.mem_left_track_9.mem_out\[0\]
rlabel metal1 25070 15062 25070 15062 0 sb_8__0_.mem_top_track_0.ccff_tail
rlabel metal2 39698 22270 39698 22270 0 sb_8__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 27784 16626 27784 16626 0 sb_8__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 20838 13804 20838 13804 0 sb_8__0_.mem_top_track_10.ccff_head
rlabel metal2 17434 10812 17434 10812 0 sb_8__0_.mem_top_track_10.ccff_tail
rlabel metal2 24058 11968 24058 11968 0 sb_8__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 21436 12750 21436 12750 0 sb_8__0_.mem_top_track_10.mem_out\[1\]
rlabel metal2 16330 9724 16330 9724 0 sb_8__0_.mem_top_track_12.ccff_tail
rlabel metal2 19228 13430 19228 13430 0 sb_8__0_.mem_top_track_12.mem_out\[0\]
rlabel metal2 14858 11186 14858 11186 0 sb_8__0_.mem_top_track_14.ccff_tail
rlabel metal1 14214 9486 14214 9486 0 sb_8__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 13294 12716 13294 12716 0 sb_8__0_.mem_top_track_16.ccff_tail
rlabel metal1 16974 10234 16974 10234 0 sb_8__0_.mem_top_track_16.mem_out\[0\]
rlabel metal2 17434 13736 17434 13736 0 sb_8__0_.mem_top_track_18.ccff_tail
rlabel metal1 17434 13192 17434 13192 0 sb_8__0_.mem_top_track_18.mem_out\[0\]
rlabel metal2 21206 9690 21206 9690 0 sb_8__0_.mem_top_track_2.ccff_tail
rlabel metal1 23920 14450 23920 14450 0 sb_8__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 24656 11866 24656 11866 0 sb_8__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 18078 15334 18078 15334 0 sb_8__0_.mem_top_track_20.ccff_tail
rlabel metal1 17940 15538 17940 15538 0 sb_8__0_.mem_top_track_20.mem_out\[0\]
rlabel metal1 15916 14926 15916 14926 0 sb_8__0_.mem_top_track_22.ccff_tail
rlabel metal1 15088 14926 15088 14926 0 sb_8__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 15870 13430 15870 13430 0 sb_8__0_.mem_top_track_24.ccff_tail
rlabel metal1 15134 13838 15134 13838 0 sb_8__0_.mem_top_track_24.mem_out\[0\]
rlabel metal1 12558 11628 12558 11628 0 sb_8__0_.mem_top_track_26.ccff_tail
rlabel metal1 12180 10438 12180 10438 0 sb_8__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 12052 11186 12052 11186 0 sb_8__0_.mem_top_track_28.ccff_tail
rlabel metal2 13202 9758 13202 9758 0 sb_8__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 13478 13974 13478 13974 0 sb_8__0_.mem_top_track_30.ccff_tail
rlabel metal1 12328 13226 12328 13226 0 sb_8__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 13064 18190 13064 18190 0 sb_8__0_.mem_top_track_32.ccff_tail
rlabel metal2 13570 15470 13570 15470 0 sb_8__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 11362 18802 11362 18802 0 sb_8__0_.mem_top_track_34.ccff_tail
rlabel metal1 13708 17782 13708 17782 0 sb_8__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 10120 20230 10120 20230 0 sb_8__0_.mem_top_track_36.ccff_tail
rlabel metal2 12558 19924 12558 19924 0 sb_8__0_.mem_top_track_36.mem_out\[0\]
rlabel metal1 5152 18666 5152 18666 0 sb_8__0_.mem_top_track_38.ccff_tail
rlabel metal1 7866 16048 7866 16048 0 sb_8__0_.mem_top_track_38.mem_out\[0\]
rlabel metal2 18952 12750 18952 12750 0 sb_8__0_.mem_top_track_4.ccff_tail
rlabel metal2 22678 10880 22678 10880 0 sb_8__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 18722 12750 18722 12750 0 sb_8__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 7084 21590 7084 21590 0 sb_8__0_.mem_top_track_40.ccff_tail
rlabel metal1 4830 19720 4830 19720 0 sb_8__0_.mem_top_track_40.mem_out\[0\]
rlabel metal2 10994 22542 10994 22542 0 sb_8__0_.mem_top_track_42.ccff_tail
rlabel metal1 12466 21420 12466 21420 0 sb_8__0_.mem_top_track_42.mem_out\[0\]
rlabel metal1 13294 21454 13294 21454 0 sb_8__0_.mem_top_track_44.ccff_tail
rlabel metal2 12650 18632 12650 18632 0 sb_8__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 15180 19890 15180 19890 0 sb_8__0_.mem_top_track_46.ccff_tail
rlabel metal1 14076 20366 14076 20366 0 sb_8__0_.mem_top_track_46.mem_out\[0\]
rlabel metal1 16652 17714 16652 17714 0 sb_8__0_.mem_top_track_48.ccff_tail
rlabel metal1 15870 20026 15870 20026 0 sb_8__0_.mem_top_track_48.mem_out\[0\]
rlabel metal2 18446 16898 18446 16898 0 sb_8__0_.mem_top_track_50.mem_out\[0\]
rlabel metal2 21482 14824 21482 14824 0 sb_8__0_.mem_top_track_6.ccff_tail
rlabel metal1 22395 14790 22395 14790 0 sb_8__0_.mem_top_track_6.mem_out\[0\]
rlabel metal2 20010 14535 20010 14535 0 sb_8__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 24012 14246 24012 14246 0 sb_8__0_.mem_top_track_8.mem_out\[0\]
rlabel metal2 22034 12687 22034 12687 0 sb_8__0_.mem_top_track_8.mem_out\[1\]
rlabel via2 12466 18411 12466 18411 0 sb_8__0_.mux_left_track_1.out
rlabel metal1 26358 19686 26358 19686 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27830 16456 27830 16456 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22770 18721 22770 18721 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 3818 12206 3818 12206 0 sb_8__0_.mux_left_track_11.out
rlabel metal2 25806 24480 25806 24480 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 1840 17850 1840 17850 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 18952 17884 18952 17884 0 sb_8__0_.mux_left_track_13.out
rlabel metal2 27186 24089 27186 24089 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17894 20519 17894 20519 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 16652 15912 16652 15912 0 sb_8__0_.mux_left_track_15.out
rlabel metal1 18814 20502 18814 20502 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20286 14994 20286 14994 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19642 13770 19642 13770 0 sb_8__0_.mux_left_track_17.out
rlabel metal2 18630 21335 18630 21335 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19872 13906 19872 13906 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16146 14620 16146 14620 0 sb_8__0_.mux_left_track_19.out
rlabel metal2 22494 21420 22494 21420 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20148 14382 20148 14382 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8188 15130 8188 15130 0 sb_8__0_.mux_left_track_29.out
rlabel metal1 23276 19482 23276 19482 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9798 13345 9798 13345 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9246 13923 9246 13923 0 sb_8__0_.mux_left_track_3.out
rlabel metal1 17296 19890 17296 19890 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16974 19992 16974 19992 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16146 15776 16146 15776 0 sb_8__0_.mux_left_track_31.out
rlabel metal1 25438 20570 25438 20570 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20746 18377 20746 18377 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 5198 10115 5198 10115 0 sb_8__0_.mux_left_track_33.out
rlabel metal1 25346 22678 25346 22678 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23414 11152 23414 11152 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 6670 17204 6670 17204 0 sb_8__0_.mux_left_track_35.out
rlabel metal2 25070 23936 25070 23936 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23874 22508 23874 22508 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4554 18734 4554 18734 0 sb_8__0_.mux_left_track_45.out
rlabel metal1 29578 21862 29578 21862 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 25622 21403 25622 21403 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10028 16558 10028 16558 0 sb_8__0_.mux_left_track_47.out
rlabel metal1 25162 21012 25162 21012 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21942 22474 21942 22474 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 6670 14756 6670 14756 0 sb_8__0_.mux_left_track_49.out
rlabel metal1 29210 18666 29210 18666 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17894 16252 17894 16252 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13478 21624 13478 21624 0 sb_8__0_.mux_left_track_5.out
rlabel metal1 21298 20468 21298 20468 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17158 20230 17158 20230 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6256 12818 6256 12818 0 sb_8__0_.mux_left_track_51.out
rlabel metal1 21643 17238 21643 17238 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19458 17000 19458 17000 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14674 19550 14674 19550 0 sb_8__0_.mux_left_track_7.out
rlabel metal1 19182 19346 19182 19346 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18722 19346 18722 19346 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14490 18836 14490 18836 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9844 8466 9844 8466 0 sb_8__0_.mux_left_track_9.out
rlabel metal2 15226 21114 15226 21114 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15502 21080 15502 21080 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel via1 21942 24157 21942 24157 0 sb_8__0_.mux_top_track_0.out
rlabel metal2 27094 17748 27094 17748 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27324 16558 27324 16558 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26036 16422 26036 16422 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21068 15878 21068 15878 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23598 19006 23598 19006 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18630 16014 18630 16014 0 sb_8__0_.mux_top_track_10.out
rlabel metal1 21206 12716 21206 12716 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21114 13464 21114 13464 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20746 12517 20746 12517 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15134 8806 15134 8806 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15410 17646 15410 17646 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 28566 16201 28566 16201 0 sb_8__0_.mux_top_track_12.out
rlabel metal1 20102 14246 20102 14246 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14306 9486 14306 9486 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19504 13294 19504 13294 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 16192 14348 16192 14348 0 sb_8__0_.mux_top_track_14.out
rlabel metal1 16928 11594 16928 11594 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13478 8330 13478 8330 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15824 17646 15824 17646 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 10258 15589 10258 15589 0 sb_8__0_.mux_top_track_16.out
rlabel metal1 18032 11866 18032 11866 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12729 12920 12729 12920 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 10994 14212 10994 14212 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32384 20842 32384 20842 0 sb_8__0_.mux_top_track_18.out
rlabel metal1 19366 16218 19366 16218 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13202 13804 13202 13804 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16698 14586 16698 14586 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18952 17850 18952 17850 0 sb_8__0_.mux_top_track_2.out
rlabel metal1 24978 13974 24978 13974 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25392 14042 25392 14042 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21574 9622 21574 9622 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 13110 8738 13110 8738 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19366 9418 19366 9418 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 32706 19023 32706 19023 0 sb_8__0_.mux_top_track_20.out
rlabel metal1 16008 15606 16008 15606 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15962 16864 15962 16864 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34224 23698 34224 23698 0 sb_8__0_.mux_top_track_22.out
rlabel metal1 15134 15606 15134 15606 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19504 15470 19504 15470 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32338 21522 32338 21522 0 sb_8__0_.mux_top_track_24.out
rlabel metal1 14398 13804 14398 13804 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 3450 13940 3450 13940 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33258 22610 33258 22610 0 sb_8__0_.mux_top_track_26.out
rlabel metal1 11132 11322 11132 11322 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12006 12036 12006 12036 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32430 17187 32430 17187 0 sb_8__0_.mux_top_track_28.out
rlabel metal2 10350 10132 10350 10132 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8786 10778 8786 10778 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 30452 22950 30452 22950 0 sb_8__0_.mux_top_track_30.out
rlabel metal1 11914 12410 11914 12410 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12098 15895 12098 15895 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 35098 21590 35098 21590 0 sb_8__0_.mux_top_track_32.out
rlabel metal1 12926 15130 12926 15130 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12098 18105 12098 18105 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33626 21658 33626 21658 0 sb_8__0_.mux_top_track_34.out
rlabel metal2 11914 17952 11914 17952 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 33442 20111 33442 20111 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 35834 19040 35834 19040 0 sb_8__0_.mux_top_track_36.out
rlabel metal2 12098 20230 12098 20230 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 3128 14212 3128 14212 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5382 9078 5382 9078 0 sb_8__0_.mux_top_track_38.out
rlabel metal1 7452 16218 7452 16218 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 4255 20740 4255 20740 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18584 16422 18584 16422 0 sb_8__0_.mux_top_track_4.out
rlabel metal1 19596 12818 19596 12818 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21206 12886 21206 12886 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17020 12954 17020 12954 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16100 13906 16100 13906 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16974 14042 16974 14042 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 5152 8602 5152 8602 0 sb_8__0_.mux_top_track_40.out
rlabel metal1 7958 17306 7958 17306 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 6417 19380 6417 19380 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7498 8364 7498 8364 0 sb_8__0_.mux_top_track_42.out
rlabel metal2 11914 21794 11914 21794 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9154 21862 9154 21862 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 34362 15929 34362 15929 0 sb_8__0_.mux_top_track_44.out
rlabel metal1 17572 18870 17572 18870 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8050 17782 8050 17782 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 33534 21471 33534 21471 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 24886 9673 24886 9673 0 sb_8__0_.mux_top_track_46.out
rlabel metal1 14812 19686 14812 19686 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12926 18428 12926 18428 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32614 20893 32614 20893 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 29992 19822 29992 19822 0 sb_8__0_.mux_top_track_48.out
rlabel metal1 17664 18394 17664 18394 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13570 17374 13570 17374 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15134 18343 15134 18343 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 31326 14977 31326 14977 0 sb_8__0_.mux_top_track_50.out
rlabel metal1 19550 17782 19550 17782 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13018 16626 13018 16626 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16882 19261 16882 19261 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9200 15470 9200 15470 0 sb_8__0_.mux_top_track_6.out
rlabel metal1 22310 15538 22310 15538 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22632 15470 22632 15470 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20746 15062 20746 15062 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 13846 13872 13846 13872 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18216 15130 18216 15130 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18722 17544 18722 17544 0 sb_8__0_.mux_top_track_8.out
rlabel metal1 23368 13362 23368 13362 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23690 13226 23690 13226 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21390 13702 21390 13702 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16146 12750 16146 12750 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19734 14042 19734 14042 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 44988 24174 44988 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal2 45494 25296 45494 25296 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 46368 24174 46368 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 46736 23698 46736 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 47564 24174 47564 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 48254 24174 48254 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal2 43654 25041 43654 25041 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 44252 23698 44252 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel via2 49082 21981 49082 21981 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 49082 23001 49082 23001 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 49082 23783 49082 23783 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 48346 24259 48346 24259 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 41446 2234 41446 2234 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 44114 2200 44114 2200 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 26128 23086 26128 23086 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 25622 22610 25622 22610 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
