magic
tech sky130A
magscale 1 2
timestamp 1680198063
<< viali >>
rect 14565 54281 14599 54315
rect 16405 54281 16439 54315
rect 24501 54281 24535 54315
rect 5825 54213 5859 54247
rect 8401 54213 8435 54247
rect 10977 54213 11011 54247
rect 14105 54213 14139 54247
rect 18429 54213 18463 54247
rect 21465 54213 21499 54247
rect 23305 54213 23339 54247
rect 2237 54145 2271 54179
rect 4629 54145 4663 54179
rect 7389 54145 7423 54179
rect 9965 54145 9999 54179
rect 11897 54145 11931 54179
rect 12357 54145 12391 54179
rect 14841 54145 14875 54179
rect 15577 54145 15611 54179
rect 16129 54145 16163 54179
rect 16865 54145 16899 54179
rect 17601 54145 17635 54179
rect 18981 54145 19015 54179
rect 19441 54145 19475 54179
rect 20177 54145 20211 54179
rect 20913 54145 20947 54179
rect 22017 54145 22051 54179
rect 22753 54145 22787 54179
rect 23765 54145 23799 54179
rect 24961 54145 24995 54179
rect 3249 54077 3283 54111
rect 12817 54077 12851 54111
rect 17785 54009 17819 54043
rect 25145 54009 25179 54043
rect 11713 53941 11747 53975
rect 15025 53941 15059 53975
rect 15761 53941 15795 53975
rect 17049 53941 17083 53975
rect 18521 53941 18555 53975
rect 19625 53941 19659 53975
rect 20361 53941 20395 53975
rect 21097 53941 21131 53975
rect 22201 53941 22235 53975
rect 22937 53941 22971 53975
rect 23949 53941 23983 53975
rect 16405 53737 16439 53771
rect 18889 53737 18923 53771
rect 21281 53669 21315 53703
rect 23121 53669 23155 53703
rect 3249 53601 3283 53635
rect 6561 53601 6595 53635
rect 8401 53601 8435 53635
rect 11069 53601 11103 53635
rect 12725 53601 12759 53635
rect 24409 53601 24443 53635
rect 2237 53533 2271 53567
rect 5549 53533 5583 53567
rect 7297 53533 7331 53567
rect 10425 53533 10459 53567
rect 12449 53533 12483 53567
rect 14289 53533 14323 53567
rect 14841 53533 14875 53567
rect 15669 53533 15703 53567
rect 16129 53533 16163 53567
rect 16681 53533 16715 53567
rect 17601 53533 17635 53567
rect 18245 53533 18279 53567
rect 18705 53533 18739 53567
rect 19441 53533 19475 53567
rect 20269 53533 20303 53567
rect 20729 53533 20763 53567
rect 21097 53533 21131 53567
rect 22017 53533 22051 53567
rect 22661 53533 22695 53567
rect 23305 53533 23339 53567
rect 23857 53533 23891 53567
rect 24593 53533 24627 53567
rect 25053 53533 25087 53567
rect 15853 53465 15887 53499
rect 20453 53465 20487 53499
rect 24041 53465 24075 53499
rect 14473 53397 14507 53431
rect 16865 53397 16899 53431
rect 17417 53397 17451 53431
rect 18337 53397 18371 53431
rect 19625 53397 19659 53431
rect 21833 53397 21867 53431
rect 22477 53397 22511 53431
rect 25237 53397 25271 53431
rect 2145 53193 2179 53227
rect 17325 53193 17359 53227
rect 19533 53193 19567 53227
rect 19717 53193 19751 53227
rect 21005 53193 21039 53227
rect 21833 53193 21867 53227
rect 22293 53193 22327 53227
rect 22569 53193 22603 53227
rect 23029 53193 23063 53227
rect 3985 53125 4019 53159
rect 5825 53125 5859 53159
rect 9137 53125 9171 53159
rect 13829 53125 13863 53159
rect 21189 53125 21223 53159
rect 1777 53057 1811 53091
rect 2973 53057 3007 53091
rect 4813 53057 4847 53091
rect 8125 53057 8159 53091
rect 9781 53057 9815 53091
rect 11897 53057 11931 53091
rect 14657 53057 14691 53091
rect 14933 53057 14967 53091
rect 16129 53057 16163 53091
rect 16405 53057 16439 53091
rect 19073 53057 19107 53091
rect 19349 53057 19383 53091
rect 20545 53057 20579 53091
rect 20821 53057 20855 53091
rect 23489 53057 23523 53091
rect 24133 53057 24167 53091
rect 24409 53057 24443 53091
rect 24777 53057 24811 53091
rect 25053 53057 25087 53091
rect 10333 52989 10367 53023
rect 12357 52989 12391 53023
rect 1593 52921 1627 52955
rect 14013 52921 14047 52955
rect 14473 52853 14507 52887
rect 15945 52853 15979 52887
rect 18889 52853 18923 52887
rect 20361 52853 20395 52887
rect 23305 52853 23339 52887
rect 23949 52853 23983 52887
rect 25237 52853 25271 52887
rect 12633 52649 12667 52683
rect 14105 52649 14139 52683
rect 24593 52649 24627 52683
rect 25237 52581 25271 52615
rect 3249 52513 3283 52547
rect 3985 52513 4019 52547
rect 4261 52513 4295 52547
rect 7757 52513 7791 52547
rect 11253 52513 11287 52547
rect 2237 52445 2271 52479
rect 5457 52445 5491 52479
rect 6561 52445 6595 52479
rect 7297 52445 7331 52479
rect 10793 52445 10827 52479
rect 12817 52445 12851 52479
rect 13645 52445 13679 52479
rect 24777 52445 24811 52479
rect 25053 52445 25087 52479
rect 13461 52377 13495 52411
rect 7021 52105 7055 52139
rect 11713 52105 11747 52139
rect 12357 52105 12391 52139
rect 13277 52105 13311 52139
rect 25237 52105 25271 52139
rect 6929 52037 6963 52071
rect 2973 51969 3007 52003
rect 4721 51969 4755 52003
rect 8033 51969 8067 52003
rect 9781 51969 9815 52003
rect 11897 51969 11931 52003
rect 12541 51969 12575 52003
rect 3341 51901 3375 51935
rect 5089 51901 5123 51935
rect 8493 51901 8527 51935
rect 10149 51901 10183 51935
rect 25513 51765 25547 51799
rect 3801 51561 3835 51595
rect 10241 51561 10275 51595
rect 2881 51425 2915 51459
rect 5733 51425 5767 51459
rect 7573 51425 7607 51459
rect 2237 51357 2271 51391
rect 5457 51357 5491 51391
rect 7113 51357 7147 51391
rect 10425 51357 10459 51391
rect 25053 51357 25087 51391
rect 25237 51221 25271 51255
rect 6929 51017 6963 51051
rect 9597 50949 9631 50983
rect 2513 50881 2547 50915
rect 4169 50881 4203 50915
rect 6837 50881 6871 50915
rect 7757 50881 7791 50915
rect 9413 50881 9447 50915
rect 24777 50881 24811 50915
rect 25053 50881 25087 50915
rect 2789 50813 2823 50847
rect 4629 50813 4663 50847
rect 7481 50813 7515 50847
rect 25237 50677 25271 50711
rect 6837 50473 6871 50507
rect 9229 50473 9263 50507
rect 3985 50337 4019 50371
rect 5089 50337 5123 50371
rect 2237 50269 2271 50303
rect 3249 50269 3283 50303
rect 4261 50269 4295 50303
rect 7021 50269 7055 50303
rect 9413 50269 9447 50303
rect 25421 50133 25455 50167
rect 25145 49929 25179 49963
rect 3157 49861 3191 49895
rect 6009 49861 6043 49895
rect 9321 49861 9355 49895
rect 2145 49793 2179 49827
rect 3985 49793 4019 49827
rect 6377 49793 6411 49827
rect 9137 49793 9171 49827
rect 25329 49793 25363 49827
rect 4242 49589 4276 49623
rect 11621 49385 11655 49419
rect 2053 49249 2087 49283
rect 1777 49181 1811 49215
rect 11805 49181 11839 49215
rect 24869 49181 24903 49215
rect 25329 49181 25363 49215
rect 25145 49045 25179 49079
rect 12725 48841 12759 48875
rect 12909 48705 12943 48739
rect 25513 48501 25547 48535
rect 17785 48229 17819 48263
rect 24869 48093 24903 48127
rect 25329 48093 25363 48127
rect 1685 48025 1719 48059
rect 1869 48025 1903 48059
rect 2145 47957 2179 47991
rect 25145 47957 25179 47991
rect 9137 47753 9171 47787
rect 17233 47753 17267 47787
rect 17325 47753 17359 47787
rect 18429 47753 18463 47787
rect 18521 47685 18555 47719
rect 19073 47685 19107 47719
rect 9321 47617 9355 47651
rect 24501 47617 24535 47651
rect 17417 47549 17451 47583
rect 18705 47549 18739 47583
rect 24777 47549 24811 47583
rect 16865 47413 16899 47447
rect 18061 47413 18095 47447
rect 15932 47209 15966 47243
rect 19349 47209 19383 47243
rect 21649 47209 21683 47243
rect 18153 47141 18187 47175
rect 25145 47141 25179 47175
rect 10241 47073 10275 47107
rect 15669 47073 15703 47107
rect 17417 47073 17451 47107
rect 18613 47073 18647 47107
rect 18797 47073 18831 47107
rect 22477 47073 22511 47107
rect 22569 47073 22603 47107
rect 18521 47005 18555 47039
rect 22385 47005 22419 47039
rect 25329 47005 25363 47039
rect 10517 46937 10551 46971
rect 24869 46937 24903 46971
rect 11989 46869 12023 46903
rect 12357 46869 12391 46903
rect 14197 46869 14231 46903
rect 17693 46869 17727 46903
rect 22017 46869 22051 46903
rect 7205 46665 7239 46699
rect 10885 46665 10919 46699
rect 18613 46665 18647 46699
rect 20821 46665 20855 46699
rect 22017 46665 22051 46699
rect 22661 46665 22695 46699
rect 22753 46665 22787 46699
rect 12633 46597 12667 46631
rect 21097 46597 21131 46631
rect 7389 46529 7423 46563
rect 11069 46529 11103 46563
rect 12357 46461 12391 46495
rect 14565 46461 14599 46495
rect 14841 46461 14875 46495
rect 16865 46461 16899 46495
rect 17141 46461 17175 46495
rect 19073 46461 19107 46495
rect 19349 46461 19383 46495
rect 22845 46461 22879 46495
rect 24501 46461 24535 46495
rect 24777 46461 24811 46495
rect 14105 46325 14139 46359
rect 16313 46325 16347 46359
rect 22293 46325 22327 46359
rect 8125 46121 8159 46155
rect 9137 46121 9171 46155
rect 10701 46121 10735 46155
rect 25421 46121 25455 46155
rect 10057 46053 10091 46087
rect 1869 45985 1903 46019
rect 11345 45985 11379 46019
rect 11897 45985 11931 46019
rect 12173 45985 12207 46019
rect 20177 45985 20211 46019
rect 20361 45985 20395 46019
rect 21373 45985 21407 46019
rect 21557 45985 21591 46019
rect 1593 45917 1627 45951
rect 9321 45917 9355 45951
rect 10241 45917 10275 45951
rect 21281 45917 21315 45951
rect 23213 45917 23247 45951
rect 23489 45917 23523 45951
rect 8033 45849 8067 45883
rect 8493 45849 8527 45883
rect 11069 45849 11103 45883
rect 20085 45849 20119 45883
rect 11161 45781 11195 45815
rect 13645 45781 13679 45815
rect 14197 45781 14231 45815
rect 16405 45781 16439 45815
rect 18705 45781 18739 45815
rect 19349 45781 19383 45815
rect 19717 45781 19751 45815
rect 20913 45781 20947 45815
rect 24501 45781 24535 45815
rect 1409 45577 1443 45611
rect 20177 45577 20211 45611
rect 23765 45577 23799 45611
rect 9505 45509 9539 45543
rect 16405 45509 16439 45543
rect 24777 45441 24811 45475
rect 9229 45373 9263 45407
rect 14381 45373 14415 45407
rect 14657 45373 14691 45407
rect 18429 45373 18463 45407
rect 18705 45373 18739 45407
rect 22017 45373 22051 45407
rect 22293 45373 22327 45407
rect 24501 45373 24535 45407
rect 10977 45305 11011 45339
rect 8861 45237 8895 45271
rect 11253 45237 11287 45271
rect 12173 45237 12207 45271
rect 16129 45237 16163 45271
rect 20545 45237 20579 45271
rect 20821 45237 20855 45271
rect 24041 45237 24075 45271
rect 7849 45033 7883 45067
rect 11621 45033 11655 45067
rect 13001 45033 13035 45067
rect 17141 45033 17175 45067
rect 9413 44965 9447 44999
rect 12541 44897 12575 44931
rect 13553 44897 13587 44931
rect 21649 44897 21683 44931
rect 12357 44829 12391 44863
rect 13369 44829 13403 44863
rect 15117 44829 15151 44863
rect 19533 44829 19567 44863
rect 22293 44829 22327 44863
rect 24501 44829 24535 44863
rect 7757 44761 7791 44795
rect 8217 44761 8251 44795
rect 9229 44761 9263 44795
rect 11161 44761 11195 44795
rect 11529 44761 11563 44795
rect 15393 44761 15427 44795
rect 19809 44761 19843 44795
rect 22569 44761 22603 44795
rect 6469 44693 6503 44727
rect 7205 44693 7239 44727
rect 9689 44693 9723 44727
rect 13461 44693 13495 44727
rect 16865 44693 16899 44727
rect 21281 44693 21315 44727
rect 24041 44693 24075 44727
rect 25513 44693 25547 44727
rect 5825 44489 5859 44523
rect 6745 44489 6779 44523
rect 7481 44489 7515 44523
rect 8033 44489 8067 44523
rect 11069 44489 11103 44523
rect 11897 44489 11931 44523
rect 12265 44489 12299 44523
rect 18889 44489 18923 44523
rect 21281 44489 21315 44523
rect 21557 44489 21591 44523
rect 24041 44489 24075 44523
rect 9137 44421 9171 44455
rect 6009 44353 6043 44387
rect 6653 44353 6687 44387
rect 7389 44353 7423 44387
rect 8217 44353 8251 44387
rect 8953 44353 8987 44387
rect 9413 44353 9447 44387
rect 10977 44353 11011 44387
rect 13185 44353 13219 44387
rect 24501 44353 24535 44387
rect 12357 44285 12391 44319
rect 12449 44285 12483 44319
rect 14933 44285 14967 44319
rect 16865 44285 16899 44319
rect 17141 44285 17175 44319
rect 19533 44285 19567 44319
rect 19809 44285 19843 44319
rect 22293 44285 22327 44319
rect 22569 44285 22603 44319
rect 24777 44285 24811 44319
rect 11529 44149 11563 44183
rect 13448 44149 13482 44183
rect 15209 44149 15243 44183
rect 18613 44149 18647 44183
rect 6837 43945 6871 43979
rect 8401 43945 8435 43979
rect 11621 43945 11655 43979
rect 9413 43809 9447 43843
rect 22477 43809 22511 43843
rect 22661 43809 22695 43843
rect 8585 43741 8619 43775
rect 9137 43741 9171 43775
rect 6745 43673 6779 43707
rect 7205 43673 7239 43707
rect 11529 43673 11563 43707
rect 11989 43673 12023 43707
rect 22385 43673 22419 43707
rect 25421 43673 25455 43707
rect 10885 43605 10919 43639
rect 17969 43605 18003 43639
rect 21649 43605 21683 43639
rect 22017 43605 22051 43639
rect 24225 43605 24259 43639
rect 25329 43605 25363 43639
rect 7757 43401 7791 43435
rect 9505 43401 9539 43435
rect 10609 43401 10643 43435
rect 14105 43401 14139 43435
rect 15025 43401 15059 43435
rect 16773 43401 16807 43435
rect 17509 43401 17543 43435
rect 20085 43401 20119 43435
rect 22477 43401 22511 43435
rect 8677 43333 8711 43367
rect 12633 43333 12667 43367
rect 17417 43333 17451 43367
rect 23857 43333 23891 43367
rect 1685 43265 1719 43299
rect 2145 43265 2179 43299
rect 7941 43265 7975 43299
rect 8493 43265 8527 43299
rect 10517 43265 10551 43299
rect 12357 43265 12391 43299
rect 15117 43265 15151 43299
rect 22385 43265 22419 43299
rect 9597 43197 9631 43231
rect 9689 43197 9723 43231
rect 15209 43197 15243 43231
rect 17601 43197 17635 43231
rect 18337 43197 18371 43231
rect 18613 43197 18647 43231
rect 22661 43197 22695 43231
rect 23581 43197 23615 43231
rect 1869 43129 1903 43163
rect 9137 43129 9171 43163
rect 11069 43061 11103 43095
rect 14657 43061 14691 43095
rect 15669 43061 15703 43095
rect 17049 43061 17083 43095
rect 20453 43061 20487 43095
rect 21373 43061 21407 43095
rect 21649 43061 21683 43095
rect 22017 43061 22051 43095
rect 25329 43061 25363 43095
rect 8309 42857 8343 42891
rect 19796 42857 19830 42891
rect 17141 42789 17175 42823
rect 4997 42721 5031 42755
rect 10793 42721 10827 42755
rect 14841 42721 14875 42755
rect 17693 42721 17727 42755
rect 18153 42721 18187 42755
rect 19533 42721 19567 42755
rect 22293 42721 22327 42755
rect 22477 42721 22511 42755
rect 23213 42653 23247 42687
rect 23489 42653 23523 42687
rect 4813 42585 4847 42619
rect 9321 42585 9355 42619
rect 11069 42585 11103 42619
rect 15117 42585 15151 42619
rect 17509 42585 17543 42619
rect 25329 42585 25363 42619
rect 5273 42517 5307 42551
rect 8953 42517 8987 42551
rect 10333 42517 10367 42551
rect 12541 42517 12575 42551
rect 12817 42517 12851 42551
rect 14289 42517 14323 42551
rect 16589 42517 16623 42551
rect 17601 42517 17635 42551
rect 21281 42517 21315 42551
rect 21833 42517 21867 42551
rect 22201 42517 22235 42551
rect 24501 42517 24535 42551
rect 4353 42313 4387 42347
rect 5089 42313 5123 42347
rect 6745 42313 6779 42347
rect 11805 42313 11839 42347
rect 13001 42313 13035 42347
rect 15393 42313 15427 42347
rect 15853 42313 15887 42347
rect 16865 42313 16899 42347
rect 17233 42313 17267 42347
rect 20729 42313 20763 42347
rect 21281 42313 21315 42347
rect 25237 42313 25271 42347
rect 6653 42245 6687 42279
rect 12265 42245 12299 42279
rect 3893 42177 3927 42211
rect 4261 42177 4295 42211
rect 4997 42177 5031 42211
rect 7481 42177 7515 42211
rect 10057 42177 10091 42211
rect 12173 42177 12207 42211
rect 13369 42177 13403 42211
rect 14197 42177 14231 42211
rect 15761 42177 15795 42211
rect 18889 42177 18923 42211
rect 20637 42177 20671 42211
rect 22017 42177 22051 42211
rect 7757 42109 7791 42143
rect 10149 42109 10183 42143
rect 10241 42109 10275 42143
rect 12449 42109 12483 42143
rect 13461 42109 13495 42143
rect 13645 42109 13679 42143
rect 15945 42109 15979 42143
rect 17325 42109 17359 42143
rect 17417 42109 17451 42143
rect 19625 42109 19659 42143
rect 20821 42109 20855 42143
rect 22845 42109 22879 42143
rect 23489 42109 23523 42143
rect 23765 42109 23799 42143
rect 21557 42041 21591 42075
rect 5549 41973 5583 42007
rect 7205 41973 7239 42007
rect 9229 41973 9263 42007
rect 9689 41973 9723 42007
rect 10793 41973 10827 42007
rect 16405 41973 16439 42007
rect 18521 41973 18555 42007
rect 20269 41973 20303 42007
rect 5181 41769 5215 41803
rect 7665 41769 7699 41803
rect 8033 41769 8067 41803
rect 10701 41769 10735 41803
rect 17325 41769 17359 41803
rect 21189 41769 21223 41803
rect 21649 41701 21683 41735
rect 22845 41701 22879 41735
rect 5917 41633 5951 41667
rect 10149 41633 10183 41667
rect 11253 41633 11287 41667
rect 12725 41633 12759 41667
rect 16773 41633 16807 41667
rect 18613 41633 18647 41667
rect 18797 41633 18831 41667
rect 19441 41633 19475 41667
rect 22293 41633 22327 41667
rect 23305 41633 23339 41667
rect 23397 41633 23431 41667
rect 16681 41565 16715 41599
rect 24685 41565 24719 41599
rect 25329 41565 25363 41599
rect 5089 41497 5123 41531
rect 6193 41497 6227 41531
rect 9321 41497 9355 41531
rect 11989 41497 12023 41531
rect 13277 41497 13311 41531
rect 19717 41497 19751 41531
rect 22109 41497 22143 41531
rect 23213 41497 23247 41531
rect 24501 41497 24535 41531
rect 5641 41429 5675 41463
rect 11069 41429 11103 41463
rect 11161 41429 11195 41463
rect 16221 41429 16255 41463
rect 16589 41429 16623 41463
rect 18153 41429 18187 41463
rect 18521 41429 18555 41463
rect 22017 41429 22051 41463
rect 24869 41429 24903 41463
rect 25145 41429 25179 41463
rect 3341 41225 3375 41259
rect 11713 41225 11747 41259
rect 12173 41225 12207 41259
rect 19809 41225 19843 41259
rect 22017 41225 22051 41259
rect 24685 41225 24719 41259
rect 18889 41157 18923 41191
rect 19901 41157 19935 41191
rect 23213 41157 23247 41191
rect 1777 41089 1811 41123
rect 2053 41089 2087 41123
rect 3249 41089 3283 41123
rect 3709 41089 3743 41123
rect 8953 41089 8987 41123
rect 12081 41089 12115 41123
rect 13645 41089 13679 41123
rect 16865 41089 16899 41123
rect 21097 41089 21131 41123
rect 25329 41089 25363 41123
rect 9229 41021 9263 41055
rect 12265 41021 12299 41055
rect 13921 41021 13955 41055
rect 17141 41021 17175 41055
rect 19993 41021 20027 41055
rect 21189 41021 21223 41055
rect 21281 41021 21315 41055
rect 22937 41021 22971 41055
rect 1593 40885 1627 40919
rect 10701 40885 10735 40919
rect 11069 40885 11103 40919
rect 15393 40885 15427 40919
rect 15761 40885 15795 40919
rect 18613 40885 18647 40919
rect 19073 40885 19107 40919
rect 19441 40885 19475 40919
rect 20729 40885 20763 40919
rect 25145 40885 25179 40919
rect 8309 40681 8343 40715
rect 20913 40681 20947 40715
rect 9229 40613 9263 40647
rect 10701 40613 10735 40647
rect 12633 40613 12667 40647
rect 13737 40613 13771 40647
rect 22109 40613 22143 40647
rect 22477 40613 22511 40647
rect 6469 40545 6503 40579
rect 9781 40545 9815 40579
rect 11897 40545 11931 40579
rect 11989 40545 12023 40579
rect 13277 40545 13311 40579
rect 15761 40545 15795 40579
rect 17141 40545 17175 40579
rect 17233 40545 17267 40579
rect 21373 40545 21407 40579
rect 21557 40545 21591 40579
rect 23029 40545 23063 40579
rect 6193 40477 6227 40511
rect 13001 40477 13035 40511
rect 13093 40477 13127 40511
rect 15577 40477 15611 40511
rect 22845 40477 22879 40511
rect 22937 40477 22971 40511
rect 24409 40477 24443 40511
rect 24685 40477 24719 40511
rect 25329 40477 25363 40511
rect 9597 40409 9631 40443
rect 11345 40409 11379 40443
rect 11805 40409 11839 40443
rect 15669 40409 15703 40443
rect 20361 40409 20395 40443
rect 22017 40409 22051 40443
rect 24869 40409 24903 40443
rect 7941 40341 7975 40375
rect 9689 40341 9723 40375
rect 11437 40341 11471 40375
rect 15209 40341 15243 40375
rect 16681 40341 16715 40375
rect 17049 40341 17083 40375
rect 21281 40341 21315 40375
rect 24041 40341 24075 40375
rect 24225 40341 24259 40375
rect 25145 40341 25179 40375
rect 7297 40137 7331 40171
rect 15025 40137 15059 40171
rect 15577 40137 15611 40171
rect 19809 40137 19843 40171
rect 25237 40137 25271 40171
rect 7665 40069 7699 40103
rect 10517 40069 10551 40103
rect 15945 40069 15979 40103
rect 18613 40069 18647 40103
rect 20177 40069 20211 40103
rect 22293 40069 22327 40103
rect 8493 40001 8527 40035
rect 12909 40001 12943 40035
rect 21097 40001 21131 40035
rect 23489 40001 23523 40035
rect 7757 39933 7791 39967
rect 7849 39933 7883 39967
rect 8769 39933 8803 39967
rect 10977 39933 11011 39967
rect 13185 39933 13219 39967
rect 16037 39933 16071 39967
rect 16129 39933 16163 39967
rect 18705 39933 18739 39967
rect 18797 39933 18831 39967
rect 20269 39933 20303 39967
rect 20361 39933 20395 39967
rect 23765 39933 23799 39967
rect 20821 39865 20855 39899
rect 14657 39797 14691 39831
rect 18245 39797 18279 39831
rect 6653 39593 6687 39627
rect 9781 39593 9815 39627
rect 13093 39593 13127 39627
rect 14381 39593 14415 39627
rect 21281 39593 21315 39627
rect 15577 39525 15611 39559
rect 22661 39525 22695 39559
rect 4905 39457 4939 39491
rect 10241 39457 10275 39491
rect 10333 39457 10367 39491
rect 10977 39457 11011 39491
rect 15025 39457 15059 39491
rect 16221 39457 16255 39491
rect 19901 39457 19935 39491
rect 20085 39457 20119 39491
rect 21833 39457 21867 39491
rect 23305 39457 23339 39491
rect 25053 39457 25087 39491
rect 25237 39457 25271 39491
rect 23121 39389 23155 39423
rect 24961 39389 24995 39423
rect 5181 39321 5215 39355
rect 11253 39321 11287 39355
rect 14841 39321 14875 39355
rect 19809 39321 19843 39355
rect 20453 39321 20487 39355
rect 21741 39321 21775 39355
rect 22293 39321 22327 39355
rect 23029 39321 23063 39355
rect 23857 39321 23891 39355
rect 7021 39253 7055 39287
rect 9137 39253 9171 39287
rect 10149 39253 10183 39287
rect 12725 39253 12759 39287
rect 13829 39253 13863 39287
rect 14749 39253 14783 39287
rect 15945 39253 15979 39287
rect 16037 39253 16071 39287
rect 18797 39253 18831 39287
rect 19441 39253 19475 39287
rect 21649 39253 21683 39287
rect 24593 39253 24627 39287
rect 7389 39049 7423 39083
rect 8769 39049 8803 39083
rect 9505 39049 9539 39083
rect 10793 39049 10827 39083
rect 14289 39049 14323 39083
rect 15301 39049 15335 39083
rect 19165 39049 19199 39083
rect 20729 39049 20763 39083
rect 24501 39049 24535 39083
rect 10885 38981 10919 39015
rect 11529 38981 11563 39015
rect 19625 38981 19659 39015
rect 24133 38981 24167 39015
rect 12081 38913 12115 38947
rect 18337 38913 18371 38947
rect 19533 38913 19567 38947
rect 24685 38913 24719 38947
rect 25329 38913 25363 38947
rect 8585 38845 8619 38879
rect 9597 38845 9631 38879
rect 9689 38845 9723 38879
rect 10977 38845 11011 38879
rect 12357 38845 12391 38879
rect 15393 38845 15427 38879
rect 15577 38845 15611 38879
rect 16865 38845 16899 38879
rect 18429 38845 18463 38879
rect 18613 38845 18647 38879
rect 19717 38845 19751 38879
rect 20821 38845 20855 38879
rect 20913 38845 20947 38879
rect 22109 38845 22143 38879
rect 22385 38845 22419 38879
rect 10425 38777 10459 38811
rect 14933 38777 14967 38811
rect 9137 38709 9171 38743
rect 13829 38709 13863 38743
rect 16037 38709 16071 38743
rect 17969 38709 18003 38743
rect 20361 38709 20395 38743
rect 23857 38709 23891 38743
rect 25145 38709 25179 38743
rect 7849 38505 7883 38539
rect 10425 38505 10459 38539
rect 14289 38505 14323 38539
rect 18153 38505 18187 38539
rect 19441 38505 19475 38539
rect 11897 38437 11931 38471
rect 5457 38369 5491 38403
rect 7205 38369 7239 38403
rect 8493 38369 8527 38403
rect 9689 38369 9723 38403
rect 9781 38369 9815 38403
rect 10977 38369 11011 38403
rect 12357 38369 12391 38403
rect 12449 38369 12483 38403
rect 14841 38369 14875 38403
rect 16221 38369 16255 38403
rect 18705 38369 18739 38403
rect 19993 38369 20027 38403
rect 21097 38369 21131 38403
rect 21189 38369 21223 38403
rect 22477 38369 22511 38403
rect 22569 38369 22603 38403
rect 23765 38369 23799 38403
rect 25145 38369 25179 38403
rect 1777 38301 1811 38335
rect 2053 38301 2087 38335
rect 8217 38301 8251 38335
rect 13921 38301 13955 38335
rect 14749 38301 14783 38335
rect 15945 38301 15979 38335
rect 25053 38301 25087 38335
rect 5733 38233 5767 38267
rect 9597 38233 9631 38267
rect 18613 38233 18647 38267
rect 19901 38233 19935 38267
rect 22385 38233 22419 38267
rect 1593 38165 1627 38199
rect 7573 38165 7607 38199
rect 8309 38165 8343 38199
rect 9229 38165 9263 38199
rect 10793 38165 10827 38199
rect 10885 38165 10919 38199
rect 12265 38165 12299 38199
rect 14657 38165 14691 38199
rect 17693 38165 17727 38199
rect 18521 38165 18555 38199
rect 19809 38165 19843 38199
rect 20637 38165 20671 38199
rect 21005 38165 21039 38199
rect 22017 38165 22051 38199
rect 23213 38165 23247 38199
rect 23581 38165 23615 38199
rect 23673 38165 23707 38199
rect 24593 38165 24627 38199
rect 24961 38165 24995 38199
rect 5273 37961 5307 37995
rect 5733 37961 5767 37995
rect 9045 37961 9079 37995
rect 11713 37961 11747 37995
rect 12817 37961 12851 37995
rect 14105 37961 14139 37995
rect 16405 37961 16439 37995
rect 17233 37961 17267 37995
rect 17969 37961 18003 37995
rect 18981 37961 19015 37995
rect 19441 37961 19475 37995
rect 20269 37961 20303 37995
rect 22017 37961 22051 37995
rect 6837 37893 6871 37927
rect 17325 37893 17359 37927
rect 21373 37893 21407 37927
rect 23857 37893 23891 37927
rect 5641 37825 5675 37859
rect 9413 37825 9447 37859
rect 10425 37825 10459 37859
rect 12725 37825 12759 37859
rect 14381 37825 14415 37859
rect 15393 37825 15427 37859
rect 15485 37825 15519 37859
rect 18705 37825 18739 37859
rect 19349 37825 19383 37859
rect 20637 37825 20671 37859
rect 21557 37825 21591 37859
rect 22385 37825 22419 37859
rect 22477 37825 22511 37859
rect 23121 37825 23155 37859
rect 5825 37757 5859 37791
rect 6561 37757 6595 37791
rect 8585 37757 8619 37791
rect 10517 37757 10551 37791
rect 10609 37757 10643 37791
rect 13001 37757 13035 37791
rect 13553 37757 13587 37791
rect 15669 37757 15703 37791
rect 17509 37757 17543 37791
rect 19625 37757 19659 37791
rect 20729 37757 20763 37791
rect 20913 37757 20947 37791
rect 22569 37757 22603 37791
rect 23213 37757 23247 37791
rect 23581 37757 23615 37791
rect 25329 37757 25363 37791
rect 10057 37689 10091 37723
rect 16865 37689 16899 37723
rect 8861 37621 8895 37655
rect 12357 37621 12391 37655
rect 15025 37621 15059 37655
rect 8585 37417 8619 37451
rect 10425 37417 10459 37451
rect 14381 37417 14415 37451
rect 17325 37417 17359 37451
rect 23949 37417 23983 37451
rect 14657 37349 14691 37383
rect 18981 37349 19015 37383
rect 23857 37349 23891 37383
rect 24685 37349 24719 37383
rect 7113 37281 7147 37315
rect 11805 37281 11839 37315
rect 12449 37281 12483 37315
rect 13369 37281 13403 37315
rect 13461 37281 13495 37315
rect 15485 37281 15519 37315
rect 16589 37281 16623 37315
rect 16681 37281 16715 37315
rect 17877 37281 17911 37315
rect 20637 37281 20671 37315
rect 24593 37281 24627 37315
rect 6837 37213 6871 37247
rect 9137 37213 9171 37247
rect 11713 37213 11747 37247
rect 13277 37213 13311 37247
rect 16497 37213 16531 37247
rect 17785 37213 17819 37247
rect 19441 37213 19475 37247
rect 21097 37213 21131 37247
rect 21465 37213 21499 37247
rect 22201 37213 22235 37247
rect 25329 37213 25363 37247
rect 9873 37145 9907 37179
rect 11621 37145 11655 37179
rect 14197 37145 14231 37179
rect 17693 37145 17727 37179
rect 20177 37145 20211 37179
rect 24225 37145 24259 37179
rect 11253 37077 11287 37111
rect 12633 37077 12667 37111
rect 12909 37077 12943 37111
rect 14933 37077 14967 37111
rect 15301 37077 15335 37111
rect 15393 37077 15427 37111
rect 16129 37077 16163 37111
rect 18521 37077 18555 37111
rect 25145 37077 25179 37111
rect 7481 36873 7515 36907
rect 7941 36873 7975 36907
rect 9045 36873 9079 36907
rect 11621 36873 11655 36907
rect 17049 36873 17083 36907
rect 17417 36873 17451 36907
rect 20453 36873 20487 36907
rect 24593 36873 24627 36907
rect 6101 36805 6135 36839
rect 8677 36805 8711 36839
rect 10241 36805 10275 36839
rect 12633 36805 12667 36839
rect 13829 36805 13863 36839
rect 15577 36805 15611 36839
rect 20361 36805 20395 36839
rect 23121 36805 23155 36839
rect 3985 36737 4019 36771
rect 7849 36737 7883 36771
rect 9413 36737 9447 36771
rect 9505 36737 9539 36771
rect 12081 36737 12115 36771
rect 12541 36737 12575 36771
rect 13737 36737 13771 36771
rect 14933 36737 14967 36771
rect 16773 36737 16807 36771
rect 17509 36737 17543 36771
rect 22845 36737 22879 36771
rect 25329 36737 25363 36771
rect 4261 36669 4295 36703
rect 5733 36669 5767 36703
rect 8033 36669 8067 36703
rect 9597 36669 9631 36703
rect 10977 36669 11011 36703
rect 12817 36669 12851 36703
rect 13921 36669 13955 36703
rect 15025 36669 15059 36703
rect 15117 36669 15151 36703
rect 17693 36669 17727 36703
rect 20545 36669 20579 36703
rect 12173 36533 12207 36567
rect 13369 36533 13403 36567
rect 14565 36533 14599 36567
rect 15853 36533 15887 36567
rect 19993 36533 20027 36567
rect 25145 36533 25179 36567
rect 7665 36329 7699 36363
rect 9137 36329 9171 36363
rect 12173 36329 12207 36363
rect 12725 36329 12759 36363
rect 14289 36329 14323 36363
rect 16129 36261 16163 36295
rect 19441 36261 19475 36295
rect 25145 36261 25179 36295
rect 8217 36193 8251 36227
rect 9689 36193 9723 36227
rect 13277 36193 13311 36227
rect 13829 36193 13863 36227
rect 14749 36193 14783 36227
rect 14841 36193 14875 36227
rect 16773 36193 16807 36227
rect 19993 36193 20027 36227
rect 21281 36193 21315 36227
rect 21373 36193 21407 36227
rect 23765 36193 23799 36227
rect 23949 36193 23983 36227
rect 1777 36125 1811 36159
rect 2053 36125 2087 36159
rect 9597 36125 9631 36159
rect 13185 36125 13219 36159
rect 16589 36125 16623 36159
rect 24869 36125 24903 36159
rect 25329 36125 25363 36159
rect 9505 36057 9539 36091
rect 16497 36057 16531 36091
rect 17325 36057 17359 36091
rect 19901 36057 19935 36091
rect 1593 35989 1627 36023
rect 8033 35989 8067 36023
rect 8125 35989 8159 36023
rect 12449 35989 12483 36023
rect 13093 35989 13127 36023
rect 14657 35989 14691 36023
rect 15761 35989 15795 36023
rect 19809 35989 19843 36023
rect 20821 35989 20855 36023
rect 21189 35989 21223 36023
rect 23305 35989 23339 36023
rect 23673 35989 23707 36023
rect 24041 35989 24075 36023
rect 25145 35989 25179 36023
rect 6009 35785 6043 35819
rect 6469 35785 6503 35819
rect 13829 35785 13863 35819
rect 14473 35785 14507 35819
rect 20177 35785 20211 35819
rect 17877 35717 17911 35751
rect 20269 35717 20303 35751
rect 4261 35649 4295 35683
rect 23121 35649 23155 35683
rect 4537 35581 4571 35615
rect 8125 35581 8159 35615
rect 8401 35581 8435 35615
rect 11713 35581 11747 35615
rect 11989 35581 12023 35615
rect 17601 35581 17635 35615
rect 20361 35581 20395 35615
rect 22477 35581 22511 35615
rect 23397 35581 23431 35615
rect 25237 35581 25271 35615
rect 13461 35513 13495 35547
rect 19349 35513 19383 35547
rect 9873 35445 9907 35479
rect 10241 35445 10275 35479
rect 19809 35445 19843 35479
rect 20913 35445 20947 35479
rect 24869 35445 24903 35479
rect 25421 35445 25455 35479
rect 7849 35241 7883 35275
rect 8217 35241 8251 35275
rect 9321 35241 9355 35275
rect 13001 35241 13035 35275
rect 17141 35241 17175 35275
rect 17509 35241 17543 35275
rect 19704 35241 19738 35275
rect 6101 35105 6135 35139
rect 6377 35105 6411 35139
rect 9873 35105 9907 35139
rect 13553 35105 13587 35139
rect 15393 35105 15427 35139
rect 19441 35105 19475 35139
rect 24409 35105 24443 35139
rect 13461 35037 13495 35071
rect 22293 35037 22327 35071
rect 25329 35037 25363 35071
rect 9689 34969 9723 35003
rect 15669 34969 15703 35003
rect 22569 34969 22603 35003
rect 9781 34901 9815 34935
rect 13369 34901 13403 34935
rect 21189 34901 21223 34935
rect 21557 34901 21591 34935
rect 24041 34901 24075 34935
rect 25145 34901 25179 34935
rect 10609 34697 10643 34731
rect 13829 34697 13863 34731
rect 15577 34697 15611 34731
rect 15945 34697 15979 34731
rect 21097 34697 21131 34731
rect 21189 34697 21223 34731
rect 22385 34697 22419 34731
rect 22477 34697 22511 34731
rect 23581 34697 23615 34731
rect 24409 34697 24443 34731
rect 25145 34697 25179 34731
rect 6837 34629 6871 34663
rect 16037 34629 16071 34663
rect 6561 34561 6595 34595
rect 8868 34561 8902 34595
rect 24593 34561 24627 34595
rect 25329 34561 25363 34595
rect 8309 34493 8343 34527
rect 11713 34493 11747 34527
rect 13461 34493 13495 34527
rect 16129 34493 16163 34527
rect 21281 34493 21315 34527
rect 22569 34493 22603 34527
rect 23673 34493 23707 34527
rect 23765 34493 23799 34527
rect 10885 34425 10919 34459
rect 23213 34425 23247 34459
rect 9124 34357 9158 34391
rect 11976 34357 12010 34391
rect 20729 34357 20763 34391
rect 22017 34357 22051 34391
rect 7573 34153 7607 34187
rect 8493 34153 8527 34187
rect 9137 34153 9171 34187
rect 12173 34153 12207 34187
rect 17693 34153 17727 34187
rect 20453 34153 20487 34187
rect 25329 34153 25363 34187
rect 25421 34153 25455 34187
rect 21097 34085 21131 34119
rect 5549 34017 5583 34051
rect 7297 34017 7331 34051
rect 9689 34017 9723 34051
rect 10701 34017 10735 34051
rect 13461 34017 13495 34051
rect 13553 34017 13587 34051
rect 15945 34017 15979 34051
rect 19993 34017 20027 34051
rect 21649 34017 21683 34051
rect 22753 34017 22787 34051
rect 22937 34017 22971 34051
rect 10425 33949 10459 33983
rect 14105 33949 14139 33983
rect 17969 33949 18003 33983
rect 19901 33949 19935 33983
rect 21557 33949 21591 33983
rect 24777 33949 24811 33983
rect 5825 33881 5859 33915
rect 9505 33881 9539 33915
rect 16221 33881 16255 33915
rect 19809 33881 19843 33915
rect 22661 33881 22695 33915
rect 9597 33813 9631 33847
rect 12449 33813 12483 33847
rect 13001 33813 13035 33847
rect 13369 33813 13403 33847
rect 19441 33813 19475 33847
rect 20637 33813 20671 33847
rect 21465 33813 21499 33847
rect 22293 33813 22327 33847
rect 24593 33813 24627 33847
rect 7205 33609 7239 33643
rect 10425 33609 10459 33643
rect 10885 33609 10919 33643
rect 12909 33609 12943 33643
rect 13369 33609 13403 33643
rect 16221 33609 16255 33643
rect 19809 33609 19843 33643
rect 20269 33609 20303 33643
rect 20637 33609 20671 33643
rect 22661 33609 22695 33643
rect 1777 33473 1811 33507
rect 2053 33473 2087 33507
rect 10793 33473 10827 33507
rect 13277 33473 13311 33507
rect 14105 33473 14139 33507
rect 18061 33473 18095 33507
rect 20729 33473 20763 33507
rect 23489 33473 23523 33507
rect 5365 33405 5399 33439
rect 9781 33405 9815 33439
rect 10977 33405 11011 33439
rect 12541 33405 12575 33439
rect 13553 33405 13587 33439
rect 14381 33405 14415 33439
rect 18337 33405 18371 33439
rect 20913 33405 20947 33439
rect 22017 33405 22051 33439
rect 23765 33405 23799 33439
rect 1593 33269 1627 33303
rect 15853 33269 15887 33303
rect 21281 33269 21315 33303
rect 25237 33269 25271 33303
rect 7481 33065 7515 33099
rect 9413 33065 9447 33099
rect 10609 33065 10643 33099
rect 11161 33065 11195 33099
rect 17417 33065 17451 33099
rect 19809 33065 19843 33099
rect 22201 33065 22235 33099
rect 15761 32997 15795 33031
rect 17233 32997 17267 33031
rect 5273 32929 5307 32963
rect 7021 32929 7055 32963
rect 8125 32929 8159 32963
rect 9965 32929 9999 32963
rect 11713 32929 11747 32963
rect 14749 32929 14783 32963
rect 14841 32929 14875 32963
rect 16589 32929 16623 32963
rect 16773 32929 16807 32963
rect 20453 32929 20487 32963
rect 21465 32929 21499 32963
rect 21557 32929 21591 32963
rect 9781 32861 9815 32895
rect 16497 32861 16531 32895
rect 20177 32861 20211 32895
rect 22385 32861 22419 32895
rect 22753 32861 22787 32895
rect 24869 32861 24903 32895
rect 25329 32861 25363 32895
rect 5549 32793 5583 32827
rect 7941 32793 7975 32827
rect 10885 32793 10919 32827
rect 11621 32793 11655 32827
rect 19441 32793 19475 32827
rect 20269 32793 20303 32827
rect 7849 32725 7883 32759
rect 9873 32725 9907 32759
rect 11529 32725 11563 32759
rect 14289 32725 14323 32759
rect 14657 32725 14691 32759
rect 16129 32725 16163 32759
rect 21005 32725 21039 32759
rect 21373 32725 21407 32759
rect 22845 32725 22879 32759
rect 25145 32725 25179 32759
rect 4629 32521 4663 32555
rect 4997 32521 5031 32555
rect 5365 32521 5399 32555
rect 6929 32521 6963 32555
rect 9321 32521 9355 32555
rect 11989 32521 12023 32555
rect 17325 32521 17359 32555
rect 21189 32521 21223 32555
rect 21925 32521 21959 32555
rect 22201 32521 22235 32555
rect 22845 32521 22879 32555
rect 24869 32521 24903 32555
rect 5457 32453 5491 32487
rect 18429 32453 18463 32487
rect 18521 32453 18555 32487
rect 7573 32385 7607 32419
rect 12357 32385 12391 32419
rect 13185 32385 13219 32419
rect 14565 32385 14599 32419
rect 17233 32385 17267 32419
rect 20269 32385 20303 32419
rect 21097 32385 21131 32419
rect 22385 32385 22419 32419
rect 23029 32385 23063 32419
rect 25329 32385 25363 32419
rect 5549 32317 5583 32351
rect 7849 32317 7883 32351
rect 9873 32317 9907 32351
rect 11713 32317 11747 32351
rect 12449 32317 12483 32351
rect 12541 32317 12575 32351
rect 14841 32317 14875 32351
rect 17509 32317 17543 32351
rect 18705 32317 18739 32351
rect 21373 32317 21407 32351
rect 23305 32317 23339 32351
rect 16313 32249 16347 32283
rect 25145 32249 25179 32283
rect 10425 32181 10459 32215
rect 16865 32181 16899 32215
rect 18061 32181 18095 32215
rect 20085 32181 20119 32215
rect 20729 32181 20763 32215
rect 7941 31977 7975 32011
rect 9676 31977 9710 32011
rect 11161 31977 11195 32011
rect 16405 31977 16439 32011
rect 24133 31977 24167 32011
rect 25145 31977 25179 32011
rect 14289 31909 14323 31943
rect 21925 31909 21959 31943
rect 6193 31841 6227 31875
rect 6469 31841 6503 31875
rect 8309 31841 8343 31875
rect 14933 31841 14967 31875
rect 16957 31841 16991 31875
rect 19993 31841 20027 31875
rect 21189 31841 21223 31875
rect 22385 31841 22419 31875
rect 22569 31841 22603 31875
rect 9413 31773 9447 31807
rect 11529 31773 11563 31807
rect 14749 31773 14783 31807
rect 16865 31773 16899 31807
rect 18061 31773 18095 31807
rect 19901 31773 19935 31807
rect 21097 31773 21131 31807
rect 24869 31773 24903 31807
rect 25329 31773 25363 31807
rect 19809 31705 19843 31739
rect 21005 31705 21039 31739
rect 13921 31637 13955 31671
rect 14657 31637 14691 31671
rect 16773 31637 16807 31671
rect 19441 31637 19475 31671
rect 20637 31637 20671 31671
rect 22293 31637 22327 31671
rect 7481 31433 7515 31467
rect 8677 31433 8711 31467
rect 9045 31433 9079 31467
rect 15025 31433 15059 31467
rect 17601 31433 17635 31467
rect 18337 31433 18371 31467
rect 19533 31433 19567 31467
rect 21557 31433 21591 31467
rect 25145 31433 25179 31467
rect 19901 31365 19935 31399
rect 22477 31365 22511 31399
rect 1777 31297 1811 31331
rect 7849 31297 7883 31331
rect 7941 31297 7975 31331
rect 17509 31297 17543 31331
rect 18705 31297 18739 31331
rect 20729 31297 20763 31331
rect 24593 31297 24627 31331
rect 25329 31297 25363 31331
rect 2053 31229 2087 31263
rect 7205 31229 7239 31263
rect 8125 31229 8159 31263
rect 9137 31229 9171 31263
rect 9229 31229 9263 31263
rect 12909 31229 12943 31263
rect 13185 31229 13219 31263
rect 16773 31229 16807 31263
rect 17785 31229 17819 31263
rect 18797 31229 18831 31263
rect 18889 31229 18923 31263
rect 19993 31229 20027 31263
rect 20177 31229 20211 31263
rect 22201 31229 22235 31263
rect 14657 31093 14691 31127
rect 17141 31093 17175 31127
rect 20545 31093 20579 31127
rect 23949 31093 23983 31127
rect 24409 31093 24443 31127
rect 12817 30889 12851 30923
rect 15945 30889 15979 30923
rect 18245 30889 18279 30923
rect 20453 30889 20487 30923
rect 23121 30889 23155 30923
rect 24869 30889 24903 30923
rect 11621 30821 11655 30855
rect 3985 30753 4019 30787
rect 7941 30753 7975 30787
rect 9597 30753 9631 30787
rect 9873 30753 9907 30787
rect 13369 30753 13403 30787
rect 16221 30753 16255 30787
rect 16497 30753 16531 30787
rect 19901 30753 19935 30787
rect 19993 30753 20027 30787
rect 22569 30753 22603 30787
rect 12541 30685 12575 30719
rect 13185 30685 13219 30719
rect 19809 30685 19843 30719
rect 22385 30685 22419 30719
rect 23857 30685 23891 30719
rect 25329 30685 25363 30719
rect 4169 30617 4203 30651
rect 5825 30617 5859 30651
rect 13277 30617 13311 30651
rect 8493 30549 8527 30583
rect 11345 30549 11379 30583
rect 17969 30549 18003 30583
rect 19441 30549 19475 30583
rect 22017 30549 22051 30583
rect 22477 30549 22511 30583
rect 23673 30549 23707 30583
rect 25145 30549 25179 30583
rect 12541 30345 12575 30379
rect 23673 30277 23707 30311
rect 10793 30209 10827 30243
rect 11713 30209 11747 30243
rect 14473 30209 14507 30243
rect 17969 30209 18003 30243
rect 18613 30209 18647 30243
rect 18889 30209 18923 30243
rect 19625 30209 19659 30243
rect 23397 30209 23431 30243
rect 10149 30141 10183 30175
rect 10885 30141 10919 30175
rect 10977 30141 11011 30175
rect 14749 30141 14783 30175
rect 16221 30141 16255 30175
rect 16957 30141 16991 30175
rect 18061 30141 18095 30175
rect 18245 30141 18279 30175
rect 25145 30141 25179 30175
rect 10425 30005 10459 30039
rect 12265 30005 12299 30039
rect 17601 30005 17635 30039
rect 19441 30005 19475 30039
rect 25421 30005 25455 30039
rect 7297 29801 7331 29835
rect 7849 29801 7883 29835
rect 9505 29801 9539 29835
rect 16037 29801 16071 29835
rect 8953 29733 8987 29767
rect 12633 29733 12667 29767
rect 25145 29733 25179 29767
rect 4261 29665 4295 29699
rect 8401 29665 8435 29699
rect 10057 29665 10091 29699
rect 11989 29665 12023 29699
rect 13185 29665 13219 29699
rect 17509 29665 17543 29699
rect 18797 29665 18831 29699
rect 20085 29665 20119 29699
rect 20269 29665 20303 29699
rect 22201 29665 22235 29699
rect 23397 29665 23431 29699
rect 23581 29665 23615 29699
rect 11805 29597 11839 29631
rect 13093 29597 13127 29631
rect 13737 29597 13771 29631
rect 19993 29597 20027 29631
rect 21925 29597 21959 29631
rect 25329 29597 25363 29631
rect 4445 29529 4479 29563
rect 6101 29529 6135 29563
rect 8309 29529 8343 29563
rect 9873 29529 9907 29563
rect 9965 29529 9999 29563
rect 13001 29529 13035 29563
rect 14749 29529 14783 29563
rect 17325 29529 17359 29563
rect 18613 29529 18647 29563
rect 7481 29461 7515 29495
rect 8217 29461 8251 29495
rect 9229 29461 9263 29495
rect 11437 29461 11471 29495
rect 11897 29461 11931 29495
rect 16957 29461 16991 29495
rect 17417 29461 17451 29495
rect 18153 29461 18187 29495
rect 18521 29461 18555 29495
rect 19625 29461 19659 29495
rect 20913 29461 20947 29495
rect 21557 29461 21591 29495
rect 22017 29461 22051 29495
rect 22937 29461 22971 29495
rect 23305 29461 23339 29495
rect 9781 29257 9815 29291
rect 14933 29257 14967 29291
rect 15301 29257 15335 29291
rect 15945 29257 15979 29291
rect 17233 29257 17267 29291
rect 17325 29257 17359 29291
rect 17969 29257 18003 29291
rect 20085 29257 20119 29291
rect 20545 29257 20579 29291
rect 22385 29257 22419 29291
rect 23949 29257 23983 29291
rect 25329 29257 25363 29291
rect 25513 29257 25547 29291
rect 16221 29189 16255 29223
rect 24685 29189 24719 29223
rect 12909 29121 12943 29155
rect 14105 29121 14139 29155
rect 14197 29121 14231 29155
rect 16497 29121 16531 29155
rect 19717 29121 19751 29155
rect 20453 29121 20487 29155
rect 21557 29121 21591 29155
rect 23673 29121 23707 29155
rect 24133 29121 24167 29155
rect 7757 29053 7791 29087
rect 9505 29053 9539 29087
rect 13001 29053 13035 29087
rect 13185 29053 13219 29087
rect 14381 29053 14415 29087
rect 15393 29053 15427 29087
rect 15485 29053 15519 29087
rect 17417 29053 17451 29087
rect 20637 29053 20671 29087
rect 22477 29053 22511 29087
rect 22661 29053 22695 29087
rect 12541 28985 12575 29019
rect 13737 28985 13771 29019
rect 16865 28985 16899 29019
rect 18061 28985 18095 29019
rect 21097 28985 21131 29019
rect 22017 28985 22051 29019
rect 24869 28985 24903 29019
rect 8020 28917 8054 28951
rect 12817 28713 12851 28747
rect 16773 28713 16807 28747
rect 21189 28645 21223 28679
rect 2053 28577 2087 28611
rect 4261 28577 4295 28611
rect 5917 28577 5951 28611
rect 6561 28577 6595 28611
rect 6837 28577 6871 28611
rect 8309 28577 8343 28611
rect 10885 28577 10919 28611
rect 13369 28577 13403 28611
rect 14841 28577 14875 28611
rect 16221 28577 16255 28611
rect 17693 28577 17727 28611
rect 17785 28577 17819 28611
rect 19441 28577 19475 28611
rect 1777 28509 1811 28543
rect 10609 28509 10643 28543
rect 14657 28509 14691 28543
rect 16037 28509 16071 28543
rect 16129 28509 16163 28543
rect 17601 28509 17635 28543
rect 24041 28509 24075 28543
rect 24777 28509 24811 28543
rect 4445 28441 4479 28475
rect 13277 28441 13311 28475
rect 19717 28441 19751 28475
rect 21465 28441 21499 28475
rect 8677 28373 8711 28407
rect 12357 28373 12391 28407
rect 13185 28373 13219 28407
rect 13921 28373 13955 28407
rect 14289 28373 14323 28407
rect 14749 28373 14783 28407
rect 15301 28373 15335 28407
rect 15669 28373 15703 28407
rect 17233 28373 17267 28407
rect 23857 28373 23891 28407
rect 24593 28373 24627 28407
rect 2053 28169 2087 28203
rect 3755 28169 3789 28203
rect 12633 28169 12667 28203
rect 15945 28169 15979 28203
rect 16681 28169 16715 28203
rect 18337 28169 18371 28203
rect 19533 28169 19567 28203
rect 20177 28169 20211 28203
rect 23765 28169 23799 28203
rect 24225 28169 24259 28203
rect 24685 28101 24719 28135
rect 2237 28033 2271 28067
rect 3652 28033 3686 28067
rect 10333 28033 10367 28067
rect 18245 28033 18279 28067
rect 19441 28033 19475 28067
rect 22017 28033 22051 28067
rect 8309 27965 8343 27999
rect 8585 27965 8619 27999
rect 16037 27965 16071 27999
rect 16221 27965 16255 27999
rect 18521 27965 18555 27999
rect 19717 27965 19751 27999
rect 22293 27965 22327 27999
rect 10057 27897 10091 27931
rect 17509 27897 17543 27931
rect 24869 27897 24903 27931
rect 13093 27829 13127 27863
rect 13369 27829 13403 27863
rect 15117 27829 15151 27863
rect 15577 27829 15611 27863
rect 16957 27829 16991 27863
rect 17877 27829 17911 27863
rect 19073 27829 19107 27863
rect 6456 27625 6490 27659
rect 18705 27625 18739 27659
rect 24225 27625 24259 27659
rect 7941 27557 7975 27591
rect 16405 27557 16439 27591
rect 20085 27557 20119 27591
rect 25145 27557 25179 27591
rect 6193 27489 6227 27523
rect 8309 27489 8343 27523
rect 8401 27489 8435 27523
rect 15669 27489 15703 27523
rect 20637 27489 20671 27523
rect 21925 27489 21959 27523
rect 11161 27421 11195 27455
rect 18337 27421 18371 27455
rect 24685 27421 24719 27455
rect 11437 27353 11471 27387
rect 13277 27353 13311 27387
rect 15577 27353 15611 27387
rect 16129 27353 16163 27387
rect 18889 27353 18923 27387
rect 20545 27353 20579 27387
rect 22201 27353 22235 27387
rect 24869 27353 24903 27387
rect 12909 27285 12943 27319
rect 15117 27285 15151 27319
rect 15485 27285 15519 27319
rect 18153 27285 18187 27319
rect 19809 27285 19843 27319
rect 20453 27285 20487 27319
rect 23673 27285 23707 27319
rect 3203 27081 3237 27115
rect 15209 27081 15243 27115
rect 17601 27081 17635 27115
rect 19993 27081 20027 27115
rect 10517 27013 10551 27047
rect 18061 27013 18095 27047
rect 23121 27013 23155 27047
rect 25145 27013 25179 27047
rect 3132 26945 3166 26979
rect 3709 26945 3743 26979
rect 6561 26945 6595 26979
rect 9137 26945 9171 26979
rect 12541 26945 12575 26979
rect 15117 26945 15151 26979
rect 17969 26945 18003 26979
rect 19901 26945 19935 26979
rect 20729 26945 20763 26979
rect 22385 26945 22419 26979
rect 3893 26877 3927 26911
rect 4445 26877 4479 26911
rect 6837 26877 6871 26911
rect 9229 26877 9263 26911
rect 9413 26877 9447 26911
rect 12817 26877 12851 26911
rect 15301 26877 15335 26911
rect 18245 26877 18279 26911
rect 20177 26877 20211 26911
rect 22845 26877 22879 26911
rect 25329 26877 25363 26911
rect 8309 26809 8343 26843
rect 10701 26809 10735 26843
rect 14749 26809 14783 26843
rect 8769 26741 8803 26775
rect 11805 26741 11839 26775
rect 14289 26741 14323 26775
rect 17233 26741 17267 26775
rect 19533 26741 19567 26775
rect 22201 26741 22235 26775
rect 24593 26741 24627 26775
rect 4077 26537 4111 26571
rect 11713 26537 11747 26571
rect 17141 26537 17175 26571
rect 22385 26537 22419 26571
rect 19441 26469 19475 26503
rect 22845 26469 22879 26503
rect 23857 26469 23891 26503
rect 25145 26469 25179 26503
rect 6469 26401 6503 26435
rect 6745 26401 6779 26435
rect 9137 26401 9171 26435
rect 10241 26401 10275 26435
rect 12725 26401 12759 26435
rect 15669 26401 15703 26435
rect 19901 26401 19935 26435
rect 20085 26401 20119 26435
rect 20637 26401 20671 26435
rect 23305 26401 23339 26435
rect 23489 26401 23523 26435
rect 1777 26333 1811 26367
rect 9965 26333 9999 26367
rect 12633 26333 12667 26367
rect 15393 26333 15427 26367
rect 23213 26333 23247 26367
rect 24685 26333 24719 26367
rect 2789 26265 2823 26299
rect 8677 26265 8711 26299
rect 17417 26265 17451 26299
rect 19809 26265 19843 26299
rect 20913 26265 20947 26299
rect 24869 26265 24903 26299
rect 8217 26197 8251 26231
rect 12173 26197 12207 26231
rect 12541 26197 12575 26231
rect 14473 26197 14507 26231
rect 2145 25993 2179 26027
rect 8493 25993 8527 26027
rect 9229 25993 9263 26027
rect 10793 25993 10827 26027
rect 10885 25993 10919 26027
rect 15853 25993 15887 26027
rect 19349 25993 19383 26027
rect 20269 25993 20303 26027
rect 20361 25993 20395 26027
rect 22385 25993 22419 26027
rect 22477 25993 22511 26027
rect 23305 25925 23339 25959
rect 2329 25857 2363 25891
rect 3065 25857 3099 25891
rect 4169 25857 4203 25891
rect 8861 25857 8895 25891
rect 9597 25857 9631 25891
rect 12725 25857 12759 25891
rect 15761 25857 15795 25891
rect 17601 25857 17635 25891
rect 23949 25857 23983 25891
rect 3249 25789 3283 25823
rect 8033 25789 8067 25823
rect 9689 25789 9723 25823
rect 9781 25789 9815 25823
rect 10977 25789 11011 25823
rect 11989 25789 12023 25823
rect 13001 25789 13035 25823
rect 14473 25789 14507 25823
rect 16037 25789 16071 25823
rect 17877 25789 17911 25823
rect 20545 25789 20579 25823
rect 21281 25789 21315 25823
rect 22661 25789 22695 25823
rect 25145 25789 25179 25823
rect 3433 25721 3467 25755
rect 4629 25721 4663 25755
rect 10425 25721 10459 25755
rect 14841 25721 14875 25755
rect 19901 25721 19935 25755
rect 23489 25721 23523 25755
rect 4261 25653 4295 25687
rect 15393 25653 15427 25687
rect 21005 25653 21039 25687
rect 22017 25653 22051 25687
rect 7100 25449 7134 25483
rect 8953 25449 8987 25483
rect 11437 25449 11471 25483
rect 14749 25449 14783 25483
rect 18061 25449 18095 25483
rect 23121 25449 23155 25483
rect 25145 25449 25179 25483
rect 25513 25449 25547 25483
rect 10057 25381 10091 25415
rect 22109 25381 22143 25415
rect 6837 25313 6871 25347
rect 8585 25313 8619 25347
rect 9413 25313 9447 25347
rect 10609 25313 10643 25347
rect 11989 25313 12023 25347
rect 13185 25313 13219 25347
rect 15301 25313 15335 25347
rect 15945 25313 15979 25347
rect 16221 25313 16255 25347
rect 19901 25313 19935 25347
rect 20085 25313 20119 25347
rect 22569 25313 22603 25347
rect 22661 25313 22695 25347
rect 4052 25245 4086 25279
rect 10517 25245 10551 25279
rect 11805 25245 11839 25279
rect 18245 25245 18279 25279
rect 19809 25245 19843 25279
rect 22477 25245 22511 25279
rect 23857 25245 23891 25279
rect 24685 25245 24719 25279
rect 10425 25177 10459 25211
rect 13093 25177 13127 25211
rect 24041 25177 24075 25211
rect 4123 25109 4157 25143
rect 11069 25109 11103 25143
rect 11897 25109 11931 25143
rect 12633 25109 12667 25143
rect 13001 25109 13035 25143
rect 15117 25109 15151 25143
rect 15209 25109 15243 25143
rect 17693 25109 17727 25143
rect 19441 25109 19475 25143
rect 23305 25109 23339 25143
rect 24777 25109 24811 25143
rect 5457 24905 5491 24939
rect 8033 24905 8067 24939
rect 15209 24905 15243 24939
rect 16865 24905 16899 24939
rect 17233 24905 17267 24939
rect 18429 24905 18463 24939
rect 19901 24905 19935 24939
rect 20637 24905 20671 24939
rect 9229 24837 9263 24871
rect 12081 24837 12115 24871
rect 23213 24837 23247 24871
rect 5733 24769 5767 24803
rect 7389 24769 7423 24803
rect 10057 24769 10091 24803
rect 12173 24769 12207 24803
rect 13829 24769 13863 24803
rect 15301 24769 15335 24803
rect 16497 24769 16531 24803
rect 18521 24769 18555 24803
rect 25329 24769 25363 24803
rect 3709 24701 3743 24735
rect 3985 24701 4019 24735
rect 8125 24701 8159 24735
rect 8217 24701 8251 24735
rect 9321 24701 9355 24735
rect 9413 24701 9447 24735
rect 12265 24701 12299 24735
rect 13921 24701 13955 24735
rect 14105 24701 14139 24735
rect 15393 24701 15427 24735
rect 17325 24701 17359 24735
rect 17509 24701 17543 24735
rect 18613 24701 18647 24735
rect 20729 24701 20763 24735
rect 20821 24701 20855 24735
rect 22937 24701 22971 24735
rect 24685 24701 24719 24735
rect 7665 24633 7699 24667
rect 11713 24633 11747 24667
rect 13093 24633 13127 24667
rect 13461 24633 13495 24667
rect 25145 24633 25179 24667
rect 8861 24565 8895 24599
rect 12725 24565 12759 24599
rect 13001 24565 13035 24599
rect 14841 24565 14875 24599
rect 18061 24565 18095 24599
rect 20269 24565 20303 24599
rect 3249 24361 3283 24395
rect 3433 24361 3467 24395
rect 5733 24361 5767 24395
rect 6193 24361 6227 24395
rect 8769 24361 8803 24395
rect 13737 24361 13771 24395
rect 4261 24225 4295 24259
rect 6653 24225 6687 24259
rect 10057 24225 10091 24259
rect 11253 24225 11287 24259
rect 11345 24225 11379 24259
rect 12541 24225 12575 24259
rect 13185 24225 13219 24259
rect 14289 24225 14323 24259
rect 16865 24225 16899 24259
rect 17049 24225 17083 24259
rect 19717 24225 19751 24259
rect 23857 24225 23891 24259
rect 25145 24225 25179 24259
rect 2237 24157 2271 24191
rect 2973 24157 3007 24191
rect 3985 24157 4019 24191
rect 6377 24157 6411 24191
rect 11161 24157 11195 24191
rect 16773 24157 16807 24191
rect 17785 24157 17819 24191
rect 22845 24157 22879 24191
rect 2697 24089 2731 24123
rect 12449 24089 12483 24123
rect 19993 24089 20027 24123
rect 21981 24089 22015 24123
rect 22201 24089 22235 24123
rect 25053 24089 25087 24123
rect 2053 24021 2087 24055
rect 9413 24021 9447 24055
rect 9781 24021 9815 24055
rect 9873 24021 9907 24055
rect 10517 24021 10551 24055
rect 10793 24021 10827 24055
rect 11989 24021 12023 24055
rect 12357 24021 12391 24055
rect 16405 24021 16439 24055
rect 17601 24021 17635 24055
rect 21465 24021 21499 24055
rect 24593 24021 24627 24055
rect 24961 24021 24995 24055
rect 6009 23817 6043 23851
rect 9413 23817 9447 23851
rect 9873 23817 9907 23851
rect 11805 23817 11839 23851
rect 12541 23817 12575 23851
rect 25145 23817 25179 23851
rect 6377 23749 6411 23783
rect 13921 23749 13955 23783
rect 1777 23681 1811 23715
rect 20821 23681 20855 23715
rect 22937 23681 22971 23715
rect 25329 23681 25363 23715
rect 2053 23613 2087 23647
rect 4261 23613 4295 23647
rect 4537 23613 4571 23647
rect 7665 23613 7699 23647
rect 7941 23613 7975 23647
rect 10885 23613 10919 23647
rect 17049 23613 17083 23647
rect 18797 23613 18831 23647
rect 19073 23613 19107 23647
rect 23213 23613 23247 23647
rect 24685 23613 24719 23647
rect 11621 23545 11655 23579
rect 10425 23477 10459 23511
rect 12173 23477 12207 23511
rect 12449 23477 12483 23511
rect 21189 23477 21223 23511
rect 21557 23477 21591 23511
rect 2053 23273 2087 23307
rect 3157 23273 3191 23307
rect 7573 23273 7607 23307
rect 16037 23273 16071 23307
rect 18245 23273 18279 23307
rect 21189 23273 21223 23307
rect 11345 23205 11379 23239
rect 13001 23205 13035 23239
rect 2973 23137 3007 23171
rect 5825 23137 5859 23171
rect 11897 23137 11931 23171
rect 12725 23137 12759 23171
rect 13553 23137 13587 23171
rect 14289 23137 14323 23171
rect 16497 23137 16531 23171
rect 19441 23137 19475 23171
rect 22017 23137 22051 23171
rect 25145 23137 25179 23171
rect 2237 23069 2271 23103
rect 2789 23069 2823 23103
rect 4112 23069 4146 23103
rect 4215 23069 4249 23103
rect 7849 23069 7883 23103
rect 9965 23069 9999 23103
rect 11713 23069 11747 23103
rect 13369 23069 13403 23103
rect 22845 23069 22879 23103
rect 23857 23069 23891 23103
rect 24961 23069 24995 23103
rect 6101 23001 6135 23035
rect 10701 23001 10735 23035
rect 12541 23001 12575 23035
rect 13461 23001 13495 23035
rect 14565 23001 14599 23035
rect 16773 23001 16807 23035
rect 19717 23001 19751 23035
rect 25053 23001 25087 23035
rect 11805 22933 11839 22967
rect 18613 22933 18647 22967
rect 21465 22933 21499 22967
rect 24593 22933 24627 22967
rect 2053 22729 2087 22763
rect 5641 22729 5675 22763
rect 6837 22729 6871 22763
rect 7205 22729 7239 22763
rect 9321 22729 9355 22763
rect 10149 22729 10183 22763
rect 10885 22729 10919 22763
rect 12357 22729 12391 22763
rect 15209 22729 15243 22763
rect 16221 22729 16255 22763
rect 17509 22729 17543 22763
rect 23765 22729 23799 22763
rect 24225 22729 24259 22763
rect 24317 22729 24351 22763
rect 24777 22729 24811 22763
rect 25421 22729 25455 22763
rect 8033 22661 8067 22695
rect 12449 22661 12483 22695
rect 13093 22661 13127 22695
rect 17877 22661 17911 22695
rect 18613 22661 18647 22695
rect 19717 22661 19751 22695
rect 20545 22661 20579 22695
rect 2237 22593 2271 22627
rect 5733 22593 5767 22627
rect 10793 22593 10827 22627
rect 15117 22593 15151 22627
rect 19625 22593 19659 22627
rect 21373 22593 21407 22627
rect 22017 22593 22051 22627
rect 5917 22525 5951 22559
rect 7297 22525 7331 22559
rect 7481 22525 7515 22559
rect 8861 22525 8895 22559
rect 10977 22525 11011 22559
rect 12633 22525 12667 22559
rect 13921 22525 13955 22559
rect 15393 22525 15427 22559
rect 19809 22525 19843 22559
rect 22293 22525 22327 22559
rect 10425 22457 10459 22491
rect 11989 22457 12023 22491
rect 5273 22389 5307 22423
rect 11621 22389 11655 22423
rect 14749 22389 14783 22423
rect 19257 22389 19291 22423
rect 16405 22185 16439 22219
rect 19698 22185 19732 22219
rect 21465 22117 21499 22151
rect 11897 22049 11931 22083
rect 12081 22049 12115 22083
rect 14289 22049 14323 22083
rect 16037 22049 16071 22083
rect 16589 22049 16623 22083
rect 17509 22049 17543 22083
rect 18521 22049 18555 22083
rect 18705 22049 18739 22083
rect 22017 22049 22051 22083
rect 22293 22049 22327 22083
rect 24041 22049 24075 22083
rect 11805 21981 11839 22015
rect 13277 21981 13311 22015
rect 17233 21981 17267 22015
rect 17325 21981 17359 22015
rect 19441 21981 19475 22015
rect 12541 21913 12575 21947
rect 14565 21913 14599 21947
rect 18429 21913 18463 21947
rect 24685 21913 24719 21947
rect 4445 21845 4479 21879
rect 11069 21845 11103 21879
rect 11437 21845 11471 21879
rect 13093 21845 13127 21879
rect 16865 21845 16899 21879
rect 18061 21845 18095 21879
rect 21189 21845 21223 21879
rect 24777 21845 24811 21879
rect 7113 21641 7147 21675
rect 7481 21641 7515 21675
rect 8309 21641 8343 21675
rect 8677 21641 8711 21675
rect 9873 21641 9907 21675
rect 11713 21641 11747 21675
rect 12081 21641 12115 21675
rect 13553 21641 13587 21675
rect 13921 21641 13955 21675
rect 16037 21641 16071 21675
rect 22477 21641 22511 21675
rect 25421 21641 25455 21675
rect 14013 21573 14047 21607
rect 23673 21573 23707 21607
rect 1777 21505 1811 21539
rect 3433 21505 3467 21539
rect 4537 21505 4571 21539
rect 7573 21505 7607 21539
rect 12173 21505 12207 21539
rect 15209 21505 15243 21539
rect 16221 21505 16255 21539
rect 17049 21505 17083 21539
rect 18705 21505 18739 21539
rect 23397 21505 23431 21539
rect 2053 21437 2087 21471
rect 3617 21437 3651 21471
rect 4997 21437 5031 21471
rect 7665 21437 7699 21471
rect 8769 21437 8803 21471
rect 8861 21437 8895 21471
rect 9965 21437 9999 21471
rect 10057 21437 10091 21471
rect 12265 21437 12299 21471
rect 14197 21437 14231 21471
rect 15301 21437 15335 21471
rect 15485 21437 15519 21471
rect 17693 21437 17727 21471
rect 22569 21437 22603 21471
rect 22753 21437 22787 21471
rect 3801 21369 3835 21403
rect 9505 21369 9539 21403
rect 16865 21369 16899 21403
rect 4813 21301 4847 21335
rect 14841 21301 14875 21335
rect 18521 21301 18555 21335
rect 20453 21301 20487 21335
rect 22109 21301 22143 21335
rect 25145 21301 25179 21335
rect 3157 21097 3191 21131
rect 7849 21097 7883 21131
rect 16865 21097 16899 21131
rect 4077 21029 4111 21063
rect 16129 21029 16163 21063
rect 17233 21029 17267 21063
rect 21925 21029 21959 21063
rect 2789 20961 2823 20995
rect 8493 20961 8527 20995
rect 11529 20961 11563 20995
rect 14933 20961 14967 20995
rect 16313 20961 16347 20995
rect 17877 20961 17911 20995
rect 19901 20961 19935 20995
rect 23857 20961 23891 20995
rect 2237 20893 2271 20927
rect 2973 20893 3007 20927
rect 4261 20893 4295 20927
rect 9781 20893 9815 20927
rect 11989 20893 12023 20927
rect 14749 20893 14783 20927
rect 15761 20893 15795 20927
rect 17601 20893 17635 20927
rect 18889 20893 18923 20927
rect 22661 20893 22695 20927
rect 10057 20825 10091 20859
rect 14841 20825 14875 20859
rect 20177 20825 20211 20859
rect 2053 20757 2087 20791
rect 7481 20757 7515 20791
rect 8217 20757 8251 20791
rect 8309 20757 8343 20791
rect 13921 20757 13955 20791
rect 14381 20757 14415 20791
rect 15577 20757 15611 20791
rect 17693 20757 17727 20791
rect 18705 20757 18739 20791
rect 21649 20757 21683 20791
rect 9965 20553 9999 20587
rect 12541 20553 12575 20587
rect 17325 20553 17359 20587
rect 19349 20553 19383 20587
rect 19441 20553 19475 20587
rect 4261 20485 4295 20519
rect 6009 20485 6043 20519
rect 10425 20485 10459 20519
rect 17693 20485 17727 20519
rect 23305 20485 23339 20519
rect 3985 20417 4019 20451
rect 6561 20417 6595 20451
rect 9137 20417 9171 20451
rect 10333 20417 10367 20451
rect 12449 20417 12483 20451
rect 13277 20417 13311 20451
rect 15669 20417 15703 20451
rect 18521 20417 18555 20451
rect 22293 20417 22327 20451
rect 24133 20417 24167 20451
rect 6837 20349 6871 20383
rect 9229 20349 9263 20383
rect 9413 20349 9447 20383
rect 10517 20349 10551 20383
rect 12725 20349 12759 20383
rect 19625 20349 19659 20383
rect 24409 20349 24443 20383
rect 8769 20281 8803 20315
rect 5733 20213 5767 20247
rect 8309 20213 8343 20247
rect 12081 20213 12115 20247
rect 13737 20213 13771 20247
rect 14749 20213 14783 20247
rect 15485 20213 15519 20247
rect 17785 20213 17819 20247
rect 18337 20213 18371 20247
rect 18981 20213 19015 20247
rect 5089 20009 5123 20043
rect 11713 20009 11747 20043
rect 14289 20009 14323 20043
rect 20361 20009 20395 20043
rect 15393 19941 15427 19975
rect 5733 19873 5767 19907
rect 6009 19873 6043 19907
rect 9137 19873 9171 19907
rect 11161 19873 11195 19907
rect 12265 19873 12299 19907
rect 14841 19873 14875 19907
rect 23857 19873 23891 19907
rect 5273 19805 5307 19839
rect 7757 19805 7791 19839
rect 8401 19805 8435 19839
rect 12081 19805 12115 19839
rect 14657 19805 14691 19839
rect 17233 19805 17267 19839
rect 17785 19805 17819 19839
rect 18705 19805 18739 19839
rect 22017 19805 22051 19839
rect 22845 19805 22879 19839
rect 9413 19737 9447 19771
rect 13829 19737 13863 19771
rect 14749 19737 14783 19771
rect 17325 19737 17359 19771
rect 17969 19737 18003 19771
rect 22201 19737 22235 19771
rect 7481 19669 7515 19703
rect 8677 19669 8711 19703
rect 12173 19669 12207 19703
rect 18521 19669 18555 19703
rect 19349 19669 19383 19703
rect 2053 19465 2087 19499
rect 4261 19465 4295 19499
rect 8769 19465 8803 19499
rect 9229 19465 9263 19499
rect 11713 19465 11747 19499
rect 13921 19465 13955 19499
rect 16865 19465 16899 19499
rect 17877 19465 17911 19499
rect 19441 19465 19475 19499
rect 19809 19465 19843 19499
rect 19901 19465 19935 19499
rect 21189 19465 21223 19499
rect 23765 19465 23799 19499
rect 18797 19397 18831 19431
rect 2237 19329 2271 19363
rect 4445 19329 4479 19363
rect 6561 19329 6595 19363
rect 9137 19329 9171 19363
rect 12081 19329 12115 19363
rect 14013 19329 14047 19363
rect 17049 19329 17083 19363
rect 21097 19329 21131 19363
rect 6837 19261 6871 19295
rect 9321 19261 9355 19295
rect 12173 19261 12207 19295
rect 12265 19261 12299 19295
rect 14197 19261 14231 19295
rect 14565 19261 14599 19295
rect 17969 19261 18003 19295
rect 18153 19261 18187 19295
rect 20085 19261 20119 19295
rect 21373 19261 21407 19295
rect 22017 19261 22051 19295
rect 22293 19261 22327 19295
rect 13553 19193 13587 19227
rect 17509 19193 17543 19227
rect 8309 19125 8343 19159
rect 10885 19125 10919 19159
rect 11069 19125 11103 19159
rect 11253 19125 11287 19159
rect 13185 19125 13219 19159
rect 18889 19125 18923 19159
rect 20729 19125 20763 19159
rect 24041 19125 24075 19159
rect 8401 18921 8435 18955
rect 12173 18921 12207 18955
rect 14289 18921 14323 18955
rect 18337 18921 18371 18955
rect 18981 18921 19015 18955
rect 24041 18921 24075 18955
rect 24409 18921 24443 18955
rect 18613 18853 18647 18887
rect 2053 18785 2087 18819
rect 13461 18785 13495 18819
rect 13553 18785 13587 18819
rect 14841 18785 14875 18819
rect 17969 18785 18003 18819
rect 1777 18717 1811 18751
rect 9781 18717 9815 18751
rect 11897 18717 11931 18751
rect 14657 18717 14691 18751
rect 16221 18717 16255 18751
rect 19625 18717 19659 18751
rect 20361 18717 20395 18751
rect 21557 18717 21591 18751
rect 22293 18717 22327 18751
rect 10057 18649 10091 18683
rect 14749 18649 14783 18683
rect 16497 18649 16531 18683
rect 21189 18649 21223 18683
rect 22569 18649 22603 18683
rect 8585 18581 8619 18615
rect 9413 18581 9447 18615
rect 11529 18581 11563 18615
rect 13001 18581 13035 18615
rect 13369 18581 13403 18615
rect 19717 18581 19751 18615
rect 7757 18377 7791 18411
rect 10425 18377 10459 18411
rect 10793 18377 10827 18411
rect 14289 18377 14323 18411
rect 14657 18377 14691 18411
rect 15393 18377 15427 18411
rect 9321 18309 9355 18343
rect 12081 18309 12115 18343
rect 13921 18309 13955 18343
rect 17233 18309 17267 18343
rect 17509 18309 17543 18343
rect 19165 18309 19199 18343
rect 7665 18241 7699 18275
rect 8493 18241 8527 18275
rect 14749 18241 14783 18275
rect 21281 18241 21315 18275
rect 22109 18241 22143 18275
rect 24041 18241 24075 18275
rect 7849 18173 7883 18207
rect 10885 18173 10919 18207
rect 11069 18173 11103 18207
rect 12173 18173 12207 18207
rect 12265 18173 12299 18207
rect 13553 18173 13587 18207
rect 13829 18173 13863 18207
rect 14933 18173 14967 18207
rect 18337 18173 18371 18207
rect 18889 18173 18923 18207
rect 23305 18173 23339 18207
rect 24777 18173 24811 18207
rect 6929 18105 6963 18139
rect 11713 18105 11747 18139
rect 21465 18105 21499 18139
rect 7297 18037 7331 18071
rect 9781 18037 9815 18071
rect 10057 18037 10091 18071
rect 20637 18037 20671 18071
rect 6285 17833 6319 17867
rect 9137 17833 9171 17867
rect 21649 17833 21683 17867
rect 23857 17833 23891 17867
rect 8677 17765 8711 17799
rect 12725 17765 12759 17799
rect 17233 17765 17267 17799
rect 6837 17697 6871 17731
rect 7941 17697 7975 17731
rect 8125 17697 8159 17731
rect 9689 17697 9723 17731
rect 12449 17697 12483 17731
rect 13461 17697 13495 17731
rect 13645 17697 13679 17731
rect 14749 17697 14783 17731
rect 14841 17697 14875 17731
rect 16681 17697 16715 17731
rect 16865 17697 16899 17731
rect 22109 17697 22143 17731
rect 22385 17697 22419 17731
rect 10517 17629 10551 17663
rect 14657 17629 14691 17663
rect 15577 17629 15611 17663
rect 19901 17629 19935 17663
rect 24869 17629 24903 17663
rect 6653 17561 6687 17595
rect 11345 17561 11379 17595
rect 13369 17561 13403 17595
rect 20177 17561 20211 17595
rect 6745 17493 6779 17527
rect 7481 17493 7515 17527
rect 7849 17493 7883 17527
rect 9505 17493 9539 17527
rect 9597 17493 9631 17527
rect 11897 17493 11931 17527
rect 13001 17493 13035 17527
rect 14289 17493 14323 17527
rect 15669 17493 15703 17527
rect 16221 17493 16255 17527
rect 16589 17493 16623 17527
rect 24133 17493 24167 17527
rect 24685 17493 24719 17527
rect 10057 17289 10091 17323
rect 10425 17289 10459 17323
rect 14381 17289 14415 17323
rect 14841 17289 14875 17323
rect 22109 17221 22143 17255
rect 6561 17153 6595 17187
rect 9045 17153 9079 17187
rect 17049 17153 17083 17187
rect 17693 17153 17727 17187
rect 19809 17153 19843 17187
rect 20913 17153 20947 17187
rect 21557 17153 21591 17187
rect 22845 17153 22879 17187
rect 23949 17153 23983 17187
rect 6837 17085 6871 17119
rect 8585 17085 8619 17119
rect 10517 17085 10551 17119
rect 10701 17085 10735 17119
rect 12633 17085 12667 17119
rect 12909 17085 12943 17119
rect 14933 17085 14967 17119
rect 17969 17085 18003 17119
rect 19441 17085 19475 17119
rect 20453 17085 20487 17119
rect 24685 17085 24719 17119
rect 22293 17017 22327 17051
rect 23029 17017 23063 17051
rect 9229 16949 9263 16983
rect 9505 16949 9539 16983
rect 16037 16949 16071 16983
rect 16865 16949 16899 16983
rect 5628 16745 5662 16779
rect 7113 16745 7147 16779
rect 7481 16745 7515 16779
rect 8769 16745 8803 16779
rect 5365 16609 5399 16643
rect 9689 16609 9723 16643
rect 11069 16609 11103 16643
rect 12265 16609 12299 16643
rect 12357 16609 12391 16643
rect 15761 16609 15795 16643
rect 15945 16609 15979 16643
rect 20637 16609 20671 16643
rect 22017 16609 22051 16643
rect 23765 16609 23799 16643
rect 1593 16541 1627 16575
rect 9505 16541 9539 16575
rect 10885 16541 10919 16575
rect 12173 16541 12207 16575
rect 20453 16541 20487 16575
rect 20545 16541 20579 16575
rect 21741 16541 21775 16575
rect 2513 16473 2547 16507
rect 9137 16405 9171 16439
rect 9597 16405 9631 16439
rect 10517 16405 10551 16439
rect 10977 16405 11011 16439
rect 11805 16405 11839 16439
rect 15301 16405 15335 16439
rect 15669 16405 15703 16439
rect 16405 16405 16439 16439
rect 20085 16405 20119 16439
rect 23489 16405 23523 16439
rect 8953 16201 8987 16235
rect 10149 16201 10183 16235
rect 10609 16201 10643 16235
rect 11713 16201 11747 16235
rect 13737 16201 13771 16235
rect 16405 16201 16439 16235
rect 18613 16201 18647 16235
rect 19257 16201 19291 16235
rect 2513 16133 2547 16167
rect 9321 16133 9355 16167
rect 12081 16133 12115 16167
rect 15945 16133 15979 16167
rect 17141 16133 17175 16167
rect 19717 16133 19751 16167
rect 6653 16065 6687 16099
rect 10517 16065 10551 16099
rect 12173 16065 12207 16099
rect 14197 16065 14231 16099
rect 14657 16065 14691 16099
rect 16865 16065 16899 16099
rect 18889 16065 18923 16099
rect 19625 16065 19659 16099
rect 20453 16065 20487 16099
rect 21281 16065 21315 16099
rect 22385 16065 22419 16099
rect 23397 16065 23431 16099
rect 24133 16065 24167 16099
rect 6929 15997 6963 16031
rect 8401 15997 8435 16031
rect 9413 15997 9447 16031
rect 9505 15997 9539 16031
rect 10701 15997 10735 16031
rect 12265 15997 12299 16031
rect 19901 15997 19935 16031
rect 22477 15997 22511 16031
rect 22661 15997 22695 16031
rect 24777 15997 24811 16031
rect 21465 15929 21499 15963
rect 2605 15861 2639 15895
rect 13001 15861 13035 15895
rect 14289 15861 14323 15895
rect 16037 15861 16071 15895
rect 22017 15861 22051 15895
rect 23213 15861 23247 15895
rect 8493 15657 8527 15691
rect 14289 15657 14323 15691
rect 13645 15589 13679 15623
rect 17325 15589 17359 15623
rect 21097 15589 21131 15623
rect 11069 15521 11103 15555
rect 14841 15521 14875 15555
rect 17877 15521 17911 15555
rect 20085 15521 20119 15555
rect 13461 15453 13495 15487
rect 14657 15453 14691 15487
rect 17785 15453 17819 15487
rect 18337 15453 18371 15487
rect 19901 15453 19935 15487
rect 20821 15453 20855 15487
rect 22845 15453 22879 15487
rect 11345 15385 11379 15419
rect 21833 15385 21867 15419
rect 23857 15385 23891 15419
rect 12817 15317 12851 15351
rect 14749 15317 14783 15351
rect 17693 15317 17727 15351
rect 18705 15317 18739 15351
rect 19441 15317 19475 15351
rect 19809 15317 19843 15351
rect 20637 15317 20671 15351
rect 21925 15317 21959 15351
rect 11529 15113 11563 15147
rect 13001 15113 13035 15147
rect 14197 15113 14231 15147
rect 18797 15113 18831 15147
rect 18889 15113 18923 15147
rect 22293 15113 22327 15147
rect 9413 15045 9447 15079
rect 11161 15045 11195 15079
rect 13461 15045 13495 15079
rect 17233 15045 17267 15079
rect 17693 15045 17727 15079
rect 13369 14977 13403 15011
rect 14565 14977 14599 15011
rect 14657 14977 14691 15011
rect 15669 14977 15703 15011
rect 16221 14977 16255 15011
rect 19809 14977 19843 15011
rect 23949 14977 23983 15011
rect 9137 14909 9171 14943
rect 13645 14909 13679 14943
rect 14841 14909 14875 14943
rect 15301 14909 15335 14943
rect 18981 14909 19015 14943
rect 24685 14909 24719 14943
rect 15853 14841 15887 14875
rect 17325 14773 17359 14807
rect 18429 14773 18463 14807
rect 19625 14773 19659 14807
rect 13001 14569 13035 14603
rect 17141 14569 17175 14603
rect 11989 14501 12023 14535
rect 14105 14501 14139 14535
rect 9965 14433 9999 14467
rect 13461 14433 13495 14467
rect 13553 14433 13587 14467
rect 15393 14433 15427 14467
rect 21189 14433 21223 14467
rect 12725 14365 12759 14399
rect 18245 14365 18279 14399
rect 18613 14365 18647 14399
rect 20913 14365 20947 14399
rect 10241 14297 10275 14331
rect 13369 14297 13403 14331
rect 15669 14297 15703 14331
rect 18797 14297 18831 14331
rect 11713 14229 11747 14263
rect 17509 14229 17543 14263
rect 19441 14229 19475 14263
rect 19993 14229 20027 14263
rect 22661 14229 22695 14263
rect 22937 14229 22971 14263
rect 12265 14025 12299 14059
rect 12725 14025 12759 14059
rect 21833 14025 21867 14059
rect 23029 14025 23063 14059
rect 10057 13957 10091 13991
rect 13553 13957 13587 13991
rect 14013 13957 14047 13991
rect 17417 13957 17451 13991
rect 19717 13957 19751 13991
rect 21373 13957 21407 13991
rect 25145 13957 25179 13991
rect 1777 13889 1811 13923
rect 8033 13889 8067 13923
rect 12633 13889 12667 13923
rect 17141 13889 17175 13923
rect 20453 13889 20487 13923
rect 21189 13889 21223 13923
rect 23213 13889 23247 13923
rect 23949 13889 23983 13923
rect 2053 13821 2087 13855
rect 9781 13821 9815 13855
rect 12817 13821 12851 13855
rect 13737 13821 13771 13855
rect 18889 13821 18923 13855
rect 19257 13821 19291 13855
rect 19901 13821 19935 13855
rect 20637 13821 20671 13855
rect 8296 13685 8330 13719
rect 11621 13481 11655 13515
rect 11989 13481 12023 13515
rect 12357 13481 12391 13515
rect 13461 13481 13495 13515
rect 16313 13481 16347 13515
rect 20729 13481 20763 13515
rect 9045 13413 9079 13447
rect 6837 13345 6871 13379
rect 7113 13345 7147 13379
rect 9873 13345 9907 13379
rect 10149 13345 10183 13379
rect 12909 13345 12943 13379
rect 14565 13345 14599 13379
rect 18245 13345 18279 13379
rect 18429 13345 18463 13379
rect 19901 13345 19935 13379
rect 19993 13345 20027 13379
rect 12817 13277 12851 13311
rect 18797 13277 18831 13311
rect 19809 13277 19843 13311
rect 22661 13277 22695 13311
rect 12725 13209 12759 13243
rect 14841 13209 14875 13243
rect 18153 13209 18187 13243
rect 23857 13209 23891 13243
rect 8585 13141 8619 13175
rect 16865 13141 16899 13175
rect 17785 13141 17819 13175
rect 19441 13141 19475 13175
rect 21557 13141 21591 13175
rect 8677 12937 8711 12971
rect 11161 12937 11195 12971
rect 15853 12937 15887 12971
rect 16497 12937 16531 12971
rect 17233 12937 17267 12971
rect 21465 12937 21499 12971
rect 11621 12869 11655 12903
rect 14473 12869 14507 12903
rect 14933 12869 14967 12903
rect 15393 12869 15427 12903
rect 17325 12869 17359 12903
rect 18981 12869 19015 12903
rect 8585 12801 8619 12835
rect 9413 12801 9447 12835
rect 13737 12801 13771 12835
rect 18521 12801 18555 12835
rect 22845 12801 22879 12835
rect 23949 12801 23983 12835
rect 8769 12733 8803 12767
rect 9689 12733 9723 12767
rect 17417 12733 17451 12767
rect 19717 12733 19751 12767
rect 19993 12733 20027 12767
rect 22017 12733 22051 12767
rect 24777 12733 24811 12767
rect 13921 12665 13955 12699
rect 14657 12665 14691 12699
rect 15577 12665 15611 12699
rect 8217 12597 8251 12631
rect 16865 12597 16899 12631
rect 18613 12597 18647 12631
rect 22661 12597 22695 12631
rect 14105 12393 14139 12427
rect 14473 12393 14507 12427
rect 15669 12393 15703 12427
rect 18889 12393 18923 12427
rect 20453 12325 20487 12359
rect 11805 12257 11839 12291
rect 15117 12257 15151 12291
rect 16221 12257 16255 12291
rect 17141 12257 17175 12291
rect 17417 12257 17451 12291
rect 21557 12257 21591 12291
rect 21741 12257 21775 12291
rect 11529 12189 11563 12223
rect 16037 12189 16071 12223
rect 20637 12189 20671 12223
rect 21465 12189 21499 12223
rect 23397 12189 23431 12223
rect 13645 12121 13679 12155
rect 14841 12121 14875 12155
rect 13277 12053 13311 12087
rect 13921 12053 13955 12087
rect 14933 12053 14967 12087
rect 16129 12053 16163 12087
rect 19349 12053 19383 12087
rect 21097 12053 21131 12087
rect 23213 12053 23247 12087
rect 14565 11849 14599 11883
rect 16129 11849 16163 11883
rect 17509 11849 17543 11883
rect 19993 11849 20027 11883
rect 15485 11781 15519 11815
rect 16957 11781 16991 11815
rect 18521 11781 18555 11815
rect 20913 11781 20947 11815
rect 21373 11781 21407 11815
rect 25145 11781 25179 11815
rect 12817 11713 12851 11747
rect 15393 11713 15427 11747
rect 18245 11713 18279 11747
rect 23949 11713 23983 11747
rect 13093 11645 13127 11679
rect 15577 11645 15611 11679
rect 21097 11577 21131 11611
rect 15025 11509 15059 11543
rect 17049 11509 17083 11543
rect 20361 11509 20395 11543
rect 15485 11305 15519 11339
rect 14749 11169 14783 11203
rect 16037 11169 16071 11203
rect 15945 11101 15979 11135
rect 15853 11033 15887 11067
rect 20821 11033 20855 11067
rect 21005 11033 21039 11067
rect 19625 10965 19659 10999
rect 19533 10761 19567 10795
rect 20361 10761 20395 10795
rect 12081 10625 12115 10659
rect 14841 10625 14875 10659
rect 18429 10625 18463 10659
rect 20545 10625 20579 10659
rect 23397 10625 23431 10659
rect 23949 10625 23983 10659
rect 19625 10557 19659 10591
rect 19809 10557 19843 10591
rect 24777 10557 24811 10591
rect 12265 10489 12299 10523
rect 14657 10489 14691 10523
rect 18245 10421 18279 10455
rect 19165 10421 19199 10455
rect 23213 10421 23247 10455
rect 21281 10149 21315 10183
rect 14657 10013 14691 10047
rect 14841 10013 14875 10047
rect 21465 10013 21499 10047
rect 22201 10013 22235 10047
rect 22661 10013 22695 10047
rect 23857 10013 23891 10047
rect 16773 9945 16807 9979
rect 24685 9945 24719 9979
rect 16865 9877 16899 9911
rect 22017 9877 22051 9911
rect 24777 9877 24811 9911
rect 16957 9605 16991 9639
rect 19073 9605 19107 9639
rect 5825 9537 5859 9571
rect 6929 9537 6963 9571
rect 22937 9537 22971 9571
rect 23949 9537 23983 9571
rect 7021 9469 7055 9503
rect 7113 9469 7147 9503
rect 24685 9469 24719 9503
rect 6561 9401 6595 9435
rect 17141 9401 17175 9435
rect 19257 9401 19291 9435
rect 22753 9333 22787 9367
rect 24685 9061 24719 9095
rect 21741 8925 21775 8959
rect 23949 8925 23983 8959
rect 24869 8925 24903 8959
rect 21557 8789 21591 8823
rect 23765 8789 23799 8823
rect 19165 8517 19199 8551
rect 20729 8517 20763 8551
rect 25145 8517 25179 8551
rect 22293 8449 22327 8483
rect 23949 8449 23983 8483
rect 20913 8381 20947 8415
rect 22569 8381 22603 8415
rect 19349 8313 19383 8347
rect 6469 8041 6503 8075
rect 4077 7905 4111 7939
rect 23397 7905 23431 7939
rect 20453 7837 20487 7871
rect 21281 7837 21315 7871
rect 22845 7837 22879 7871
rect 24869 7837 24903 7871
rect 4353 7769 4387 7803
rect 6101 7769 6135 7803
rect 20269 7701 20303 7735
rect 21097 7701 21131 7735
rect 24685 7701 24719 7735
rect 18797 7429 18831 7463
rect 25145 7429 25179 7463
rect 20269 7361 20303 7395
rect 22109 7361 22143 7395
rect 23949 7361 23983 7395
rect 21281 7293 21315 7327
rect 22569 7293 22603 7327
rect 18981 7225 19015 7259
rect 19717 6749 19751 6783
rect 20821 6749 20855 6783
rect 22845 6749 22879 6783
rect 22017 6681 22051 6715
rect 23857 6681 23891 6715
rect 19533 6613 19567 6647
rect 21281 6341 21315 6375
rect 25145 6341 25179 6375
rect 18429 6273 18463 6307
rect 20269 6273 20303 6307
rect 22109 6273 22143 6307
rect 24041 6273 24075 6307
rect 19257 6205 19291 6239
rect 22477 6205 22511 6239
rect 24777 5865 24811 5899
rect 21005 5729 21039 5763
rect 22845 5729 22879 5763
rect 20545 5661 20579 5695
rect 22385 5661 22419 5695
rect 24685 5661 24719 5695
rect 18797 5253 18831 5287
rect 17785 5185 17819 5219
rect 19533 5185 19567 5219
rect 22017 5185 22051 5219
rect 24133 5185 24167 5219
rect 19901 5117 19935 5151
rect 22477 5117 22511 5151
rect 24777 5117 24811 5151
rect 24869 4709 24903 4743
rect 19901 4641 19935 4675
rect 21741 4641 21775 4675
rect 23213 4641 23247 4675
rect 23489 4641 23523 4675
rect 17693 4573 17727 4607
rect 19441 4573 19475 4607
rect 21281 4573 21315 4607
rect 24685 4573 24719 4607
rect 18705 4505 18739 4539
rect 1777 4097 1811 4131
rect 13553 4097 13587 4131
rect 16129 4097 16163 4131
rect 16865 4097 16899 4131
rect 18705 4097 18739 4131
rect 22109 4097 22143 4131
rect 23857 4097 23891 4131
rect 11345 4029 11379 4063
rect 11713 4029 11747 4063
rect 11989 4029 12023 4063
rect 14013 4029 14047 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 22477 4029 22511 4063
rect 24317 4029 24351 4063
rect 1593 3961 1627 3995
rect 9965 3961 9999 3995
rect 16313 3961 16347 3995
rect 2053 3893 2087 3927
rect 6377 3893 6411 3927
rect 9505 3893 9539 3927
rect 9781 3893 9815 3927
rect 11069 3893 11103 3927
rect 5273 3689 5307 3723
rect 6745 3689 6779 3723
rect 8217 3689 8251 3723
rect 9321 3689 9355 3723
rect 10057 3689 10091 3723
rect 1777 3621 1811 3655
rect 5917 3621 5951 3655
rect 7573 3553 7607 3587
rect 11253 3553 11287 3587
rect 12817 3553 12851 3587
rect 15485 3553 15519 3587
rect 17325 3553 17359 3587
rect 19901 3553 19935 3587
rect 21741 3553 21775 3587
rect 1961 3485 1995 3519
rect 2421 3485 2455 3519
rect 5089 3485 5123 3519
rect 6101 3485 6135 3519
rect 6561 3485 6595 3519
rect 8033 3485 8067 3519
rect 9137 3485 9171 3519
rect 9873 3485 9907 3519
rect 10517 3485 10551 3519
rect 10977 3485 11011 3519
rect 12449 3485 12483 3519
rect 15117 3485 15151 3519
rect 16865 3485 16899 3519
rect 19441 3485 19475 3519
rect 21281 3485 21315 3519
rect 3157 3417 3191 3451
rect 2237 3349 2271 3383
rect 2881 3349 2915 3383
rect 3249 3349 3283 3383
rect 3617 3349 3651 3383
rect 4813 3349 4847 3383
rect 7205 3349 7239 3383
rect 7757 3349 7791 3383
rect 8677 3349 8711 3383
rect 10701 3349 10735 3383
rect 25421 3349 25455 3383
rect 2697 3145 2731 3179
rect 5181 3145 5215 3179
rect 5917 3145 5951 3179
rect 7021 3145 7055 3179
rect 7757 3145 7791 3179
rect 8493 3145 8527 3179
rect 11897 3145 11931 3179
rect 24869 3145 24903 3179
rect 23581 3077 23615 3111
rect 1869 3009 1903 3043
rect 2513 3009 2547 3043
rect 3525 3009 3559 3043
rect 4721 3009 4755 3043
rect 4997 3009 5031 3043
rect 5733 3009 5767 3043
rect 6837 3009 6871 3043
rect 7573 3009 7607 3043
rect 8309 3009 8343 3043
rect 9321 3009 9355 3043
rect 10609 3009 10643 3043
rect 11713 3009 11747 3043
rect 12633 3009 12667 3043
rect 14289 3009 14323 3043
rect 16865 3009 16899 3043
rect 18705 3009 18739 3043
rect 3249 2941 3283 2975
rect 9045 2941 9079 2975
rect 10333 2941 10367 2975
rect 13369 2941 13403 2975
rect 14749 2941 14783 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 2053 2873 2087 2907
rect 1501 2805 1535 2839
rect 4353 2805 4387 2839
rect 6469 2805 6503 2839
rect 1869 2601 1903 2635
rect 2605 2601 2639 2635
rect 4169 2601 4203 2635
rect 7113 2601 7147 2635
rect 9781 2601 9815 2635
rect 3341 2533 3375 2567
rect 4997 2465 5031 2499
rect 7941 2465 7975 2499
rect 10609 2465 10643 2499
rect 14105 2465 14139 2499
rect 15209 2465 15243 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 22477 2465 22511 2499
rect 1685 2397 1719 2431
rect 2421 2397 2455 2431
rect 3157 2397 3191 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 5825 2397 5859 2431
rect 6469 2397 6503 2431
rect 6929 2397 6963 2431
rect 7665 2397 7699 2431
rect 9137 2397 9171 2431
rect 9597 2397 9631 2431
rect 10333 2397 10367 2431
rect 11897 2397 11931 2431
rect 12541 2397 12575 2431
rect 14657 2397 14691 2431
rect 16865 2397 16899 2431
rect 19441 2397 19475 2431
rect 22017 2397 22051 2431
rect 25329 2397 25363 2431
rect 6101 2329 6135 2363
rect 6653 2329 6687 2363
rect 9321 2329 9355 2363
rect 13553 2329 13587 2363
rect 11713 2261 11747 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 9950 54272 9956 54324
rect 10008 54272 10014 54324
rect 14553 54315 14611 54321
rect 14553 54281 14565 54315
rect 14599 54312 14611 54315
rect 14734 54312 14740 54324
rect 14599 54284 14740 54312
rect 14599 54281 14611 54284
rect 14553 54275 14611 54281
rect 14734 54272 14740 54284
rect 14792 54272 14798 54324
rect 16206 54272 16212 54324
rect 16264 54312 16270 54324
rect 16393 54315 16451 54321
rect 16393 54312 16405 54315
rect 16264 54284 16405 54312
rect 16264 54272 16270 54284
rect 16393 54281 16405 54284
rect 16439 54312 16451 54315
rect 16439 54284 16574 54312
rect 16439 54281 16451 54284
rect 16393 54275 16451 54281
rect 5813 54247 5871 54253
rect 5813 54213 5825 54247
rect 5859 54244 5871 54247
rect 7834 54244 7840 54256
rect 5859 54216 7840 54244
rect 5859 54213 5871 54216
rect 5813 54207 5871 54213
rect 7834 54204 7840 54216
rect 7892 54204 7898 54256
rect 8389 54247 8447 54253
rect 8389 54213 8401 54247
rect 8435 54244 8447 54247
rect 9968 54244 9996 54272
rect 8435 54216 9996 54244
rect 10965 54247 11023 54253
rect 8435 54213 8447 54216
rect 8389 54207 8447 54213
rect 10965 54213 10977 54247
rect 11011 54244 11023 54247
rect 11422 54244 11428 54256
rect 11011 54216 11428 54244
rect 11011 54213 11023 54216
rect 10965 54207 11023 54213
rect 11422 54204 11428 54216
rect 11480 54204 11486 54256
rect 12894 54244 12900 54256
rect 11900 54216 12900 54244
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 4522 54176 4528 54188
rect 2271 54148 4528 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 4522 54136 4528 54148
rect 4580 54136 4586 54188
rect 4614 54136 4620 54188
rect 4672 54136 4678 54188
rect 7377 54179 7435 54185
rect 7377 54145 7389 54179
rect 7423 54145 7435 54179
rect 7377 54139 7435 54145
rect 3237 54111 3295 54117
rect 3237 54077 3249 54111
rect 3283 54108 3295 54111
rect 5902 54108 5908 54120
rect 3283 54080 5908 54108
rect 3283 54077 3295 54080
rect 3237 54071 3295 54077
rect 5902 54068 5908 54080
rect 5960 54068 5966 54120
rect 7392 54108 7420 54139
rect 9950 54136 9956 54188
rect 10008 54136 10014 54188
rect 11900 54185 11928 54216
rect 12894 54204 12900 54216
rect 12952 54244 12958 54256
rect 14093 54247 14151 54253
rect 14093 54244 14105 54247
rect 12952 54216 14105 54244
rect 12952 54204 12958 54216
rect 14093 54213 14105 54216
rect 14139 54213 14151 54247
rect 14093 54207 14151 54213
rect 11885 54179 11943 54185
rect 11885 54145 11897 54179
rect 11931 54145 11943 54179
rect 11885 54139 11943 54145
rect 12342 54136 12348 54188
rect 12400 54136 12406 54188
rect 14752 54176 14780 54272
rect 14829 54179 14887 54185
rect 14829 54176 14841 54179
rect 14752 54148 14841 54176
rect 14829 54145 14841 54148
rect 14875 54145 14887 54179
rect 14829 54139 14887 54145
rect 15194 54136 15200 54188
rect 15252 54176 15258 54188
rect 15565 54179 15623 54185
rect 15565 54176 15577 54179
rect 15252 54148 15577 54176
rect 15252 54136 15258 54148
rect 15565 54145 15577 54148
rect 15611 54176 15623 54179
rect 16117 54179 16175 54185
rect 16117 54176 16129 54179
rect 15611 54148 16129 54176
rect 15611 54145 15623 54148
rect 15565 54139 15623 54145
rect 16117 54145 16129 54148
rect 16163 54145 16175 54179
rect 16546 54176 16574 54284
rect 24486 54272 24492 54324
rect 24544 54272 24550 54324
rect 17678 54204 17684 54256
rect 17736 54244 17742 54256
rect 18417 54247 18475 54253
rect 18417 54244 18429 54247
rect 17736 54216 18429 54244
rect 17736 54204 17742 54216
rect 18417 54213 18429 54216
rect 18463 54244 18475 54247
rect 18874 54244 18880 54256
rect 18463 54216 18880 54244
rect 18463 54213 18475 54216
rect 18417 54207 18475 54213
rect 18874 54204 18880 54216
rect 18932 54204 18938 54256
rect 21453 54247 21511 54253
rect 21453 54244 21465 54247
rect 20180 54216 21465 54244
rect 16853 54179 16911 54185
rect 16853 54176 16865 54179
rect 16546 54148 16865 54176
rect 16117 54139 16175 54145
rect 16853 54145 16865 54148
rect 16899 54145 16911 54179
rect 16853 54139 16911 54145
rect 16942 54136 16948 54188
rect 17000 54176 17006 54188
rect 17589 54179 17647 54185
rect 17589 54176 17601 54179
rect 17000 54148 17601 54176
rect 17000 54136 17006 54148
rect 17589 54145 17601 54148
rect 17635 54176 17647 54179
rect 18969 54179 19027 54185
rect 18969 54176 18981 54179
rect 17635 54148 18981 54176
rect 17635 54145 17647 54148
rect 17589 54139 17647 54145
rect 18969 54145 18981 54148
rect 19015 54145 19027 54179
rect 18969 54139 19027 54145
rect 19429 54179 19487 54185
rect 19429 54145 19441 54179
rect 19475 54145 19487 54179
rect 19429 54139 19487 54145
rect 11238 54108 11244 54120
rect 7392 54080 11244 54108
rect 11238 54068 11244 54080
rect 11296 54068 11302 54120
rect 12526 54068 12532 54120
rect 12584 54108 12590 54120
rect 12805 54111 12863 54117
rect 12805 54108 12817 54111
rect 12584 54080 12817 54108
rect 12584 54068 12590 54080
rect 12805 54077 12817 54080
rect 12851 54077 12863 54111
rect 12805 54071 12863 54077
rect 18414 54068 18420 54120
rect 18472 54108 18478 54120
rect 19444 54108 19472 54139
rect 19518 54136 19524 54188
rect 19576 54176 19582 54188
rect 20180 54185 20208 54216
rect 21453 54213 21465 54216
rect 21499 54213 21511 54247
rect 23293 54247 23351 54253
rect 23293 54244 23305 54247
rect 21453 54207 21511 54213
rect 22020 54216 23305 54244
rect 20165 54179 20223 54185
rect 20165 54176 20177 54179
rect 19576 54148 20177 54176
rect 19576 54136 19582 54148
rect 20165 54145 20177 54148
rect 20211 54145 20223 54179
rect 20165 54139 20223 54145
rect 20714 54136 20720 54188
rect 20772 54176 20778 54188
rect 20901 54179 20959 54185
rect 20901 54176 20913 54179
rect 20772 54148 20913 54176
rect 20772 54136 20778 54148
rect 20901 54145 20913 54148
rect 20947 54145 20959 54179
rect 20901 54139 20959 54145
rect 21358 54136 21364 54188
rect 21416 54176 21422 54188
rect 22020 54185 22048 54216
rect 23293 54213 23305 54216
rect 23339 54213 23351 54247
rect 23293 54207 23351 54213
rect 22005 54179 22063 54185
rect 22005 54176 22017 54179
rect 21416 54148 22017 54176
rect 21416 54136 21422 54148
rect 22005 54145 22017 54148
rect 22051 54145 22063 54179
rect 22005 54139 22063 54145
rect 22462 54136 22468 54188
rect 22520 54176 22526 54188
rect 22741 54179 22799 54185
rect 22741 54176 22753 54179
rect 22520 54148 22753 54176
rect 22520 54136 22526 54148
rect 22741 54145 22753 54148
rect 22787 54145 22799 54179
rect 22741 54139 22799 54145
rect 23753 54179 23811 54185
rect 23753 54145 23765 54179
rect 23799 54176 23811 54179
rect 24504 54176 24532 54272
rect 23799 54148 24532 54176
rect 23799 54145 23811 54148
rect 23753 54139 23811 54145
rect 24946 54136 24952 54188
rect 25004 54136 25010 54188
rect 19702 54108 19708 54120
rect 18472 54080 19708 54108
rect 18472 54068 18478 54080
rect 19702 54068 19708 54080
rect 19760 54068 19766 54120
rect 15378 54000 15384 54052
rect 15436 54040 15442 54052
rect 17773 54043 17831 54049
rect 17773 54040 17785 54043
rect 15436 54012 17785 54040
rect 15436 54000 15442 54012
rect 17773 54009 17785 54012
rect 17819 54009 17831 54043
rect 17773 54003 17831 54009
rect 25130 54000 25136 54052
rect 25188 54000 25194 54052
rect 11698 53932 11704 53984
rect 11756 53932 11762 53984
rect 14090 53932 14096 53984
rect 14148 53972 14154 53984
rect 15013 53975 15071 53981
rect 15013 53972 15025 53975
rect 14148 53944 15025 53972
rect 14148 53932 14154 53944
rect 15013 53941 15025 53944
rect 15059 53941 15071 53975
rect 15013 53935 15071 53941
rect 15286 53932 15292 53984
rect 15344 53972 15350 53984
rect 15749 53975 15807 53981
rect 15749 53972 15761 53975
rect 15344 53944 15761 53972
rect 15344 53932 15350 53944
rect 15749 53941 15761 53944
rect 15795 53941 15807 53975
rect 15749 53935 15807 53941
rect 17034 53932 17040 53984
rect 17092 53932 17098 53984
rect 18506 53932 18512 53984
rect 18564 53932 18570 53984
rect 19334 53932 19340 53984
rect 19392 53972 19398 53984
rect 19613 53975 19671 53981
rect 19613 53972 19625 53975
rect 19392 53944 19625 53972
rect 19392 53932 19398 53944
rect 19613 53941 19625 53944
rect 19659 53941 19671 53975
rect 19613 53935 19671 53941
rect 20349 53975 20407 53981
rect 20349 53941 20361 53975
rect 20395 53972 20407 53975
rect 20898 53972 20904 53984
rect 20395 53944 20904 53972
rect 20395 53941 20407 53944
rect 20349 53935 20407 53941
rect 20898 53932 20904 53944
rect 20956 53932 20962 53984
rect 21085 53975 21143 53981
rect 21085 53941 21097 53975
rect 21131 53972 21143 53975
rect 21542 53972 21548 53984
rect 21131 53944 21548 53972
rect 21131 53941 21143 53944
rect 21085 53935 21143 53941
rect 21542 53932 21548 53944
rect 21600 53932 21606 53984
rect 22186 53932 22192 53984
rect 22244 53932 22250 53984
rect 22738 53932 22744 53984
rect 22796 53972 22802 53984
rect 22925 53975 22983 53981
rect 22925 53972 22937 53975
rect 22796 53944 22937 53972
rect 22796 53932 22802 53944
rect 22925 53941 22937 53944
rect 22971 53941 22983 53975
rect 22925 53935 22983 53941
rect 23937 53975 23995 53981
rect 23937 53941 23949 53975
rect 23983 53972 23995 53975
rect 24118 53972 24124 53984
rect 23983 53944 24124 53972
rect 23983 53941 23995 53944
rect 23937 53935 23995 53941
rect 24118 53932 24124 53944
rect 24176 53932 24182 53984
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 16393 53771 16451 53777
rect 16393 53737 16405 53771
rect 16439 53768 16451 53771
rect 16574 53768 16580 53780
rect 16439 53740 16580 53768
rect 16439 53737 16451 53740
rect 16393 53731 16451 53737
rect 16574 53728 16580 53740
rect 16632 53728 16638 53780
rect 18874 53728 18880 53780
rect 18932 53728 18938 53780
rect 5534 53660 5540 53712
rect 5592 53660 5598 53712
rect 21269 53703 21327 53709
rect 21269 53669 21281 53703
rect 21315 53700 21327 53703
rect 21634 53700 21640 53712
rect 21315 53672 21640 53700
rect 21315 53669 21327 53672
rect 21269 53663 21327 53669
rect 21634 53660 21640 53672
rect 21692 53660 21698 53712
rect 22370 53660 22376 53712
rect 22428 53700 22434 53712
rect 23109 53703 23167 53709
rect 23109 53700 23121 53703
rect 22428 53672 23121 53700
rect 22428 53660 22434 53672
rect 23109 53669 23121 53672
rect 23155 53669 23167 53703
rect 23109 53663 23167 53669
rect 3237 53635 3295 53641
rect 3237 53601 3249 53635
rect 3283 53632 3295 53635
rect 5552 53632 5580 53660
rect 3283 53604 5580 53632
rect 6549 53635 6607 53641
rect 3283 53601 3295 53604
rect 3237 53595 3295 53601
rect 6549 53601 6561 53635
rect 6595 53632 6607 53635
rect 7374 53632 7380 53644
rect 6595 53604 7380 53632
rect 6595 53601 6607 53604
rect 6549 53595 6607 53601
rect 7374 53592 7380 53604
rect 7432 53592 7438 53644
rect 8389 53635 8447 53641
rect 8389 53601 8401 53635
rect 8435 53632 8447 53635
rect 8846 53632 8852 53644
rect 8435 53604 8852 53632
rect 8435 53601 8447 53604
rect 8389 53595 8447 53601
rect 8846 53592 8852 53604
rect 8904 53592 8910 53644
rect 11054 53592 11060 53644
rect 11112 53592 11118 53644
rect 12158 53592 12164 53644
rect 12216 53632 12222 53644
rect 12713 53635 12771 53641
rect 12713 53632 12725 53635
rect 12216 53604 12725 53632
rect 12216 53592 12222 53604
rect 12713 53601 12725 53604
rect 12759 53601 12771 53635
rect 24397 53635 24455 53641
rect 24397 53632 24409 53635
rect 12713 53595 12771 53601
rect 23308 53604 24409 53632
rect 2225 53567 2283 53573
rect 2225 53533 2237 53567
rect 2271 53564 2283 53567
rect 5537 53567 5595 53573
rect 2271 53536 4476 53564
rect 2271 53533 2283 53536
rect 2225 53527 2283 53533
rect 4448 53496 4476 53536
rect 5537 53533 5549 53567
rect 5583 53564 5595 53567
rect 6822 53564 6828 53576
rect 5583 53536 6828 53564
rect 5583 53533 5595 53536
rect 5537 53527 5595 53533
rect 6822 53524 6828 53536
rect 6880 53524 6886 53576
rect 7285 53567 7343 53573
rect 7285 53533 7297 53567
rect 7331 53564 7343 53567
rect 9122 53564 9128 53576
rect 7331 53536 9128 53564
rect 7331 53533 7343 53536
rect 7285 53527 7343 53533
rect 9122 53524 9128 53536
rect 9180 53524 9186 53576
rect 10410 53524 10416 53576
rect 10468 53524 10474 53576
rect 12437 53567 12495 53573
rect 12437 53533 12449 53567
rect 12483 53564 12495 53567
rect 12618 53564 12624 53576
rect 12483 53536 12624 53564
rect 12483 53533 12495 53536
rect 12437 53527 12495 53533
rect 12618 53524 12624 53536
rect 12676 53524 12682 53576
rect 13998 53524 14004 53576
rect 14056 53564 14062 53576
rect 14277 53567 14335 53573
rect 14277 53564 14289 53567
rect 14056 53536 14289 53564
rect 14056 53524 14062 53536
rect 14277 53533 14289 53536
rect 14323 53564 14335 53567
rect 14829 53567 14887 53573
rect 14829 53564 14841 53567
rect 14323 53536 14841 53564
rect 14323 53533 14335 53536
rect 14277 53527 14335 53533
rect 14829 53533 14841 53536
rect 14875 53533 14887 53567
rect 14829 53527 14887 53533
rect 15470 53524 15476 53576
rect 15528 53564 15534 53576
rect 15657 53567 15715 53573
rect 15657 53564 15669 53567
rect 15528 53536 15669 53564
rect 15528 53524 15534 53536
rect 15657 53533 15669 53536
rect 15703 53564 15715 53567
rect 16117 53567 16175 53573
rect 16117 53564 16129 53567
rect 15703 53536 16129 53564
rect 15703 53533 15715 53536
rect 15657 53527 15715 53533
rect 16117 53533 16129 53536
rect 16163 53533 16175 53567
rect 16117 53527 16175 53533
rect 16574 53524 16580 53576
rect 16632 53564 16638 53576
rect 16669 53567 16727 53573
rect 16669 53564 16681 53567
rect 16632 53536 16681 53564
rect 16632 53524 16638 53536
rect 16669 53533 16681 53536
rect 16715 53533 16727 53567
rect 16669 53527 16727 53533
rect 17310 53524 17316 53576
rect 17368 53564 17374 53576
rect 17589 53567 17647 53573
rect 17589 53564 17601 53567
rect 17368 53536 17601 53564
rect 17368 53524 17374 53536
rect 17589 53533 17601 53536
rect 17635 53533 17647 53567
rect 17589 53527 17647 53533
rect 18233 53567 18291 53573
rect 18233 53533 18245 53567
rect 18279 53564 18291 53567
rect 18322 53564 18328 53576
rect 18279 53536 18328 53564
rect 18279 53533 18291 53536
rect 18233 53527 18291 53533
rect 18322 53524 18328 53536
rect 18380 53564 18386 53576
rect 18693 53567 18751 53573
rect 18693 53564 18705 53567
rect 18380 53536 18705 53564
rect 18380 53524 18386 53536
rect 18693 53533 18705 53536
rect 18739 53533 18751 53567
rect 18693 53527 18751 53533
rect 19150 53524 19156 53576
rect 19208 53564 19214 53576
rect 19429 53567 19487 53573
rect 19429 53564 19441 53567
rect 19208 53536 19441 53564
rect 19208 53524 19214 53536
rect 19429 53533 19441 53536
rect 19475 53533 19487 53567
rect 19429 53527 19487 53533
rect 19886 53524 19892 53576
rect 19944 53564 19950 53576
rect 20257 53567 20315 53573
rect 20257 53564 20269 53567
rect 19944 53536 20269 53564
rect 19944 53524 19950 53536
rect 20257 53533 20269 53536
rect 20303 53564 20315 53567
rect 20717 53567 20775 53573
rect 20717 53564 20729 53567
rect 20303 53536 20729 53564
rect 20303 53533 20315 53536
rect 20257 53527 20315 53533
rect 20717 53533 20729 53536
rect 20763 53533 20775 53567
rect 20717 53527 20775 53533
rect 20990 53524 20996 53576
rect 21048 53564 21054 53576
rect 21085 53567 21143 53573
rect 21085 53564 21097 53567
rect 21048 53536 21097 53564
rect 21048 53524 21054 53536
rect 21085 53533 21097 53536
rect 21131 53533 21143 53567
rect 21085 53527 21143 53533
rect 21726 53524 21732 53576
rect 21784 53564 21790 53576
rect 22005 53567 22063 53573
rect 22005 53564 22017 53567
rect 21784 53536 22017 53564
rect 21784 53524 21790 53536
rect 22005 53533 22017 53536
rect 22051 53533 22063 53567
rect 22005 53527 22063 53533
rect 22094 53524 22100 53576
rect 22152 53564 22158 53576
rect 22649 53567 22707 53573
rect 22649 53564 22661 53567
rect 22152 53536 22661 53564
rect 22152 53524 22158 53536
rect 22649 53533 22661 53536
rect 22695 53533 22707 53567
rect 22649 53527 22707 53533
rect 22830 53524 22836 53576
rect 22888 53564 22894 53576
rect 23308 53573 23336 53604
rect 24397 53601 24409 53604
rect 24443 53601 24455 53635
rect 24397 53595 24455 53601
rect 23293 53567 23351 53573
rect 23293 53564 23305 53567
rect 22888 53536 23305 53564
rect 22888 53524 22894 53536
rect 23293 53533 23305 53536
rect 23339 53533 23351 53567
rect 23293 53527 23351 53533
rect 23382 53524 23388 53576
rect 23440 53564 23446 53576
rect 23845 53567 23903 53573
rect 23845 53564 23857 53567
rect 23440 53536 23857 53564
rect 23440 53524 23446 53536
rect 23845 53533 23857 53536
rect 23891 53564 23903 53567
rect 24581 53567 24639 53573
rect 24581 53564 24593 53567
rect 23891 53536 24593 53564
rect 23891 53533 23903 53536
rect 23845 53527 23903 53533
rect 24581 53533 24593 53536
rect 24627 53533 24639 53567
rect 24581 53527 24639 53533
rect 24762 53524 24768 53576
rect 24820 53564 24826 53576
rect 25041 53567 25099 53573
rect 25041 53564 25053 53567
rect 24820 53536 25053 53564
rect 24820 53524 24826 53536
rect 25041 53533 25053 53536
rect 25087 53533 25099 53567
rect 25041 53527 25099 53533
rect 7374 53496 7380 53508
rect 4448 53468 7380 53496
rect 7374 53456 7380 53468
rect 7432 53456 7438 53508
rect 15841 53499 15899 53505
rect 15841 53465 15853 53499
rect 15887 53496 15899 53499
rect 16390 53496 16396 53508
rect 15887 53468 16396 53496
rect 15887 53465 15899 53468
rect 15841 53459 15899 53465
rect 16390 53456 16396 53468
rect 16448 53456 16454 53508
rect 20438 53456 20444 53508
rect 20496 53456 20502 53508
rect 24029 53499 24087 53505
rect 24029 53465 24041 53499
rect 24075 53496 24087 53499
rect 24210 53496 24216 53508
rect 24075 53468 24216 53496
rect 24075 53465 24087 53468
rect 24029 53459 24087 53465
rect 24210 53456 24216 53468
rect 24268 53456 24274 53508
rect 14458 53388 14464 53440
rect 14516 53388 14522 53440
rect 16850 53388 16856 53440
rect 16908 53388 16914 53440
rect 17402 53388 17408 53440
rect 17460 53388 17466 53440
rect 18322 53388 18328 53440
rect 18380 53388 18386 53440
rect 19610 53388 19616 53440
rect 19668 53388 19674 53440
rect 21358 53388 21364 53440
rect 21416 53428 21422 53440
rect 21821 53431 21879 53437
rect 21821 53428 21833 53431
rect 21416 53400 21833 53428
rect 21416 53388 21422 53400
rect 21821 53397 21833 53400
rect 21867 53397 21879 53431
rect 21821 53391 21879 53397
rect 22462 53388 22468 53440
rect 22520 53388 22526 53440
rect 25225 53431 25283 53437
rect 25225 53397 25237 53431
rect 25271 53428 25283 53431
rect 25866 53428 25872 53440
rect 25271 53400 25872 53428
rect 25271 53397 25283 53400
rect 25225 53391 25283 53397
rect 25866 53388 25872 53400
rect 25924 53388 25930 53440
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 2133 53227 2191 53233
rect 2133 53193 2145 53227
rect 2179 53224 2191 53227
rect 2774 53224 2780 53236
rect 2179 53196 2780 53224
rect 2179 53193 2191 53196
rect 2133 53187 2191 53193
rect 1765 53091 1823 53097
rect 1765 53057 1777 53091
rect 1811 53088 1823 53091
rect 2148 53088 2176 53187
rect 2774 53184 2780 53196
rect 2832 53184 2838 53236
rect 17310 53184 17316 53236
rect 17368 53184 17374 53236
rect 19150 53184 19156 53236
rect 19208 53224 19214 53236
rect 19521 53227 19579 53233
rect 19521 53224 19533 53227
rect 19208 53196 19533 53224
rect 19208 53184 19214 53196
rect 19521 53193 19533 53196
rect 19567 53193 19579 53227
rect 19521 53187 19579 53193
rect 19702 53184 19708 53236
rect 19760 53184 19766 53236
rect 20990 53184 20996 53236
rect 21048 53184 21054 53236
rect 21726 53184 21732 53236
rect 21784 53224 21790 53236
rect 21821 53227 21879 53233
rect 21821 53224 21833 53227
rect 21784 53196 21833 53224
rect 21784 53184 21790 53196
rect 21821 53193 21833 53196
rect 21867 53193 21879 53227
rect 21821 53187 21879 53193
rect 22094 53184 22100 53236
rect 22152 53224 22158 53236
rect 22281 53227 22339 53233
rect 22281 53224 22293 53227
rect 22152 53196 22293 53224
rect 22152 53184 22158 53196
rect 22281 53193 22293 53196
rect 22327 53193 22339 53227
rect 22281 53187 22339 53193
rect 22554 53184 22560 53236
rect 22612 53184 22618 53236
rect 23017 53227 23075 53233
rect 23017 53193 23029 53227
rect 23063 53224 23075 53227
rect 23290 53224 23296 53236
rect 23063 53196 23296 53224
rect 23063 53193 23075 53196
rect 23017 53187 23075 53193
rect 23290 53184 23296 53196
rect 23348 53184 23354 53236
rect 3973 53159 4031 53165
rect 3973 53125 3985 53159
rect 4019 53156 4031 53159
rect 4430 53156 4436 53168
rect 4019 53128 4436 53156
rect 4019 53125 4031 53128
rect 3973 53119 4031 53125
rect 4430 53116 4436 53128
rect 4488 53116 4494 53168
rect 5813 53159 5871 53165
rect 5813 53125 5825 53159
rect 5859 53156 5871 53159
rect 6270 53156 6276 53168
rect 5859 53128 6276 53156
rect 5859 53125 5871 53128
rect 5813 53119 5871 53125
rect 6270 53116 6276 53128
rect 6328 53116 6334 53168
rect 9125 53159 9183 53165
rect 9125 53125 9137 53159
rect 9171 53156 9183 53159
rect 9214 53156 9220 53168
rect 9171 53128 9220 53156
rect 9171 53125 9183 53128
rect 9125 53119 9183 53125
rect 9214 53116 9220 53128
rect 9272 53116 9278 53168
rect 13630 53116 13636 53168
rect 13688 53156 13694 53168
rect 13817 53159 13875 53165
rect 13817 53156 13829 53159
rect 13688 53128 13829 53156
rect 13688 53116 13694 53128
rect 13817 53125 13829 53128
rect 13863 53125 13875 53159
rect 13817 53119 13875 53125
rect 20714 53116 20720 53168
rect 20772 53156 20778 53168
rect 21177 53159 21235 53165
rect 21177 53156 21189 53159
rect 20772 53128 21189 53156
rect 20772 53116 20778 53128
rect 21177 53125 21189 53128
rect 21223 53125 21235 53159
rect 21177 53119 21235 53125
rect 1811 53060 2176 53088
rect 2961 53091 3019 53097
rect 1811 53057 1823 53060
rect 1765 53051 1823 53057
rect 2961 53057 2973 53091
rect 3007 53057 3019 53091
rect 2961 53051 3019 53057
rect 4801 53091 4859 53097
rect 4801 53057 4813 53091
rect 4847 53088 4859 53091
rect 6362 53088 6368 53100
rect 4847 53060 6368 53088
rect 4847 53057 4859 53060
rect 4801 53051 4859 53057
rect 2976 53020 3004 53051
rect 6362 53048 6368 53060
rect 6420 53048 6426 53100
rect 8113 53091 8171 53097
rect 8113 53057 8125 53091
rect 8159 53057 8171 53091
rect 8113 53051 8171 53057
rect 5626 53020 5632 53032
rect 2976 52992 5632 53020
rect 5626 52980 5632 52992
rect 5684 52980 5690 53032
rect 8128 53020 8156 53051
rect 9674 53048 9680 53100
rect 9732 53088 9738 53100
rect 9769 53091 9827 53097
rect 9769 53088 9781 53091
rect 9732 53060 9781 53088
rect 9732 53048 9738 53060
rect 9769 53057 9781 53060
rect 9815 53057 9827 53091
rect 9769 53051 9827 53057
rect 11882 53048 11888 53100
rect 11940 53048 11946 53100
rect 14366 53048 14372 53100
rect 14424 53088 14430 53100
rect 14645 53091 14703 53097
rect 14645 53088 14657 53091
rect 14424 53060 14657 53088
rect 14424 53048 14430 53060
rect 14645 53057 14657 53060
rect 14691 53088 14703 53091
rect 14921 53091 14979 53097
rect 14921 53088 14933 53091
rect 14691 53060 14933 53088
rect 14691 53057 14703 53060
rect 14645 53051 14703 53057
rect 14921 53057 14933 53060
rect 14967 53057 14979 53091
rect 14921 53051 14979 53057
rect 15838 53048 15844 53100
rect 15896 53088 15902 53100
rect 16117 53091 16175 53097
rect 16117 53088 16129 53091
rect 15896 53060 16129 53088
rect 15896 53048 15902 53060
rect 16117 53057 16129 53060
rect 16163 53088 16175 53091
rect 16393 53091 16451 53097
rect 16393 53088 16405 53091
rect 16163 53060 16405 53088
rect 16163 53057 16175 53060
rect 16117 53051 16175 53057
rect 16393 53057 16405 53060
rect 16439 53057 16451 53091
rect 16393 53051 16451 53057
rect 18782 53048 18788 53100
rect 18840 53088 18846 53100
rect 19061 53091 19119 53097
rect 19061 53088 19073 53091
rect 18840 53060 19073 53088
rect 18840 53048 18846 53060
rect 19061 53057 19073 53060
rect 19107 53088 19119 53091
rect 19337 53091 19395 53097
rect 19337 53088 19349 53091
rect 19107 53060 19349 53088
rect 19107 53057 19119 53060
rect 19061 53051 19119 53057
rect 19337 53057 19349 53060
rect 19383 53057 19395 53091
rect 19337 53051 19395 53057
rect 20254 53048 20260 53100
rect 20312 53088 20318 53100
rect 20533 53091 20591 53097
rect 20533 53088 20545 53091
rect 20312 53060 20545 53088
rect 20312 53048 20318 53060
rect 20533 53057 20545 53060
rect 20579 53088 20591 53091
rect 20809 53091 20867 53097
rect 20809 53088 20821 53091
rect 20579 53060 20821 53088
rect 20579 53057 20591 53060
rect 20533 53051 20591 53057
rect 20809 53057 20821 53060
rect 20855 53057 20867 53091
rect 23308 53088 23336 53184
rect 23477 53091 23535 53097
rect 23477 53088 23489 53091
rect 23308 53060 23489 53088
rect 20809 53051 20867 53057
rect 23477 53057 23489 53060
rect 23523 53057 23535 53091
rect 23477 53051 23535 53057
rect 23566 53048 23572 53100
rect 23624 53088 23630 53100
rect 24121 53091 24179 53097
rect 24121 53088 24133 53091
rect 23624 53060 24133 53088
rect 23624 53048 23630 53060
rect 24121 53057 24133 53060
rect 24167 53088 24179 53091
rect 24397 53091 24455 53097
rect 24397 53088 24409 53091
rect 24167 53060 24409 53088
rect 24167 53057 24179 53060
rect 24121 53051 24179 53057
rect 24397 53057 24409 53060
rect 24443 53057 24455 53091
rect 24397 53051 24455 53057
rect 24765 53091 24823 53097
rect 24765 53057 24777 53091
rect 24811 53088 24823 53091
rect 25038 53088 25044 53100
rect 24811 53060 25044 53088
rect 24811 53057 24823 53060
rect 24765 53051 24823 53057
rect 25038 53048 25044 53060
rect 25096 53048 25102 53100
rect 10226 53020 10232 53032
rect 8128 52992 10232 53020
rect 10226 52980 10232 52992
rect 10284 52980 10290 53032
rect 10318 52980 10324 53032
rect 10376 52980 10382 53032
rect 11790 52980 11796 53032
rect 11848 53020 11854 53032
rect 12345 53023 12403 53029
rect 12345 53020 12357 53023
rect 11848 52992 12357 53020
rect 11848 52980 11854 52992
rect 12345 52989 12357 52992
rect 12391 52989 12403 53023
rect 12345 52983 12403 52989
rect 1581 52955 1639 52961
rect 1581 52921 1593 52955
rect 1627 52952 1639 52955
rect 3970 52952 3976 52964
rect 1627 52924 3976 52952
rect 1627 52921 1639 52924
rect 1581 52915 1639 52921
rect 3970 52912 3976 52924
rect 4028 52912 4034 52964
rect 13998 52912 14004 52964
rect 14056 52912 14062 52964
rect 1854 52844 1860 52896
rect 1912 52884 1918 52896
rect 3510 52884 3516 52896
rect 1912 52856 3516 52884
rect 1912 52844 1918 52856
rect 3510 52844 3516 52856
rect 3568 52844 3574 52896
rect 14458 52844 14464 52896
rect 14516 52844 14522 52896
rect 15930 52844 15936 52896
rect 15988 52844 15994 52896
rect 18598 52844 18604 52896
rect 18656 52884 18662 52896
rect 18877 52887 18935 52893
rect 18877 52884 18889 52887
rect 18656 52856 18889 52884
rect 18656 52844 18662 52856
rect 18877 52853 18889 52856
rect 18923 52853 18935 52887
rect 18877 52847 18935 52853
rect 20162 52844 20168 52896
rect 20220 52884 20226 52896
rect 20349 52887 20407 52893
rect 20349 52884 20361 52887
rect 20220 52856 20361 52884
rect 20220 52844 20226 52856
rect 20349 52853 20361 52856
rect 20395 52853 20407 52887
rect 20349 52847 20407 52853
rect 22186 52844 22192 52896
rect 22244 52884 22250 52896
rect 23293 52887 23351 52893
rect 23293 52884 23305 52887
rect 22244 52856 23305 52884
rect 22244 52844 22250 52856
rect 23293 52853 23305 52856
rect 23339 52853 23351 52887
rect 23293 52847 23351 52853
rect 23934 52844 23940 52896
rect 23992 52844 23998 52896
rect 25222 52844 25228 52896
rect 25280 52844 25286 52896
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 2222 52640 2228 52692
rect 2280 52680 2286 52692
rect 3418 52680 3424 52692
rect 2280 52652 3424 52680
rect 2280 52640 2286 52652
rect 3418 52640 3424 52652
rect 3476 52640 3482 52692
rect 12618 52640 12624 52692
rect 12676 52640 12682 52692
rect 13630 52640 13636 52692
rect 13688 52680 13694 52692
rect 14093 52683 14151 52689
rect 14093 52680 14105 52683
rect 13688 52652 14105 52680
rect 13688 52640 13694 52652
rect 14093 52649 14105 52652
rect 14139 52649 14151 52683
rect 14093 52643 14151 52649
rect 24581 52683 24639 52689
rect 24581 52649 24593 52683
rect 24627 52680 24639 52683
rect 24762 52680 24768 52692
rect 24627 52652 24768 52680
rect 24627 52649 24639 52652
rect 24581 52643 24639 52649
rect 24762 52640 24768 52652
rect 24820 52640 24826 52692
rect 1302 52572 1308 52624
rect 1360 52612 1366 52624
rect 3786 52612 3792 52624
rect 1360 52584 3792 52612
rect 1360 52572 1366 52584
rect 3786 52572 3792 52584
rect 3844 52612 3850 52624
rect 25225 52615 25283 52621
rect 3844 52584 4016 52612
rect 3844 52572 3850 52584
rect 3237 52547 3295 52553
rect 3237 52513 3249 52547
rect 3283 52544 3295 52547
rect 3694 52544 3700 52556
rect 3283 52516 3700 52544
rect 3283 52513 3295 52516
rect 3237 52507 3295 52513
rect 3694 52504 3700 52516
rect 3752 52504 3758 52556
rect 3988 52553 4016 52584
rect 25225 52581 25237 52615
rect 25271 52612 25283 52615
rect 25590 52612 25596 52624
rect 25271 52584 25596 52612
rect 25271 52581 25283 52584
rect 25225 52575 25283 52581
rect 25590 52572 25596 52584
rect 25648 52572 25654 52624
rect 3973 52547 4031 52553
rect 3973 52513 3985 52547
rect 4019 52513 4031 52547
rect 4430 52544 4436 52556
rect 3973 52507 4031 52513
rect 4249 52547 4307 52553
rect 4249 52513 4261 52547
rect 4295 52544 4307 52547
rect 4295 52516 7696 52544
rect 4295 52513 4307 52516
rect 4249 52507 4307 52513
rect 2225 52479 2283 52485
rect 2225 52445 2237 52479
rect 2271 52476 2283 52479
rect 5166 52476 5172 52488
rect 2271 52448 5172 52476
rect 2271 52445 2283 52448
rect 2225 52439 2283 52445
rect 5166 52436 5172 52448
rect 5224 52436 5230 52488
rect 5445 52479 5503 52485
rect 5445 52445 5457 52479
rect 5491 52476 5503 52479
rect 5718 52476 5724 52488
rect 5491 52448 5724 52476
rect 5491 52445 5503 52448
rect 5445 52439 5503 52445
rect 5718 52436 5724 52448
rect 5776 52436 5782 52488
rect 6549 52479 6607 52485
rect 6549 52445 6561 52479
rect 6595 52476 6607 52479
rect 6638 52476 6644 52488
rect 6595 52448 6644 52476
rect 6595 52445 6607 52448
rect 6549 52439 6607 52445
rect 6638 52436 6644 52448
rect 6696 52436 6702 52488
rect 7282 52436 7288 52488
rect 7340 52436 7346 52488
rect 7668 52476 7696 52516
rect 7742 52504 7748 52556
rect 7800 52504 7806 52556
rect 10686 52504 10692 52556
rect 10744 52544 10750 52556
rect 11241 52547 11299 52553
rect 11241 52544 11253 52547
rect 10744 52516 11253 52544
rect 10744 52504 10750 52516
rect 11241 52513 11253 52516
rect 11287 52513 11299 52547
rect 11241 52507 11299 52513
rect 8938 52476 8944 52488
rect 7668 52448 8944 52476
rect 8938 52436 8944 52448
rect 8996 52436 9002 52488
rect 10778 52436 10784 52488
rect 10836 52436 10842 52488
rect 12802 52436 12808 52488
rect 12860 52436 12866 52488
rect 13538 52436 13544 52488
rect 13596 52476 13602 52488
rect 13633 52479 13691 52485
rect 13633 52476 13645 52479
rect 13596 52448 13645 52476
rect 13596 52436 13602 52448
rect 13633 52445 13645 52448
rect 13679 52445 13691 52479
rect 13633 52439 13691 52445
rect 24762 52436 24768 52488
rect 24820 52476 24826 52488
rect 25041 52479 25099 52485
rect 25041 52476 25053 52479
rect 24820 52448 25053 52476
rect 24820 52436 24826 52448
rect 25041 52445 25053 52448
rect 25087 52445 25099 52479
rect 25041 52439 25099 52445
rect 13354 52368 13360 52420
rect 13412 52408 13418 52420
rect 13449 52411 13507 52417
rect 13449 52408 13461 52411
rect 13412 52380 13461 52408
rect 13412 52368 13418 52380
rect 13449 52377 13461 52380
rect 13495 52377 13507 52411
rect 13449 52371 13507 52377
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 5626 52096 5632 52148
rect 5684 52136 5690 52148
rect 7009 52139 7067 52145
rect 7009 52136 7021 52139
rect 5684 52108 7021 52136
rect 5684 52096 5690 52108
rect 7009 52105 7021 52108
rect 7055 52105 7067 52139
rect 7009 52099 7067 52105
rect 11701 52139 11759 52145
rect 11701 52105 11713 52139
rect 11747 52136 11759 52139
rect 11882 52136 11888 52148
rect 11747 52108 11888 52136
rect 11747 52105 11759 52108
rect 11701 52099 11759 52105
rect 11882 52096 11888 52108
rect 11940 52096 11946 52148
rect 12342 52096 12348 52148
rect 12400 52096 12406 52148
rect 13265 52139 13323 52145
rect 13265 52105 13277 52139
rect 13311 52136 13323 52139
rect 13354 52136 13360 52148
rect 13311 52108 13360 52136
rect 13311 52105 13323 52108
rect 13265 52099 13323 52105
rect 13354 52096 13360 52108
rect 13412 52096 13418 52148
rect 24946 52096 24952 52148
rect 25004 52136 25010 52148
rect 25225 52139 25283 52145
rect 25225 52136 25237 52139
rect 25004 52108 25237 52136
rect 25004 52096 25010 52108
rect 25225 52105 25237 52108
rect 25271 52105 25283 52139
rect 25225 52099 25283 52105
rect 4890 52068 4896 52080
rect 2976 52040 4896 52068
rect 2976 52009 3004 52040
rect 4890 52028 4896 52040
rect 4948 52028 4954 52080
rect 6917 52071 6975 52077
rect 6917 52037 6929 52071
rect 6963 52068 6975 52071
rect 9030 52068 9036 52080
rect 6963 52040 9036 52068
rect 6963 52037 6975 52040
rect 6917 52031 6975 52037
rect 9030 52028 9036 52040
rect 9088 52028 9094 52080
rect 10134 52068 10140 52080
rect 9140 52040 10140 52068
rect 2961 52003 3019 52009
rect 2961 51969 2973 52003
rect 3007 51969 3019 52003
rect 2961 51963 3019 51969
rect 4706 51960 4712 52012
rect 4764 51960 4770 52012
rect 8021 52003 8079 52009
rect 8021 51969 8033 52003
rect 8067 52000 8079 52003
rect 9140 52000 9168 52040
rect 10134 52028 10140 52040
rect 10192 52028 10198 52080
rect 8067 51972 9168 52000
rect 8067 51969 8079 51972
rect 8021 51963 8079 51969
rect 9766 51960 9772 52012
rect 9824 51960 9830 52012
rect 10870 51960 10876 52012
rect 10928 52000 10934 52012
rect 11885 52003 11943 52009
rect 11885 52000 11897 52003
rect 10928 51972 11897 52000
rect 10928 51960 10934 51972
rect 11885 51969 11897 51972
rect 11931 51969 11943 52003
rect 11885 51963 11943 51969
rect 11974 51960 11980 52012
rect 12032 52000 12038 52012
rect 12529 52003 12587 52009
rect 12529 52000 12541 52003
rect 12032 51972 12541 52000
rect 12032 51960 12038 51972
rect 12529 51969 12541 51972
rect 12575 51969 12587 52003
rect 12529 51963 12587 51969
rect 3326 51892 3332 51944
rect 3384 51892 3390 51944
rect 4798 51892 4804 51944
rect 4856 51932 4862 51944
rect 5077 51935 5135 51941
rect 5077 51932 5089 51935
rect 4856 51904 5089 51932
rect 4856 51892 4862 51904
rect 5077 51901 5089 51904
rect 5123 51901 5135 51935
rect 5077 51895 5135 51901
rect 8478 51892 8484 51944
rect 8536 51892 8542 51944
rect 9858 51892 9864 51944
rect 9916 51932 9922 51944
rect 10137 51935 10195 51941
rect 10137 51932 10149 51935
rect 9916 51904 10149 51932
rect 9916 51892 9922 51904
rect 10137 51901 10149 51904
rect 10183 51901 10195 51935
rect 10137 51895 10195 51901
rect 25498 51756 25504 51808
rect 25556 51756 25562 51808
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 3786 51552 3792 51604
rect 3844 51552 3850 51604
rect 9950 51552 9956 51604
rect 10008 51592 10014 51604
rect 10229 51595 10287 51601
rect 10229 51592 10241 51595
rect 10008 51564 10241 51592
rect 10008 51552 10014 51564
rect 10229 51561 10241 51564
rect 10275 51561 10287 51595
rect 10229 51555 10287 51561
rect 2866 51416 2872 51468
rect 2924 51416 2930 51468
rect 5534 51416 5540 51468
rect 5592 51456 5598 51468
rect 5721 51459 5779 51465
rect 5721 51456 5733 51459
rect 5592 51428 5733 51456
rect 5592 51416 5598 51428
rect 5721 51425 5733 51428
rect 5767 51425 5779 51459
rect 5721 51419 5779 51425
rect 7006 51416 7012 51468
rect 7064 51456 7070 51468
rect 7561 51459 7619 51465
rect 7561 51456 7573 51459
rect 7064 51428 7573 51456
rect 7064 51416 7070 51428
rect 7561 51425 7573 51428
rect 7607 51425 7619 51459
rect 7561 51419 7619 51425
rect 2225 51391 2283 51397
rect 2225 51357 2237 51391
rect 2271 51357 2283 51391
rect 2225 51351 2283 51357
rect 5445 51391 5503 51397
rect 5445 51357 5457 51391
rect 5491 51388 5503 51391
rect 6730 51388 6736 51400
rect 5491 51360 6736 51388
rect 5491 51357 5503 51360
rect 5445 51351 5503 51357
rect 2240 51320 2268 51351
rect 6730 51348 6736 51360
rect 6788 51348 6794 51400
rect 7098 51348 7104 51400
rect 7156 51348 7162 51400
rect 9214 51348 9220 51400
rect 9272 51388 9278 51400
rect 10413 51391 10471 51397
rect 10413 51388 10425 51391
rect 9272 51360 10425 51388
rect 9272 51348 9278 51360
rect 10413 51357 10425 51360
rect 10459 51357 10471 51391
rect 10413 51351 10471 51357
rect 25041 51391 25099 51397
rect 25041 51357 25053 51391
rect 25087 51388 25099 51391
rect 25498 51388 25504 51400
rect 25087 51360 25504 51388
rect 25087 51357 25099 51360
rect 25041 51351 25099 51357
rect 25498 51348 25504 51360
rect 25556 51348 25562 51400
rect 5534 51320 5540 51332
rect 2240 51292 5540 51320
rect 5534 51280 5540 51292
rect 5592 51280 5598 51332
rect 25225 51255 25283 51261
rect 25225 51221 25237 51255
rect 25271 51252 25283 51255
rect 25682 51252 25688 51264
rect 25271 51224 25688 51252
rect 25271 51221 25283 51224
rect 25225 51215 25283 51221
rect 25682 51212 25688 51224
rect 25740 51212 25746 51264
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 5534 51008 5540 51060
rect 5592 51048 5598 51060
rect 6917 51051 6975 51057
rect 6917 51048 6929 51051
rect 5592 51020 6929 51048
rect 5592 51008 5598 51020
rect 6917 51017 6929 51020
rect 6963 51017 6975 51051
rect 6917 51011 6975 51017
rect 4338 50980 4344 50992
rect 2516 50952 4344 50980
rect 2516 50921 2544 50952
rect 4338 50940 4344 50952
rect 4396 50940 4402 50992
rect 4522 50940 4528 50992
rect 4580 50980 4586 50992
rect 9585 50983 9643 50989
rect 4580 50952 7788 50980
rect 4580 50940 4586 50952
rect 2501 50915 2559 50921
rect 2501 50881 2513 50915
rect 2547 50881 2559 50915
rect 2501 50875 2559 50881
rect 4154 50872 4160 50924
rect 4212 50872 4218 50924
rect 6825 50915 6883 50921
rect 6825 50881 6837 50915
rect 6871 50912 6883 50915
rect 7650 50912 7656 50924
rect 6871 50884 7656 50912
rect 6871 50881 6883 50884
rect 6825 50875 6883 50881
rect 7650 50872 7656 50884
rect 7708 50872 7714 50924
rect 7760 50921 7788 50952
rect 9585 50949 9597 50983
rect 9631 50980 9643 50983
rect 10778 50980 10784 50992
rect 9631 50952 10784 50980
rect 9631 50949 9643 50952
rect 9585 50943 9643 50949
rect 10778 50940 10784 50952
rect 10836 50940 10842 50992
rect 7745 50915 7803 50921
rect 7745 50881 7757 50915
rect 7791 50881 7803 50915
rect 7745 50875 7803 50881
rect 7834 50872 7840 50924
rect 7892 50912 7898 50924
rect 9401 50915 9459 50921
rect 9401 50912 9413 50915
rect 7892 50884 9413 50912
rect 7892 50872 7898 50884
rect 9401 50881 9413 50884
rect 9447 50881 9459 50915
rect 9401 50875 9459 50881
rect 24765 50915 24823 50921
rect 24765 50881 24777 50915
rect 24811 50912 24823 50915
rect 25038 50912 25044 50924
rect 24811 50884 25044 50912
rect 24811 50881 24823 50884
rect 24765 50875 24823 50881
rect 25038 50872 25044 50884
rect 25096 50872 25102 50924
rect 2774 50804 2780 50856
rect 2832 50804 2838 50856
rect 4246 50804 4252 50856
rect 4304 50844 4310 50856
rect 4617 50847 4675 50853
rect 4617 50844 4629 50847
rect 4304 50816 4629 50844
rect 4304 50804 4310 50816
rect 4617 50813 4629 50816
rect 4663 50813 4675 50847
rect 4617 50807 4675 50813
rect 7466 50804 7472 50856
rect 7524 50804 7530 50856
rect 15838 50804 15844 50856
rect 15896 50844 15902 50856
rect 16850 50844 16856 50856
rect 15896 50816 16856 50844
rect 15896 50804 15902 50816
rect 16850 50804 16856 50816
rect 16908 50804 16914 50856
rect 25225 50711 25283 50717
rect 25225 50677 25237 50711
rect 25271 50708 25283 50711
rect 25406 50708 25412 50720
rect 25271 50680 25412 50708
rect 25271 50677 25283 50680
rect 25225 50671 25283 50677
rect 25406 50668 25412 50680
rect 25464 50668 25470 50720
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 6822 50464 6828 50516
rect 6880 50464 6886 50516
rect 9122 50464 9128 50516
rect 9180 50504 9186 50516
rect 9217 50507 9275 50513
rect 9217 50504 9229 50507
rect 9180 50476 9229 50504
rect 9180 50464 9186 50476
rect 9217 50473 9229 50476
rect 9263 50473 9275 50507
rect 9217 50467 9275 50473
rect 1302 50328 1308 50380
rect 1360 50368 1366 50380
rect 3973 50371 4031 50377
rect 3973 50368 3985 50371
rect 1360 50340 3985 50368
rect 1360 50328 1366 50340
rect 3973 50337 3985 50340
rect 4019 50368 4031 50371
rect 5077 50371 5135 50377
rect 5077 50368 5089 50371
rect 4019 50340 5089 50368
rect 4019 50337 4031 50340
rect 3973 50331 4031 50337
rect 5077 50337 5089 50340
rect 5123 50337 5135 50371
rect 5077 50331 5135 50337
rect 2225 50303 2283 50309
rect 2225 50269 2237 50303
rect 2271 50269 2283 50303
rect 2225 50263 2283 50269
rect 3237 50303 3295 50309
rect 3237 50269 3249 50303
rect 3283 50300 3295 50303
rect 3418 50300 3424 50312
rect 3283 50272 3424 50300
rect 3283 50269 3295 50272
rect 3237 50263 3295 50269
rect 2240 50164 2268 50263
rect 3418 50260 3424 50272
rect 3476 50260 3482 50312
rect 4249 50303 4307 50309
rect 4249 50269 4261 50303
rect 4295 50269 4307 50303
rect 4249 50263 4307 50269
rect 4264 50232 4292 50263
rect 5810 50260 5816 50312
rect 5868 50300 5874 50312
rect 7009 50303 7067 50309
rect 7009 50300 7021 50303
rect 5868 50272 7021 50300
rect 5868 50260 5874 50272
rect 7009 50269 7021 50272
rect 7055 50269 7067 50303
rect 7009 50263 7067 50269
rect 8386 50260 8392 50312
rect 8444 50300 8450 50312
rect 9401 50303 9459 50309
rect 9401 50300 9413 50303
rect 8444 50272 9413 50300
rect 8444 50260 8450 50272
rect 9401 50269 9413 50272
rect 9447 50269 9459 50303
rect 9401 50263 9459 50269
rect 7558 50232 7564 50244
rect 4264 50204 7564 50232
rect 7558 50192 7564 50204
rect 7616 50192 7622 50244
rect 5074 50164 5080 50176
rect 2240 50136 5080 50164
rect 5074 50124 5080 50136
rect 5132 50124 5138 50176
rect 25314 50124 25320 50176
rect 25372 50164 25378 50176
rect 25409 50167 25467 50173
rect 25409 50164 25421 50167
rect 25372 50136 25421 50164
rect 25372 50124 25378 50136
rect 25409 50133 25421 50136
rect 25455 50133 25467 50167
rect 25409 50127 25467 50133
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 10226 49960 10232 49972
rect 3988 49932 10232 49960
rect 3145 49895 3203 49901
rect 3145 49861 3157 49895
rect 3191 49892 3203 49895
rect 3510 49892 3516 49904
rect 3191 49864 3516 49892
rect 3191 49861 3203 49864
rect 3145 49855 3203 49861
rect 3510 49852 3516 49864
rect 3568 49852 3574 49904
rect 2133 49827 2191 49833
rect 2133 49793 2145 49827
rect 2179 49824 2191 49827
rect 3326 49824 3332 49836
rect 2179 49796 3332 49824
rect 2179 49793 2191 49796
rect 2133 49787 2191 49793
rect 3326 49784 3332 49796
rect 3384 49784 3390 49836
rect 3988 49833 4016 49932
rect 10226 49920 10232 49932
rect 10284 49920 10290 49972
rect 20990 49920 20996 49972
rect 21048 49960 21054 49972
rect 25133 49963 25191 49969
rect 25133 49960 25145 49963
rect 21048 49932 25145 49960
rect 21048 49920 21054 49932
rect 25133 49929 25145 49932
rect 25179 49929 25191 49963
rect 25133 49923 25191 49929
rect 5997 49895 6055 49901
rect 5997 49861 6009 49895
rect 6043 49892 6055 49895
rect 9309 49895 9367 49901
rect 6043 49864 9260 49892
rect 6043 49861 6055 49864
rect 5997 49855 6055 49861
rect 3973 49827 4031 49833
rect 3973 49793 3985 49827
rect 4019 49793 4031 49827
rect 6365 49827 6423 49833
rect 6365 49824 6377 49827
rect 5382 49796 6377 49824
rect 3973 49787 4031 49793
rect 6365 49793 6377 49796
rect 6411 49824 6423 49827
rect 6411 49796 6914 49824
rect 6411 49793 6423 49796
rect 6365 49787 6423 49793
rect 6886 49756 6914 49796
rect 7742 49784 7748 49836
rect 7800 49824 7806 49836
rect 9125 49827 9183 49833
rect 9125 49824 9137 49827
rect 7800 49796 9137 49824
rect 7800 49784 7806 49796
rect 9125 49793 9137 49796
rect 9171 49793 9183 49827
rect 9232 49824 9260 49864
rect 9309 49861 9321 49895
rect 9355 49892 9367 49895
rect 9674 49892 9680 49904
rect 9355 49864 9680 49892
rect 9355 49861 9367 49864
rect 9309 49855 9367 49861
rect 9674 49852 9680 49864
rect 9732 49852 9738 49904
rect 9490 49824 9496 49836
rect 9232 49796 9496 49824
rect 9125 49787 9183 49793
rect 9490 49784 9496 49796
rect 9548 49784 9554 49836
rect 25314 49784 25320 49836
rect 25372 49784 25378 49836
rect 8846 49756 8852 49768
rect 6886 49728 8852 49756
rect 8846 49716 8852 49728
rect 8904 49716 8910 49768
rect 11698 49716 11704 49768
rect 11756 49756 11762 49768
rect 12710 49756 12716 49768
rect 11756 49728 12716 49756
rect 11756 49716 11762 49728
rect 12710 49716 12716 49728
rect 12768 49716 12774 49768
rect 3970 49580 3976 49632
rect 4028 49620 4034 49632
rect 4230 49623 4288 49629
rect 4230 49620 4242 49623
rect 4028 49592 4242 49620
rect 4028 49580 4034 49592
rect 4230 49589 4242 49592
rect 4276 49589 4288 49623
rect 4230 49583 4288 49589
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 11609 49419 11667 49425
rect 11609 49385 11621 49419
rect 11655 49416 11667 49419
rect 11974 49416 11980 49428
rect 11655 49388 11980 49416
rect 11655 49385 11667 49388
rect 11609 49379 11667 49385
rect 11974 49376 11980 49388
rect 12032 49376 12038 49428
rect 1486 49240 1492 49292
rect 1544 49280 1550 49292
rect 2041 49283 2099 49289
rect 2041 49280 2053 49283
rect 1544 49252 2053 49280
rect 1544 49240 1550 49252
rect 2041 49249 2053 49252
rect 2087 49249 2099 49283
rect 2041 49243 2099 49249
rect 1765 49215 1823 49221
rect 1765 49181 1777 49215
rect 1811 49212 1823 49215
rect 10594 49212 10600 49224
rect 1811 49184 10600 49212
rect 1811 49181 1823 49184
rect 1765 49175 1823 49181
rect 10594 49172 10600 49184
rect 10652 49172 10658 49224
rect 10686 49172 10692 49224
rect 10744 49212 10750 49224
rect 11793 49215 11851 49221
rect 11793 49212 11805 49215
rect 10744 49184 11805 49212
rect 10744 49172 10750 49184
rect 11793 49181 11805 49184
rect 11839 49181 11851 49215
rect 11793 49175 11851 49181
rect 24857 49215 24915 49221
rect 24857 49181 24869 49215
rect 24903 49212 24915 49215
rect 25314 49212 25320 49224
rect 24903 49184 25320 49212
rect 24903 49181 24915 49184
rect 24857 49175 24915 49181
rect 25314 49172 25320 49184
rect 25372 49172 25378 49224
rect 25130 49036 25136 49088
rect 25188 49036 25194 49088
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 12713 48875 12771 48881
rect 12713 48841 12725 48875
rect 12759 48872 12771 48875
rect 12802 48872 12808 48884
rect 12759 48844 12808 48872
rect 12759 48841 12771 48844
rect 12713 48835 12771 48841
rect 12802 48832 12808 48844
rect 12860 48832 12866 48884
rect 12526 48696 12532 48748
rect 12584 48736 12590 48748
rect 12897 48739 12955 48745
rect 12897 48736 12909 48739
rect 12584 48708 12909 48736
rect 12584 48696 12590 48708
rect 12897 48705 12909 48708
rect 12943 48705 12955 48739
rect 12897 48699 12955 48705
rect 25501 48535 25559 48541
rect 25501 48501 25513 48535
rect 25547 48532 25559 48535
rect 25774 48532 25780 48544
rect 25547 48504 25780 48532
rect 25547 48501 25559 48504
rect 25501 48495 25559 48501
rect 25774 48492 25780 48504
rect 25832 48492 25838 48544
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 17310 48220 17316 48272
rect 17368 48260 17374 48272
rect 17678 48260 17684 48272
rect 17368 48232 17684 48260
rect 17368 48220 17374 48232
rect 17678 48220 17684 48232
rect 17736 48260 17742 48272
rect 17773 48263 17831 48269
rect 17773 48260 17785 48263
rect 17736 48232 17785 48260
rect 17736 48220 17742 48232
rect 17773 48229 17785 48232
rect 17819 48260 17831 48263
rect 18506 48260 18512 48272
rect 17819 48232 18512 48260
rect 17819 48229 17831 48232
rect 17773 48223 17831 48229
rect 18506 48220 18512 48232
rect 18564 48220 18570 48272
rect 24857 48127 24915 48133
rect 24857 48093 24869 48127
rect 24903 48124 24915 48127
rect 25314 48124 25320 48136
rect 24903 48096 25320 48124
rect 24903 48093 24915 48096
rect 24857 48087 24915 48093
rect 25314 48084 25320 48096
rect 25372 48084 25378 48136
rect 1302 48016 1308 48068
rect 1360 48056 1366 48068
rect 1673 48059 1731 48065
rect 1673 48056 1685 48059
rect 1360 48028 1685 48056
rect 1360 48016 1366 48028
rect 1673 48025 1685 48028
rect 1719 48056 1731 48059
rect 2133 48059 2191 48065
rect 2133 48056 2145 48059
rect 1719 48028 2145 48056
rect 1719 48025 1731 48028
rect 1673 48019 1731 48025
rect 1857 48059 1915 48065
rect 1857 48025 1869 48059
rect 1903 48056 1915 48059
rect 8294 48056 8300 48068
rect 1903 48028 8300 48056
rect 1903 48025 1915 48028
rect 1857 48019 1915 48025
rect 1688 47988 1716 48019
rect 8294 48016 8300 48028
rect 8352 48016 8358 48068
rect 2133 47991 2191 47997
rect 2133 47988 2145 47991
rect 1688 47960 2145 47988
rect 2133 47957 2145 47960
rect 2179 47957 2191 47991
rect 2133 47951 2191 47957
rect 24854 47948 24860 48000
rect 24912 47988 24918 48000
rect 25133 47991 25191 47997
rect 25133 47988 25145 47991
rect 24912 47960 25145 47988
rect 24912 47948 24918 47960
rect 25133 47957 25145 47960
rect 25179 47957 25191 47991
rect 25133 47951 25191 47957
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 9030 47744 9036 47796
rect 9088 47784 9094 47796
rect 9125 47787 9183 47793
rect 9125 47784 9137 47787
rect 9088 47756 9137 47784
rect 9088 47744 9094 47756
rect 9125 47753 9137 47756
rect 9171 47753 9183 47787
rect 9125 47747 9183 47753
rect 15930 47744 15936 47796
rect 15988 47784 15994 47796
rect 17221 47787 17279 47793
rect 17221 47784 17233 47787
rect 15988 47756 17233 47784
rect 15988 47744 15994 47756
rect 17221 47753 17233 47756
rect 17267 47753 17279 47787
rect 17221 47747 17279 47753
rect 17310 47744 17316 47796
rect 17368 47744 17374 47796
rect 17402 47744 17408 47796
rect 17460 47784 17466 47796
rect 18417 47787 18475 47793
rect 18417 47784 18429 47787
rect 17460 47756 18429 47784
rect 17460 47744 17466 47756
rect 18417 47753 18429 47756
rect 18463 47753 18475 47787
rect 18417 47747 18475 47753
rect 18322 47676 18328 47728
rect 18380 47716 18386 47728
rect 18509 47719 18567 47725
rect 18509 47716 18521 47719
rect 18380 47688 18521 47716
rect 18380 47676 18386 47688
rect 18509 47685 18521 47688
rect 18555 47716 18567 47719
rect 18782 47716 18788 47728
rect 18555 47688 18788 47716
rect 18555 47685 18567 47688
rect 18509 47679 18567 47685
rect 18782 47676 18788 47688
rect 18840 47716 18846 47728
rect 19061 47719 19119 47725
rect 19061 47716 19073 47719
rect 18840 47688 19073 47716
rect 18840 47676 18846 47688
rect 19061 47685 19073 47688
rect 19107 47685 19119 47719
rect 19061 47679 19119 47685
rect 9309 47651 9367 47657
rect 9309 47617 9321 47651
rect 9355 47648 9367 47651
rect 11790 47648 11796 47660
rect 9355 47620 11796 47648
rect 9355 47617 9367 47620
rect 9309 47611 9367 47617
rect 11790 47608 11796 47620
rect 11848 47608 11854 47660
rect 24489 47651 24547 47657
rect 24489 47617 24501 47651
rect 24535 47648 24547 47651
rect 25774 47648 25780 47660
rect 24535 47620 25780 47648
rect 24535 47617 24547 47620
rect 24489 47611 24547 47617
rect 25774 47608 25780 47620
rect 25832 47608 25838 47660
rect 17405 47583 17463 47589
rect 17405 47549 17417 47583
rect 17451 47549 17463 47583
rect 17405 47543 17463 47549
rect 16298 47472 16304 47524
rect 16356 47512 16362 47524
rect 17420 47512 17448 47543
rect 18690 47540 18696 47592
rect 18748 47540 18754 47592
rect 23842 47540 23848 47592
rect 23900 47580 23906 47592
rect 24765 47583 24823 47589
rect 24765 47580 24777 47583
rect 23900 47552 24777 47580
rect 23900 47540 23906 47552
rect 24765 47549 24777 47552
rect 24811 47549 24823 47583
rect 24765 47543 24823 47549
rect 16356 47484 17448 47512
rect 16356 47472 16362 47484
rect 16574 47404 16580 47456
rect 16632 47444 16638 47456
rect 16853 47447 16911 47453
rect 16853 47444 16865 47447
rect 16632 47416 16865 47444
rect 16632 47404 16638 47416
rect 16853 47413 16865 47416
rect 16899 47413 16911 47447
rect 16853 47407 16911 47413
rect 17494 47404 17500 47456
rect 17552 47444 17558 47456
rect 18049 47447 18107 47453
rect 18049 47444 18061 47447
rect 17552 47416 18061 47444
rect 17552 47404 17558 47416
rect 18049 47413 18061 47416
rect 18095 47413 18107 47447
rect 18049 47407 18107 47413
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 15920 47243 15978 47249
rect 15920 47209 15932 47243
rect 15966 47240 15978 47243
rect 18690 47240 18696 47252
rect 15966 47212 18696 47240
rect 15966 47209 15978 47212
rect 15920 47203 15978 47209
rect 18690 47200 18696 47212
rect 18748 47200 18754 47252
rect 19334 47200 19340 47252
rect 19392 47200 19398 47252
rect 20438 47200 20444 47252
rect 20496 47240 20502 47252
rect 21637 47243 21695 47249
rect 21637 47240 21649 47243
rect 20496 47212 21649 47240
rect 20496 47200 20502 47212
rect 21637 47209 21649 47212
rect 21683 47240 21695 47243
rect 21683 47212 22416 47240
rect 21683 47209 21695 47212
rect 21637 47203 21695 47209
rect 18141 47175 18199 47181
rect 18141 47141 18153 47175
rect 18187 47172 18199 47175
rect 18506 47172 18512 47184
rect 18187 47144 18512 47172
rect 18187 47141 18199 47144
rect 18141 47135 18199 47141
rect 18506 47132 18512 47144
rect 18564 47132 18570 47184
rect 19352 47172 19380 47200
rect 18708 47144 19380 47172
rect 10226 47064 10232 47116
rect 10284 47064 10290 47116
rect 15657 47107 15715 47113
rect 15657 47073 15669 47107
rect 15703 47104 15715 47107
rect 16666 47104 16672 47116
rect 15703 47076 16672 47104
rect 15703 47073 15715 47076
rect 15657 47067 15715 47073
rect 16666 47064 16672 47076
rect 16724 47064 16730 47116
rect 17218 47064 17224 47116
rect 17276 47104 17282 47116
rect 17405 47107 17463 47113
rect 17405 47104 17417 47107
rect 17276 47076 17417 47104
rect 17276 47064 17282 47076
rect 17405 47073 17417 47076
rect 17451 47073 17463 47107
rect 17405 47067 17463 47073
rect 18598 47064 18604 47116
rect 18656 47064 18662 47116
rect 18509 47039 18567 47045
rect 18509 47005 18521 47039
rect 18555 47036 18567 47039
rect 18708 47036 18736 47144
rect 18785 47107 18843 47113
rect 18785 47073 18797 47107
rect 18831 47104 18843 47107
rect 19334 47104 19340 47116
rect 18831 47076 19340 47104
rect 18831 47073 18843 47076
rect 18785 47067 18843 47073
rect 19334 47064 19340 47076
rect 19392 47064 19398 47116
rect 22388 47045 22416 47212
rect 25133 47175 25191 47181
rect 25133 47141 25145 47175
rect 25179 47172 25191 47175
rect 25590 47172 25596 47184
rect 25179 47144 25596 47172
rect 25179 47141 25191 47144
rect 25133 47135 25191 47141
rect 25590 47132 25596 47144
rect 25648 47132 25654 47184
rect 22462 47064 22468 47116
rect 22520 47064 22526 47116
rect 22554 47064 22560 47116
rect 22612 47064 22618 47116
rect 18555 47008 18736 47036
rect 22373 47039 22431 47045
rect 18555 47005 18567 47008
rect 18509 46999 18567 47005
rect 18616 46980 18644 47008
rect 22373 47005 22385 47039
rect 22419 47005 22431 47039
rect 25317 47039 25375 47045
rect 25317 47036 25329 47039
rect 22373 46999 22431 47005
rect 24872 47008 25329 47036
rect 10505 46971 10563 46977
rect 10505 46937 10517 46971
rect 10551 46968 10563 46971
rect 10778 46968 10784 46980
rect 10551 46940 10784 46968
rect 10551 46937 10563 46940
rect 10505 46931 10563 46937
rect 10778 46928 10784 46940
rect 10836 46928 10842 46980
rect 11730 46940 12388 46968
rect 11977 46903 12035 46909
rect 11977 46869 11989 46903
rect 12023 46900 12035 46903
rect 12158 46900 12164 46912
rect 12023 46872 12164 46900
rect 12023 46869 12035 46872
rect 11977 46863 12035 46869
rect 12158 46860 12164 46872
rect 12216 46860 12222 46912
rect 12360 46909 12388 46940
rect 16390 46928 16396 46980
rect 16448 46928 16454 46980
rect 18598 46928 18604 46980
rect 18656 46928 18662 46980
rect 24762 46928 24768 46980
rect 24820 46968 24826 46980
rect 24872 46977 24900 47008
rect 25317 47005 25329 47008
rect 25363 47005 25375 47039
rect 25317 46999 25375 47005
rect 24857 46971 24915 46977
rect 24857 46968 24869 46971
rect 24820 46940 24869 46968
rect 24820 46928 24826 46940
rect 24857 46937 24869 46940
rect 24903 46937 24915 46971
rect 24857 46931 24915 46937
rect 12345 46903 12403 46909
rect 12345 46869 12357 46903
rect 12391 46900 12403 46903
rect 13906 46900 13912 46912
rect 12391 46872 13912 46900
rect 12391 46869 12403 46872
rect 12345 46863 12403 46869
rect 13906 46860 13912 46872
rect 13964 46900 13970 46912
rect 14185 46903 14243 46909
rect 14185 46900 14197 46903
rect 13964 46872 14197 46900
rect 13964 46860 13970 46872
rect 14185 46869 14197 46872
rect 14231 46869 14243 46903
rect 14185 46863 14243 46869
rect 17586 46860 17592 46912
rect 17644 46900 17650 46912
rect 17681 46903 17739 46909
rect 17681 46900 17693 46903
rect 17644 46872 17693 46900
rect 17644 46860 17650 46872
rect 17681 46869 17693 46872
rect 17727 46869 17739 46903
rect 17681 46863 17739 46869
rect 22002 46860 22008 46912
rect 22060 46860 22066 46912
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 7193 46699 7251 46705
rect 7193 46665 7205 46699
rect 7239 46696 7251 46699
rect 7466 46696 7472 46708
rect 7239 46668 7472 46696
rect 7239 46665 7251 46668
rect 7193 46659 7251 46665
rect 7466 46656 7472 46668
rect 7524 46656 7530 46708
rect 10870 46656 10876 46708
rect 10928 46656 10934 46708
rect 14182 46696 14188 46708
rect 12636 46668 14188 46696
rect 12636 46637 12664 46668
rect 14182 46656 14188 46668
rect 14240 46656 14246 46708
rect 18601 46699 18659 46705
rect 18601 46665 18613 46699
rect 18647 46696 18659 46699
rect 18690 46696 18696 46708
rect 18647 46668 18696 46696
rect 18647 46665 18659 46668
rect 18601 46659 18659 46665
rect 18690 46656 18696 46668
rect 18748 46656 18754 46708
rect 18966 46656 18972 46708
rect 19024 46696 19030 46708
rect 20809 46699 20867 46705
rect 20809 46696 20821 46699
rect 19024 46668 20821 46696
rect 19024 46656 19030 46668
rect 20809 46665 20821 46668
rect 20855 46665 20867 46699
rect 20809 46659 20867 46665
rect 21910 46656 21916 46708
rect 21968 46696 21974 46708
rect 22005 46699 22063 46705
rect 22005 46696 22017 46699
rect 21968 46668 22017 46696
rect 21968 46656 21974 46668
rect 22005 46665 22017 46668
rect 22051 46696 22063 46699
rect 22094 46696 22100 46708
rect 22051 46668 22100 46696
rect 22051 46665 22063 46668
rect 22005 46659 22063 46665
rect 22094 46656 22100 46668
rect 22152 46696 22158 46708
rect 22649 46699 22707 46705
rect 22649 46696 22661 46699
rect 22152 46668 22661 46696
rect 22152 46656 22158 46668
rect 22649 46665 22661 46668
rect 22695 46665 22707 46699
rect 22649 46659 22707 46665
rect 22741 46699 22799 46705
rect 22741 46665 22753 46699
rect 22787 46696 22799 46699
rect 23934 46696 23940 46708
rect 22787 46668 23940 46696
rect 22787 46665 22799 46668
rect 22741 46659 22799 46665
rect 23934 46656 23940 46668
rect 23992 46656 23998 46708
rect 12621 46631 12679 46637
rect 12621 46597 12633 46631
rect 12667 46597 12679 46631
rect 13906 46628 13912 46640
rect 13846 46600 13912 46628
rect 12621 46591 12679 46597
rect 13906 46588 13912 46600
rect 13964 46628 13970 46640
rect 13964 46600 15318 46628
rect 13964 46588 13970 46600
rect 17586 46588 17592 46640
rect 17644 46588 17650 46640
rect 21085 46631 21143 46637
rect 21085 46628 21097 46631
rect 20562 46614 21097 46628
rect 20548 46600 21097 46614
rect 7377 46563 7435 46569
rect 7377 46529 7389 46563
rect 7423 46560 7435 46563
rect 9306 46560 9312 46572
rect 7423 46532 9312 46560
rect 7423 46529 7435 46532
rect 7377 46523 7435 46529
rect 9306 46520 9312 46532
rect 9364 46520 9370 46572
rect 11054 46520 11060 46572
rect 11112 46520 11118 46572
rect 20548 46504 20576 46600
rect 21085 46597 21097 46600
rect 21131 46597 21143 46631
rect 21085 46591 21143 46597
rect 12345 46495 12403 46501
rect 12345 46461 12357 46495
rect 12391 46461 12403 46495
rect 14553 46495 14611 46501
rect 14553 46492 14565 46495
rect 12345 46455 12403 46461
rect 13648 46464 14565 46492
rect 11882 46316 11888 46368
rect 11940 46356 11946 46368
rect 12360 46356 12388 46455
rect 13354 46356 13360 46368
rect 11940 46328 13360 46356
rect 11940 46316 11946 46328
rect 13354 46316 13360 46328
rect 13412 46356 13418 46368
rect 13648 46356 13676 46464
rect 14553 46461 14565 46464
rect 14599 46461 14611 46495
rect 14553 46455 14611 46461
rect 14829 46495 14887 46501
rect 14829 46461 14841 46495
rect 14875 46492 14887 46495
rect 16666 46492 16672 46504
rect 14875 46464 16672 46492
rect 14875 46461 14887 46464
rect 14829 46455 14887 46461
rect 16666 46452 16672 46464
rect 16724 46452 16730 46504
rect 16850 46452 16856 46504
rect 16908 46452 16914 46504
rect 17129 46495 17187 46501
rect 17129 46461 17141 46495
rect 17175 46492 17187 46495
rect 18782 46492 18788 46504
rect 17175 46464 18788 46492
rect 17175 46461 17187 46464
rect 17129 46455 17187 46461
rect 18782 46452 18788 46464
rect 18840 46452 18846 46504
rect 19061 46495 19119 46501
rect 19061 46461 19073 46495
rect 19107 46461 19119 46495
rect 19061 46455 19119 46461
rect 13412 46328 13676 46356
rect 13412 46316 13418 46328
rect 13722 46316 13728 46368
rect 13780 46356 13786 46368
rect 14093 46359 14151 46365
rect 14093 46356 14105 46359
rect 13780 46328 14105 46356
rect 13780 46316 13786 46328
rect 14093 46325 14105 46328
rect 14139 46325 14151 46359
rect 14093 46319 14151 46325
rect 16298 46316 16304 46368
rect 16356 46316 16362 46368
rect 19076 46356 19104 46455
rect 19334 46452 19340 46504
rect 19392 46452 19398 46504
rect 20530 46452 20536 46504
rect 20588 46452 20594 46504
rect 22833 46495 22891 46501
rect 22833 46461 22845 46495
rect 22879 46461 22891 46495
rect 22833 46455 22891 46461
rect 22646 46384 22652 46436
rect 22704 46424 22710 46436
rect 22848 46424 22876 46455
rect 24486 46452 24492 46504
rect 24544 46452 24550 46504
rect 24670 46452 24676 46504
rect 24728 46492 24734 46504
rect 24765 46495 24823 46501
rect 24765 46492 24777 46495
rect 24728 46464 24777 46492
rect 24728 46452 24734 46464
rect 24765 46461 24777 46464
rect 24811 46461 24823 46495
rect 24765 46455 24823 46461
rect 22704 46396 22876 46424
rect 22704 46384 22710 46396
rect 19518 46356 19524 46368
rect 19076 46328 19524 46356
rect 19518 46316 19524 46328
rect 19576 46316 19582 46368
rect 22281 46359 22339 46365
rect 22281 46325 22293 46359
rect 22327 46356 22339 46359
rect 23290 46356 23296 46368
rect 22327 46328 23296 46356
rect 22327 46325 22339 46328
rect 22281 46319 22339 46325
rect 23290 46316 23296 46328
rect 23348 46316 23354 46368
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 5718 46112 5724 46164
rect 5776 46152 5782 46164
rect 8113 46155 8171 46161
rect 8113 46152 8125 46155
rect 5776 46124 8125 46152
rect 5776 46112 5782 46124
rect 8113 46121 8125 46124
rect 8159 46121 8171 46155
rect 8113 46115 8171 46121
rect 9125 46155 9183 46161
rect 9125 46121 9137 46155
rect 9171 46152 9183 46155
rect 9214 46152 9220 46164
rect 9171 46124 9220 46152
rect 9171 46121 9183 46124
rect 9125 46115 9183 46121
rect 9214 46112 9220 46124
rect 9272 46112 9278 46164
rect 10686 46112 10692 46164
rect 10744 46112 10750 46164
rect 24486 46112 24492 46164
rect 24544 46152 24550 46164
rect 24762 46152 24768 46164
rect 24544 46124 24768 46152
rect 24544 46112 24550 46124
rect 24762 46112 24768 46124
rect 24820 46152 24826 46164
rect 25409 46155 25467 46161
rect 25409 46152 25421 46155
rect 24820 46124 25421 46152
rect 24820 46112 24826 46124
rect 25409 46121 25421 46124
rect 25455 46121 25467 46155
rect 25409 46115 25467 46121
rect 7650 46044 7656 46096
rect 7708 46084 7714 46096
rect 10045 46087 10103 46093
rect 10045 46084 10057 46087
rect 7708 46056 10057 46084
rect 7708 46044 7714 46056
rect 10045 46053 10057 46056
rect 10091 46053 10103 46087
rect 10045 46047 10103 46053
rect 11348 46056 12020 46084
rect 1857 46019 1915 46025
rect 1857 45985 1869 46019
rect 1903 46016 1915 46019
rect 9214 46016 9220 46028
rect 1903 45988 9220 46016
rect 1903 45985 1915 45988
rect 1857 45979 1915 45985
rect 9214 45976 9220 45988
rect 9272 45976 9278 46028
rect 11348 46025 11376 46056
rect 11333 46019 11391 46025
rect 11333 45985 11345 46019
rect 11379 45985 11391 46019
rect 11333 45979 11391 45985
rect 11882 45976 11888 46028
rect 11940 45976 11946 46028
rect 11992 46016 12020 46056
rect 12158 46016 12164 46028
rect 11992 45988 12164 46016
rect 12158 45976 12164 45988
rect 12216 45976 12222 46028
rect 20162 45976 20168 46028
rect 20220 45976 20226 46028
rect 20349 46019 20407 46025
rect 20349 45985 20361 46019
rect 20395 46016 20407 46019
rect 20438 46016 20444 46028
rect 20395 45988 20444 46016
rect 20395 45985 20407 45988
rect 20349 45979 20407 45985
rect 20438 45976 20444 45988
rect 20496 45976 20502 46028
rect 21358 45976 21364 46028
rect 21416 45976 21422 46028
rect 21542 45976 21548 46028
rect 21600 45976 21606 46028
rect 1302 45908 1308 45960
rect 1360 45948 1366 45960
rect 1581 45951 1639 45957
rect 1581 45948 1593 45951
rect 1360 45920 1593 45948
rect 1360 45908 1366 45920
rect 1581 45917 1593 45920
rect 1627 45917 1639 45951
rect 1581 45911 1639 45917
rect 8662 45908 8668 45960
rect 8720 45948 8726 45960
rect 9309 45951 9367 45957
rect 9309 45948 9321 45951
rect 8720 45920 9321 45948
rect 8720 45908 8726 45920
rect 9309 45917 9321 45920
rect 9355 45917 9367 45951
rect 9309 45911 9367 45917
rect 10229 45951 10287 45957
rect 10229 45917 10241 45951
rect 10275 45948 10287 45951
rect 10962 45948 10968 45960
rect 10275 45920 10968 45948
rect 10275 45917 10287 45920
rect 10229 45911 10287 45917
rect 10962 45908 10968 45920
rect 11020 45908 11026 45960
rect 20898 45908 20904 45960
rect 20956 45948 20962 45960
rect 21269 45951 21327 45957
rect 21269 45948 21281 45951
rect 20956 45920 21281 45948
rect 20956 45908 20962 45920
rect 21269 45917 21281 45920
rect 21315 45917 21327 45951
rect 21269 45911 21327 45917
rect 23201 45951 23259 45957
rect 23201 45917 23213 45951
rect 23247 45917 23259 45951
rect 23201 45911 23259 45917
rect 7374 45840 7380 45892
rect 7432 45880 7438 45892
rect 8021 45883 8079 45889
rect 8021 45880 8033 45883
rect 7432 45852 8033 45880
rect 7432 45840 7438 45852
rect 8021 45849 8033 45852
rect 8067 45880 8079 45883
rect 8481 45883 8539 45889
rect 8481 45880 8493 45883
rect 8067 45852 8493 45880
rect 8067 45849 8079 45852
rect 8021 45843 8079 45849
rect 8481 45849 8493 45852
rect 8527 45849 8539 45883
rect 8481 45843 8539 45849
rect 11057 45883 11115 45889
rect 11057 45849 11069 45883
rect 11103 45880 11115 45883
rect 11698 45880 11704 45892
rect 11103 45852 11704 45880
rect 11103 45849 11115 45852
rect 11057 45843 11115 45849
rect 11698 45840 11704 45852
rect 11756 45840 11762 45892
rect 13906 45880 13912 45892
rect 13386 45852 13912 45880
rect 13906 45840 13912 45852
rect 13964 45880 13970 45892
rect 19610 45880 19616 45892
rect 13964 45852 14228 45880
rect 13964 45840 13970 45852
rect 11146 45772 11152 45824
rect 11204 45772 11210 45824
rect 13630 45772 13636 45824
rect 13688 45772 13694 45824
rect 14200 45821 14228 45852
rect 19352 45852 19616 45880
rect 14185 45815 14243 45821
rect 14185 45781 14197 45815
rect 14231 45812 14243 45815
rect 15010 45812 15016 45824
rect 14231 45784 15016 45812
rect 14231 45781 14243 45784
rect 14185 45775 14243 45781
rect 15010 45772 15016 45784
rect 15068 45812 15074 45824
rect 16390 45812 16396 45824
rect 15068 45784 16396 45812
rect 15068 45772 15074 45784
rect 16390 45772 16396 45784
rect 16448 45772 16454 45824
rect 17586 45772 17592 45824
rect 17644 45812 17650 45824
rect 18693 45815 18751 45821
rect 18693 45812 18705 45815
rect 17644 45784 18705 45812
rect 17644 45772 17650 45784
rect 18693 45781 18705 45784
rect 18739 45781 18751 45815
rect 18693 45775 18751 45781
rect 19058 45772 19064 45824
rect 19116 45812 19122 45824
rect 19352 45821 19380 45852
rect 19610 45840 19616 45852
rect 19668 45880 19674 45892
rect 20073 45883 20131 45889
rect 20073 45880 20085 45883
rect 19668 45852 20085 45880
rect 19668 45840 19674 45852
rect 20073 45849 20085 45852
rect 20119 45849 20131 45883
rect 20073 45843 20131 45849
rect 19337 45815 19395 45821
rect 19337 45812 19349 45815
rect 19116 45784 19349 45812
rect 19116 45772 19122 45784
rect 19337 45781 19349 45784
rect 19383 45781 19395 45815
rect 19337 45775 19395 45781
rect 19705 45815 19763 45821
rect 19705 45781 19717 45815
rect 19751 45812 19763 45815
rect 19886 45812 19892 45824
rect 19751 45784 19892 45812
rect 19751 45781 19763 45784
rect 19705 45775 19763 45781
rect 19886 45772 19892 45784
rect 19944 45772 19950 45824
rect 20714 45772 20720 45824
rect 20772 45812 20778 45824
rect 20901 45815 20959 45821
rect 20901 45812 20913 45815
rect 20772 45784 20913 45812
rect 20772 45772 20778 45784
rect 20901 45781 20913 45784
rect 20947 45781 20959 45815
rect 23216 45812 23244 45911
rect 23474 45908 23480 45960
rect 23532 45908 23538 45960
rect 24489 45815 24547 45821
rect 24489 45812 24501 45815
rect 23216 45784 24501 45812
rect 20901 45775 20959 45781
rect 24489 45781 24501 45784
rect 24535 45812 24547 45815
rect 24946 45812 24952 45824
rect 24535 45784 24952 45812
rect 24535 45781 24547 45784
rect 24489 45775 24547 45781
rect 24946 45772 24952 45784
rect 25004 45772 25010 45824
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 1302 45568 1308 45620
rect 1360 45608 1366 45620
rect 1397 45611 1455 45617
rect 1397 45608 1409 45611
rect 1360 45580 1409 45608
rect 1360 45568 1366 45580
rect 1397 45577 1409 45580
rect 1443 45577 1455 45611
rect 1397 45571 1455 45577
rect 19334 45568 19340 45620
rect 19392 45608 19398 45620
rect 20165 45611 20223 45617
rect 20165 45608 20177 45611
rect 19392 45580 20177 45608
rect 19392 45568 19398 45580
rect 20165 45577 20177 45580
rect 20211 45577 20223 45611
rect 23753 45611 23811 45617
rect 23753 45608 23765 45611
rect 20165 45571 20223 45577
rect 22664 45580 23765 45608
rect 8754 45500 8760 45552
rect 8812 45540 8818 45552
rect 9490 45540 9496 45552
rect 8812 45512 9496 45540
rect 8812 45500 8818 45512
rect 9490 45500 9496 45512
rect 9548 45500 9554 45552
rect 10870 45540 10876 45552
rect 10718 45512 10876 45540
rect 10870 45500 10876 45512
rect 10928 45500 10934 45552
rect 15930 45540 15936 45552
rect 15870 45512 15936 45540
rect 15930 45500 15936 45512
rect 15988 45540 15994 45552
rect 16393 45543 16451 45549
rect 16393 45540 16405 45543
rect 15988 45512 16405 45540
rect 15988 45500 15994 45512
rect 16393 45509 16405 45512
rect 16439 45509 16451 45543
rect 20530 45540 20536 45552
rect 19918 45512 20536 45540
rect 16393 45503 16451 45509
rect 20530 45500 20536 45512
rect 20588 45500 20594 45552
rect 21542 45500 21548 45552
rect 21600 45540 21606 45552
rect 22664 45540 22692 45580
rect 23753 45577 23765 45580
rect 23799 45577 23811 45611
rect 23753 45571 23811 45577
rect 21600 45512 22692 45540
rect 21600 45500 21606 45512
rect 24026 45472 24032 45484
rect 23414 45444 24032 45472
rect 24026 45432 24032 45444
rect 24084 45432 24090 45484
rect 24394 45432 24400 45484
rect 24452 45472 24458 45484
rect 24765 45475 24823 45481
rect 24765 45472 24777 45475
rect 24452 45444 24777 45472
rect 24452 45432 24458 45444
rect 24765 45441 24777 45444
rect 24811 45441 24823 45475
rect 24765 45435 24823 45441
rect 9217 45407 9275 45413
rect 9217 45373 9229 45407
rect 9263 45373 9275 45407
rect 9217 45367 9275 45373
rect 14369 45407 14427 45413
rect 14369 45373 14381 45407
rect 14415 45404 14427 45407
rect 14645 45407 14703 45413
rect 14415 45376 14504 45404
rect 14415 45373 14427 45376
rect 14369 45367 14427 45373
rect 8754 45228 8760 45280
rect 8812 45268 8818 45280
rect 8849 45271 8907 45277
rect 8849 45268 8861 45271
rect 8812 45240 8861 45268
rect 8812 45228 8818 45240
rect 8849 45237 8861 45240
rect 8895 45237 8907 45271
rect 9232 45268 9260 45367
rect 10778 45296 10784 45348
rect 10836 45336 10842 45348
rect 10965 45339 11023 45345
rect 10965 45336 10977 45339
rect 10836 45308 10977 45336
rect 10836 45296 10842 45308
rect 10965 45305 10977 45308
rect 11011 45336 11023 45339
rect 12250 45336 12256 45348
rect 11011 45308 12256 45336
rect 11011 45305 11023 45308
rect 10965 45299 11023 45305
rect 12250 45296 12256 45308
rect 12308 45296 12314 45348
rect 10226 45268 10232 45280
rect 9232 45240 10232 45268
rect 8849 45231 8907 45237
rect 10226 45228 10232 45240
rect 10284 45228 10290 45280
rect 10870 45228 10876 45280
rect 10928 45268 10934 45280
rect 11241 45271 11299 45277
rect 11241 45268 11253 45271
rect 10928 45240 11253 45268
rect 10928 45228 10934 45240
rect 11241 45237 11253 45240
rect 11287 45237 11299 45271
rect 11241 45231 11299 45237
rect 12161 45271 12219 45277
rect 12161 45237 12173 45271
rect 12207 45268 12219 45271
rect 12434 45268 12440 45280
rect 12207 45240 12440 45268
rect 12207 45237 12219 45240
rect 12161 45231 12219 45237
rect 12434 45228 12440 45240
rect 12492 45228 12498 45280
rect 14476 45268 14504 45376
rect 14645 45373 14657 45407
rect 14691 45404 14703 45407
rect 16298 45404 16304 45416
rect 14691 45376 16304 45404
rect 14691 45373 14703 45376
rect 14645 45367 14703 45373
rect 16298 45364 16304 45376
rect 16356 45364 16362 45416
rect 18322 45364 18328 45416
rect 18380 45404 18386 45416
rect 18417 45407 18475 45413
rect 18417 45404 18429 45407
rect 18380 45376 18429 45404
rect 18380 45364 18386 45376
rect 18417 45373 18429 45376
rect 18463 45373 18475 45407
rect 18417 45367 18475 45373
rect 18693 45407 18751 45413
rect 18693 45373 18705 45407
rect 18739 45404 18751 45407
rect 20070 45404 20076 45416
rect 18739 45376 20076 45404
rect 18739 45373 18751 45376
rect 18693 45367 18751 45373
rect 20070 45364 20076 45376
rect 20128 45364 20134 45416
rect 22005 45407 22063 45413
rect 22005 45373 22017 45407
rect 22051 45373 22063 45407
rect 22005 45367 22063 45373
rect 22281 45407 22339 45413
rect 22281 45373 22293 45407
rect 22327 45404 22339 45407
rect 22738 45404 22744 45416
rect 22327 45376 22744 45404
rect 22327 45373 22339 45376
rect 22281 45367 22339 45373
rect 14826 45268 14832 45280
rect 14476 45240 14832 45268
rect 14826 45228 14832 45240
rect 14884 45228 14890 45280
rect 16114 45228 16120 45280
rect 16172 45228 16178 45280
rect 20530 45228 20536 45280
rect 20588 45228 20594 45280
rect 20806 45228 20812 45280
rect 20864 45228 20870 45280
rect 22020 45268 22048 45367
rect 22738 45364 22744 45376
rect 22796 45364 22802 45416
rect 24486 45364 24492 45416
rect 24544 45364 24550 45416
rect 22278 45268 22284 45280
rect 22020 45240 22284 45268
rect 22278 45228 22284 45240
rect 22336 45228 22342 45280
rect 24026 45228 24032 45280
rect 24084 45228 24090 45280
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 6362 45024 6368 45076
rect 6420 45064 6426 45076
rect 7837 45067 7895 45073
rect 7837 45064 7849 45067
rect 6420 45036 7849 45064
rect 6420 45024 6426 45036
rect 7837 45033 7849 45036
rect 7883 45033 7895 45067
rect 7837 45027 7895 45033
rect 11238 45024 11244 45076
rect 11296 45064 11302 45076
rect 11609 45067 11667 45073
rect 11609 45064 11621 45067
rect 11296 45036 11621 45064
rect 11296 45024 11302 45036
rect 11609 45033 11621 45036
rect 11655 45033 11667 45067
rect 11609 45027 11667 45033
rect 12526 45024 12532 45076
rect 12584 45064 12590 45076
rect 12989 45067 13047 45073
rect 12989 45064 13001 45067
rect 12584 45036 13001 45064
rect 12584 45024 12590 45036
rect 12989 45033 13001 45036
rect 13035 45033 13047 45067
rect 12989 45027 13047 45033
rect 15930 45024 15936 45076
rect 15988 45064 15994 45076
rect 16758 45064 16764 45076
rect 15988 45036 16764 45064
rect 15988 45024 15994 45036
rect 16758 45024 16764 45036
rect 16816 45064 16822 45076
rect 17129 45067 17187 45073
rect 17129 45064 17141 45067
rect 16816 45036 17141 45064
rect 16816 45024 16822 45036
rect 17129 45033 17141 45036
rect 17175 45064 17187 45067
rect 17586 45064 17592 45076
rect 17175 45036 17592 45064
rect 17175 45033 17187 45036
rect 17129 45027 17187 45033
rect 17586 45024 17592 45036
rect 17644 45024 17650 45076
rect 22094 45024 22100 45076
rect 22152 45064 22158 45076
rect 22554 45064 22560 45076
rect 22152 45036 22560 45064
rect 22152 45024 22158 45036
rect 22554 45024 22560 45036
rect 22612 45024 22618 45076
rect 7282 44956 7288 45008
rect 7340 44996 7346 45008
rect 9401 44999 9459 45005
rect 9401 44996 9413 44999
rect 7340 44968 9413 44996
rect 7340 44956 7346 44968
rect 9401 44965 9413 44968
rect 9447 44965 9459 44999
rect 9401 44959 9459 44965
rect 10410 44888 10416 44940
rect 10468 44928 10474 44940
rect 12529 44931 12587 44937
rect 12529 44928 12541 44931
rect 10468 44900 12541 44928
rect 10468 44888 10474 44900
rect 12529 44897 12541 44900
rect 12575 44897 12587 44931
rect 12529 44891 12587 44897
rect 12618 44888 12624 44940
rect 12676 44928 12682 44940
rect 13541 44931 13599 44937
rect 13541 44928 13553 44931
rect 12676 44900 13553 44928
rect 12676 44888 12682 44900
rect 13541 44897 13553 44900
rect 13587 44928 13599 44931
rect 13722 44928 13728 44940
rect 13587 44900 13728 44928
rect 13587 44897 13599 44900
rect 13541 44891 13599 44897
rect 13722 44888 13728 44900
rect 13780 44888 13786 44940
rect 16850 44928 16856 44940
rect 15120 44900 16856 44928
rect 12345 44863 12403 44869
rect 12345 44829 12357 44863
rect 12391 44860 12403 44863
rect 12434 44860 12440 44872
rect 12391 44832 12440 44860
rect 12391 44829 12403 44832
rect 12345 44823 12403 44829
rect 12434 44820 12440 44832
rect 12492 44820 12498 44872
rect 13357 44863 13415 44869
rect 13357 44829 13369 44863
rect 13403 44860 13415 44863
rect 13446 44860 13452 44872
rect 13403 44832 13452 44860
rect 13403 44829 13415 44832
rect 13357 44823 13415 44829
rect 13446 44820 13452 44832
rect 13504 44820 13510 44872
rect 14826 44820 14832 44872
rect 14884 44860 14890 44872
rect 15120 44869 15148 44900
rect 16850 44888 16856 44900
rect 16908 44888 16914 44940
rect 20530 44888 20536 44940
rect 20588 44928 20594 44940
rect 21450 44928 21456 44940
rect 20588 44900 21456 44928
rect 20588 44888 20594 44900
rect 15105 44863 15163 44869
rect 15105 44860 15117 44863
rect 14884 44832 15117 44860
rect 14884 44820 14890 44832
rect 15105 44829 15117 44832
rect 15151 44829 15163 44863
rect 15105 44823 15163 44829
rect 19518 44820 19524 44872
rect 19576 44820 19582 44872
rect 7745 44795 7803 44801
rect 7745 44761 7757 44795
rect 7791 44792 7803 44795
rect 8205 44795 8263 44801
rect 8205 44792 8217 44795
rect 7791 44764 8217 44792
rect 7791 44761 7803 44764
rect 7745 44755 7803 44761
rect 8205 44761 8217 44764
rect 8251 44792 8263 44795
rect 8570 44792 8576 44804
rect 8251 44764 8576 44792
rect 8251 44761 8263 44764
rect 8205 44755 8263 44761
rect 8570 44752 8576 44764
rect 8628 44752 8634 44804
rect 9217 44795 9275 44801
rect 9217 44761 9229 44795
rect 9263 44792 9275 44795
rect 11149 44795 11207 44801
rect 9263 44764 9720 44792
rect 9263 44761 9275 44764
rect 9217 44755 9275 44761
rect 9692 44736 9720 44764
rect 11149 44761 11161 44795
rect 11195 44792 11207 44795
rect 11514 44792 11520 44804
rect 11195 44764 11520 44792
rect 11195 44761 11207 44764
rect 11149 44755 11207 44761
rect 11514 44752 11520 44764
rect 11572 44752 11578 44804
rect 15381 44795 15439 44801
rect 15381 44761 15393 44795
rect 15427 44792 15439 44795
rect 15654 44792 15660 44804
rect 15427 44764 15660 44792
rect 15427 44761 15439 44764
rect 15381 44755 15439 44761
rect 15654 44752 15660 44764
rect 15712 44752 15718 44804
rect 15930 44752 15936 44804
rect 15988 44752 15994 44804
rect 19794 44752 19800 44804
rect 19852 44752 19858 44804
rect 21008 44778 21036 44900
rect 21450 44888 21456 44900
rect 21508 44928 21514 44940
rect 21637 44931 21695 44937
rect 21637 44928 21649 44931
rect 21508 44900 21649 44928
rect 21508 44888 21514 44900
rect 21637 44897 21649 44900
rect 21683 44928 21695 44931
rect 21683 44900 23704 44928
rect 21683 44897 21695 44900
rect 21637 44891 21695 44897
rect 22278 44820 22284 44872
rect 22336 44820 22342 44872
rect 23676 44860 23704 44900
rect 24026 44860 24032 44872
rect 23676 44846 24032 44860
rect 23690 44832 24032 44846
rect 24026 44820 24032 44832
rect 24084 44860 24090 44872
rect 24489 44863 24547 44869
rect 24489 44860 24501 44863
rect 24084 44832 24501 44860
rect 24084 44820 24090 44832
rect 24489 44829 24501 44832
rect 24535 44860 24547 44863
rect 24578 44860 24584 44872
rect 24535 44832 24584 44860
rect 24535 44829 24547 44832
rect 24489 44823 24547 44829
rect 24578 44820 24584 44832
rect 24636 44820 24642 44872
rect 25498 44820 25504 44872
rect 25556 44860 25562 44872
rect 25774 44860 25780 44872
rect 25556 44832 25780 44860
rect 25556 44820 25562 44832
rect 25774 44820 25780 44832
rect 25832 44820 25838 44872
rect 22554 44752 22560 44804
rect 22612 44752 22618 44804
rect 6454 44684 6460 44736
rect 6512 44684 6518 44736
rect 7193 44727 7251 44733
rect 7193 44693 7205 44727
rect 7239 44724 7251 44727
rect 7374 44724 7380 44736
rect 7239 44696 7380 44724
rect 7239 44693 7251 44696
rect 7193 44687 7251 44693
rect 7374 44684 7380 44696
rect 7432 44684 7438 44736
rect 9674 44684 9680 44736
rect 9732 44684 9738 44736
rect 13449 44727 13507 44733
rect 13449 44693 13461 44727
rect 13495 44724 13507 44727
rect 15194 44724 15200 44736
rect 13495 44696 15200 44724
rect 13495 44693 13507 44696
rect 13449 44687 13507 44693
rect 15194 44684 15200 44696
rect 15252 44684 15258 44736
rect 16666 44684 16672 44736
rect 16724 44724 16730 44736
rect 16853 44727 16911 44733
rect 16853 44724 16865 44727
rect 16724 44696 16865 44724
rect 16724 44684 16730 44696
rect 16853 44693 16865 44696
rect 16899 44724 16911 44727
rect 16942 44724 16948 44736
rect 16899 44696 16948 44724
rect 16899 44693 16911 44696
rect 16853 44687 16911 44693
rect 16942 44684 16948 44696
rect 17000 44684 17006 44736
rect 20622 44684 20628 44736
rect 20680 44724 20686 44736
rect 21269 44727 21327 44733
rect 21269 44724 21281 44727
rect 20680 44696 21281 44724
rect 20680 44684 20686 44696
rect 21269 44693 21281 44696
rect 21315 44693 21327 44727
rect 21269 44687 21327 44693
rect 22738 44684 22744 44736
rect 22796 44724 22802 44736
rect 24029 44727 24087 44733
rect 24029 44724 24041 44727
rect 22796 44696 24041 44724
rect 22796 44684 22802 44696
rect 24029 44693 24041 44696
rect 24075 44693 24087 44727
rect 24029 44687 24087 44693
rect 24486 44684 24492 44736
rect 24544 44724 24550 44736
rect 25498 44724 25504 44736
rect 24544 44696 25504 44724
rect 24544 44684 24550 44696
rect 25498 44684 25504 44696
rect 25556 44684 25562 44736
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 5810 44480 5816 44532
rect 5868 44480 5874 44532
rect 6730 44480 6736 44532
rect 6788 44480 6794 44532
rect 7466 44480 7472 44532
rect 7524 44480 7530 44532
rect 7834 44480 7840 44532
rect 7892 44520 7898 44532
rect 8021 44523 8079 44529
rect 8021 44520 8033 44523
rect 7892 44492 8033 44520
rect 7892 44480 7898 44492
rect 8021 44489 8033 44492
rect 8067 44489 8079 44523
rect 8021 44483 8079 44489
rect 9766 44480 9772 44532
rect 9824 44520 9830 44532
rect 11057 44523 11115 44529
rect 11057 44520 11069 44523
rect 9824 44492 11069 44520
rect 9824 44480 9830 44492
rect 11057 44489 11069 44492
rect 11103 44489 11115 44523
rect 11057 44483 11115 44489
rect 11146 44480 11152 44532
rect 11204 44520 11210 44532
rect 11885 44523 11943 44529
rect 11885 44520 11897 44523
rect 11204 44492 11897 44520
rect 11204 44480 11210 44492
rect 11885 44489 11897 44492
rect 11931 44489 11943 44523
rect 11885 44483 11943 44489
rect 12253 44523 12311 44529
rect 12253 44489 12265 44523
rect 12299 44520 12311 44523
rect 15102 44520 15108 44532
rect 12299 44492 15108 44520
rect 12299 44489 12311 44492
rect 12253 44483 12311 44489
rect 15102 44480 15108 44492
rect 15160 44480 15166 44532
rect 18877 44523 18935 44529
rect 18877 44520 18889 44523
rect 17512 44492 18889 44520
rect 7098 44412 7104 44464
rect 7156 44452 7162 44464
rect 9125 44455 9183 44461
rect 9125 44452 9137 44455
rect 7156 44424 9137 44452
rect 7156 44412 7162 44424
rect 9125 44421 9137 44424
rect 9171 44421 9183 44455
rect 9125 44415 9183 44421
rect 10318 44412 10324 44464
rect 10376 44452 10382 44464
rect 11606 44452 11612 44464
rect 10376 44424 11612 44452
rect 10376 44412 10382 44424
rect 11606 44412 11612 44424
rect 11664 44412 11670 44464
rect 12342 44412 12348 44464
rect 12400 44452 12406 44464
rect 13354 44452 13360 44464
rect 12400 44424 13360 44452
rect 12400 44412 12406 44424
rect 5350 44344 5356 44396
rect 5408 44384 5414 44396
rect 5997 44387 6055 44393
rect 5997 44384 6009 44387
rect 5408 44356 6009 44384
rect 5408 44344 5414 44356
rect 5997 44353 6009 44356
rect 6043 44353 6055 44387
rect 5997 44347 6055 44353
rect 6454 44344 6460 44396
rect 6512 44384 6518 44396
rect 6641 44387 6699 44393
rect 6641 44384 6653 44387
rect 6512 44356 6653 44384
rect 6512 44344 6518 44356
rect 6641 44353 6653 44356
rect 6687 44353 6699 44387
rect 6641 44347 6699 44353
rect 7374 44344 7380 44396
rect 7432 44344 7438 44396
rect 7466 44344 7472 44396
rect 7524 44384 7530 44396
rect 8205 44387 8263 44393
rect 8205 44384 8217 44387
rect 7524 44356 8217 44384
rect 7524 44344 7530 44356
rect 8205 44353 8217 44356
rect 8251 44353 8263 44387
rect 8205 44347 8263 44353
rect 8941 44387 8999 44393
rect 8941 44353 8953 44387
rect 8987 44384 8999 44387
rect 9398 44384 9404 44396
rect 8987 44356 9404 44384
rect 8987 44353 8999 44356
rect 8941 44347 8999 44353
rect 9398 44344 9404 44356
rect 9456 44344 9462 44396
rect 10965 44387 11023 44393
rect 10965 44353 10977 44387
rect 11011 44384 11023 44387
rect 11514 44384 11520 44396
rect 11011 44356 11520 44384
rect 11011 44353 11023 44356
rect 10965 44347 11023 44353
rect 11514 44344 11520 44356
rect 11572 44344 11578 44396
rect 13188 44393 13216 44424
rect 13354 44412 13360 44424
rect 13412 44412 13418 44464
rect 15010 44452 15016 44464
rect 14674 44424 15016 44452
rect 15010 44412 15016 44424
rect 15068 44412 15074 44464
rect 17512 44452 17540 44492
rect 18877 44489 18889 44492
rect 18923 44520 18935 44523
rect 18923 44492 19334 44520
rect 18923 44489 18935 44492
rect 18877 44483 18935 44489
rect 17586 44452 17592 44464
rect 17512 44424 17592 44452
rect 17586 44412 17592 44424
rect 17644 44412 17650 44464
rect 19306 44452 19334 44492
rect 19794 44480 19800 44532
rect 19852 44520 19858 44532
rect 20438 44520 20444 44532
rect 19852 44492 20444 44520
rect 19852 44480 19858 44492
rect 20438 44480 20444 44492
rect 20496 44520 20502 44532
rect 21269 44523 21327 44529
rect 21269 44520 21281 44523
rect 20496 44492 21281 44520
rect 20496 44480 20502 44492
rect 21269 44489 21281 44492
rect 21315 44489 21327 44523
rect 21269 44483 21327 44489
rect 21450 44480 21456 44532
rect 21508 44520 21514 44532
rect 21545 44523 21603 44529
rect 21545 44520 21557 44523
rect 21508 44492 21557 44520
rect 21508 44480 21514 44492
rect 21545 44489 21557 44492
rect 21591 44489 21603 44523
rect 21545 44483 21603 44489
rect 22554 44480 22560 44532
rect 22612 44520 22618 44532
rect 24029 44523 24087 44529
rect 24029 44520 24041 44523
rect 22612 44492 24041 44520
rect 22612 44480 22618 44492
rect 24029 44489 24041 44492
rect 24075 44489 24087 44523
rect 24029 44483 24087 44489
rect 20254 44452 20260 44464
rect 19306 44424 20260 44452
rect 20254 44412 20260 44424
rect 20312 44412 20318 44464
rect 20530 44412 20536 44464
rect 20588 44412 20594 44464
rect 22094 44412 22100 44464
rect 22152 44452 22158 44464
rect 22646 44452 22652 44464
rect 22152 44424 22652 44452
rect 22152 44412 22158 44424
rect 22646 44412 22652 44424
rect 22704 44412 22710 44464
rect 24578 44452 24584 44464
rect 23782 44424 24584 44452
rect 24578 44412 24584 44424
rect 24636 44412 24642 44464
rect 13173 44387 13231 44393
rect 13173 44353 13185 44387
rect 13219 44353 13231 44387
rect 13173 44347 13231 44353
rect 24489 44387 24547 44393
rect 24489 44353 24501 44387
rect 24535 44384 24547 44387
rect 25314 44384 25320 44396
rect 24535 44356 25320 44384
rect 24535 44353 24547 44356
rect 24489 44347 24547 44353
rect 25314 44344 25320 44356
rect 25372 44344 25378 44396
rect 7392 44316 7420 44344
rect 10594 44316 10600 44328
rect 7392 44288 10600 44316
rect 10594 44276 10600 44288
rect 10652 44276 10658 44328
rect 11146 44276 11152 44328
rect 11204 44316 11210 44328
rect 12345 44319 12403 44325
rect 12345 44316 12357 44319
rect 11204 44288 12357 44316
rect 11204 44276 11210 44288
rect 12345 44285 12357 44288
rect 12391 44285 12403 44319
rect 12345 44279 12403 44285
rect 12437 44319 12495 44325
rect 12437 44285 12449 44319
rect 12483 44285 12495 44319
rect 12437 44279 12495 44285
rect 12250 44208 12256 44260
rect 12308 44248 12314 44260
rect 12452 44248 12480 44279
rect 14182 44276 14188 44328
rect 14240 44316 14246 44328
rect 14921 44319 14979 44325
rect 14921 44316 14933 44319
rect 14240 44288 14933 44316
rect 14240 44276 14246 44288
rect 14921 44285 14933 44288
rect 14967 44285 14979 44319
rect 14921 44279 14979 44285
rect 16850 44276 16856 44328
rect 16908 44276 16914 44328
rect 17129 44319 17187 44325
rect 17129 44285 17141 44319
rect 17175 44316 17187 44319
rect 18966 44316 18972 44328
rect 17175 44288 18972 44316
rect 17175 44285 17187 44288
rect 17129 44279 17187 44285
rect 18966 44276 18972 44288
rect 19024 44276 19030 44328
rect 19518 44276 19524 44328
rect 19576 44276 19582 44328
rect 19797 44319 19855 44325
rect 19797 44285 19809 44319
rect 19843 44316 19855 44319
rect 21174 44316 21180 44328
rect 19843 44288 21180 44316
rect 19843 44285 19855 44288
rect 19797 44279 19855 44285
rect 21174 44276 21180 44288
rect 21232 44276 21238 44328
rect 22278 44276 22284 44328
rect 22336 44276 22342 44328
rect 22557 44319 22615 44325
rect 22557 44285 22569 44319
rect 22603 44316 22615 44319
rect 22646 44316 22652 44328
rect 22603 44288 22652 44316
rect 22603 44285 22615 44288
rect 22557 44279 22615 44285
rect 22646 44276 22652 44288
rect 22704 44276 22710 44328
rect 23934 44276 23940 44328
rect 23992 44316 23998 44328
rect 24765 44319 24823 44325
rect 24765 44316 24777 44319
rect 23992 44288 24777 44316
rect 23992 44276 23998 44288
rect 24765 44285 24777 44288
rect 24811 44285 24823 44319
rect 24765 44279 24823 44285
rect 12308 44220 12480 44248
rect 12308 44208 12314 44220
rect 11514 44140 11520 44192
rect 11572 44140 11578 44192
rect 13436 44183 13494 44189
rect 13436 44149 13448 44183
rect 13482 44180 13494 44183
rect 13630 44180 13636 44192
rect 13482 44152 13636 44180
rect 13482 44149 13494 44152
rect 13436 44143 13494 44149
rect 13630 44140 13636 44152
rect 13688 44140 13694 44192
rect 15010 44140 15016 44192
rect 15068 44180 15074 44192
rect 15197 44183 15255 44189
rect 15197 44180 15209 44183
rect 15068 44152 15209 44180
rect 15068 44140 15074 44152
rect 15197 44149 15209 44152
rect 15243 44149 15255 44183
rect 16868 44180 16896 44276
rect 18322 44180 18328 44192
rect 16868 44152 18328 44180
rect 15197 44143 15255 44149
rect 18322 44140 18328 44152
rect 18380 44140 18386 44192
rect 18601 44183 18659 44189
rect 18601 44149 18613 44183
rect 18647 44180 18659 44183
rect 18782 44180 18788 44192
rect 18647 44152 18788 44180
rect 18647 44149 18659 44152
rect 18601 44143 18659 44149
rect 18782 44140 18788 44152
rect 18840 44140 18846 44192
rect 19536 44180 19564 44276
rect 22278 44180 22284 44192
rect 19536 44152 22284 44180
rect 22278 44140 22284 44152
rect 22336 44140 22342 44192
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 4706 43936 4712 43988
rect 4764 43976 4770 43988
rect 6825 43979 6883 43985
rect 6825 43976 6837 43979
rect 4764 43948 6837 43976
rect 4764 43936 4770 43948
rect 6825 43945 6837 43948
rect 6871 43945 6883 43979
rect 6825 43939 6883 43945
rect 8386 43936 8392 43988
rect 8444 43936 8450 43988
rect 11606 43936 11612 43988
rect 11664 43936 11670 43988
rect 9401 43843 9459 43849
rect 9401 43809 9413 43843
rect 9447 43840 9459 43843
rect 16022 43840 16028 43852
rect 9447 43812 16028 43840
rect 9447 43809 9459 43812
rect 9401 43803 9459 43809
rect 16022 43800 16028 43812
rect 16080 43800 16086 43852
rect 22186 43800 22192 43852
rect 22244 43840 22250 43852
rect 22465 43843 22523 43849
rect 22465 43840 22477 43843
rect 22244 43812 22477 43840
rect 22244 43800 22250 43812
rect 22465 43809 22477 43812
rect 22511 43809 22523 43843
rect 22465 43803 22523 43809
rect 22649 43843 22707 43849
rect 22649 43809 22661 43843
rect 22695 43840 22707 43843
rect 23382 43840 23388 43852
rect 22695 43812 23388 43840
rect 22695 43809 22707 43812
rect 22649 43803 22707 43809
rect 23382 43800 23388 43812
rect 23440 43800 23446 43852
rect 8573 43775 8631 43781
rect 8573 43741 8585 43775
rect 8619 43772 8631 43775
rect 9030 43772 9036 43784
rect 8619 43744 9036 43772
rect 8619 43741 8631 43744
rect 8573 43735 8631 43741
rect 9030 43732 9036 43744
rect 9088 43732 9094 43784
rect 9122 43732 9128 43784
rect 9180 43732 9186 43784
rect 6733 43707 6791 43713
rect 6733 43673 6745 43707
rect 6779 43704 6791 43707
rect 7193 43707 7251 43713
rect 7193 43704 7205 43707
rect 6779 43676 7205 43704
rect 6779 43673 6791 43676
rect 6733 43667 6791 43673
rect 7193 43673 7205 43676
rect 7239 43673 7251 43707
rect 10778 43704 10784 43716
rect 10626 43676 10784 43704
rect 7193 43667 7251 43673
rect 7208 43636 7236 43667
rect 10778 43664 10784 43676
rect 10836 43664 10842 43716
rect 11517 43707 11575 43713
rect 11517 43673 11529 43707
rect 11563 43704 11575 43707
rect 11882 43704 11888 43716
rect 11563 43676 11888 43704
rect 11563 43673 11575 43676
rect 11517 43667 11575 43673
rect 11882 43664 11888 43676
rect 11940 43704 11946 43716
rect 11977 43707 12035 43713
rect 11977 43704 11989 43707
rect 11940 43676 11989 43704
rect 11940 43664 11946 43676
rect 11977 43673 11989 43676
rect 12023 43673 12035 43707
rect 11977 43667 12035 43673
rect 17402 43664 17408 43716
rect 17460 43704 17466 43716
rect 18598 43704 18604 43716
rect 17460 43676 18604 43704
rect 17460 43664 17466 43676
rect 18598 43664 18604 43676
rect 18656 43664 18662 43716
rect 21726 43704 21732 43716
rect 21652 43676 21732 43704
rect 10318 43636 10324 43648
rect 7208 43608 10324 43636
rect 10318 43596 10324 43608
rect 10376 43596 10382 43648
rect 10686 43596 10692 43648
rect 10744 43636 10750 43648
rect 10873 43639 10931 43645
rect 10873 43636 10885 43639
rect 10744 43608 10885 43636
rect 10744 43596 10750 43608
rect 10873 43605 10885 43608
rect 10919 43636 10931 43639
rect 11238 43636 11244 43648
rect 10919 43608 11244 43636
rect 10919 43605 10931 43608
rect 10873 43599 10931 43605
rect 11238 43596 11244 43608
rect 11296 43596 11302 43648
rect 17586 43596 17592 43648
rect 17644 43636 17650 43648
rect 17957 43639 18015 43645
rect 17957 43636 17969 43639
rect 17644 43608 17969 43636
rect 17644 43596 17650 43608
rect 17957 43605 17969 43608
rect 18003 43636 18015 43639
rect 19518 43636 19524 43648
rect 18003 43608 19524 43636
rect 18003 43605 18015 43608
rect 17957 43599 18015 43605
rect 19518 43596 19524 43608
rect 19576 43596 19582 43648
rect 20806 43596 20812 43648
rect 20864 43636 20870 43648
rect 21652 43645 21680 43676
rect 21726 43664 21732 43676
rect 21784 43704 21790 43716
rect 22373 43707 22431 43713
rect 22373 43704 22385 43707
rect 21784 43676 22385 43704
rect 21784 43664 21790 43676
rect 22373 43673 22385 43676
rect 22419 43673 22431 43707
rect 25409 43707 25467 43713
rect 25409 43704 25421 43707
rect 22373 43667 22431 43673
rect 24596 43676 25421 43704
rect 24596 43648 24624 43676
rect 25409 43673 25421 43676
rect 25455 43673 25467 43707
rect 25409 43667 25467 43673
rect 21637 43639 21695 43645
rect 21637 43636 21649 43639
rect 20864 43608 21649 43636
rect 20864 43596 20870 43608
rect 21637 43605 21649 43608
rect 21683 43605 21695 43639
rect 21637 43599 21695 43605
rect 21910 43596 21916 43648
rect 21968 43636 21974 43648
rect 22005 43639 22063 43645
rect 22005 43636 22017 43639
rect 21968 43608 22017 43636
rect 21968 43596 21974 43608
rect 22005 43605 22017 43608
rect 22051 43605 22063 43639
rect 22005 43599 22063 43605
rect 24213 43639 24271 43645
rect 24213 43605 24225 43639
rect 24259 43636 24271 43639
rect 24578 43636 24584 43648
rect 24259 43608 24584 43636
rect 24259 43605 24271 43608
rect 24213 43599 24271 43605
rect 24578 43596 24584 43608
rect 24636 43596 24642 43648
rect 25314 43596 25320 43648
rect 25372 43636 25378 43648
rect 25498 43636 25504 43648
rect 25372 43608 25504 43636
rect 25372 43596 25378 43608
rect 25498 43596 25504 43608
rect 25556 43596 25562 43648
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 7742 43392 7748 43444
rect 7800 43392 7806 43444
rect 8938 43392 8944 43444
rect 8996 43432 9002 43444
rect 9490 43432 9496 43444
rect 8996 43404 9496 43432
rect 8996 43392 9002 43404
rect 9490 43392 9496 43404
rect 9548 43392 9554 43444
rect 10134 43392 10140 43444
rect 10192 43432 10198 43444
rect 10597 43435 10655 43441
rect 10597 43432 10609 43435
rect 10192 43404 10609 43432
rect 10192 43392 10198 43404
rect 10597 43401 10609 43404
rect 10643 43401 10655 43435
rect 10597 43395 10655 43401
rect 14093 43435 14151 43441
rect 14093 43401 14105 43435
rect 14139 43401 14151 43435
rect 14093 43395 14151 43401
rect 4614 43324 4620 43376
rect 4672 43364 4678 43376
rect 8665 43367 8723 43373
rect 8665 43364 8677 43367
rect 4672 43336 8677 43364
rect 4672 43324 4678 43336
rect 8665 43333 8677 43336
rect 8711 43333 8723 43367
rect 8665 43327 8723 43333
rect 12618 43324 12624 43376
rect 12676 43324 12682 43376
rect 14108 43364 14136 43395
rect 14458 43392 14464 43444
rect 14516 43432 14522 43444
rect 15013 43435 15071 43441
rect 15013 43432 15025 43435
rect 14516 43404 15025 43432
rect 14516 43392 14522 43404
rect 15013 43401 15025 43404
rect 15059 43401 15071 43435
rect 15013 43395 15071 43401
rect 16758 43392 16764 43444
rect 16816 43392 16822 43444
rect 17494 43392 17500 43444
rect 17552 43392 17558 43444
rect 20070 43392 20076 43444
rect 20128 43392 20134 43444
rect 22370 43392 22376 43444
rect 22428 43432 22434 43444
rect 22465 43435 22523 43441
rect 22465 43432 22477 43435
rect 22428 43404 22477 43432
rect 22428 43392 22434 43404
rect 22465 43401 22477 43404
rect 22511 43401 22523 43435
rect 22465 43395 22523 43401
rect 15470 43364 15476 43376
rect 14108 43336 15476 43364
rect 15470 43324 15476 43336
rect 15528 43324 15534 43376
rect 17405 43367 17463 43373
rect 17405 43333 17417 43367
rect 17451 43364 17463 43367
rect 17586 43364 17592 43376
rect 17451 43336 17592 43364
rect 17451 43333 17463 43336
rect 17405 43327 17463 43333
rect 17586 43324 17592 43336
rect 17644 43324 17650 43376
rect 20530 43364 20536 43376
rect 19826 43336 20536 43364
rect 20530 43324 20536 43336
rect 20588 43324 20594 43376
rect 23566 43324 23572 43376
rect 23624 43364 23630 43376
rect 23845 43367 23903 43373
rect 23845 43364 23857 43367
rect 23624 43336 23857 43364
rect 23624 43324 23630 43336
rect 23845 43333 23857 43336
rect 23891 43333 23903 43367
rect 23845 43327 23903 43333
rect 24578 43324 24584 43376
rect 24636 43324 24642 43376
rect 1302 43256 1308 43308
rect 1360 43296 1366 43308
rect 1673 43299 1731 43305
rect 1673 43296 1685 43299
rect 1360 43268 1685 43296
rect 1360 43256 1366 43268
rect 1673 43265 1685 43268
rect 1719 43296 1731 43299
rect 2133 43299 2191 43305
rect 2133 43296 2145 43299
rect 1719 43268 2145 43296
rect 1719 43265 1731 43268
rect 1673 43259 1731 43265
rect 2133 43265 2145 43268
rect 2179 43265 2191 43299
rect 2133 43259 2191 43265
rect 6914 43256 6920 43308
rect 6972 43296 6978 43308
rect 7929 43299 7987 43305
rect 7929 43296 7941 43299
rect 6972 43268 7941 43296
rect 6972 43256 6978 43268
rect 7929 43265 7941 43268
rect 7975 43265 7987 43299
rect 7929 43259 7987 43265
rect 8478 43256 8484 43308
rect 8536 43256 8542 43308
rect 8754 43256 8760 43308
rect 8812 43296 8818 43308
rect 8938 43296 8944 43308
rect 8812 43268 8944 43296
rect 8812 43256 8818 43268
rect 8938 43256 8944 43268
rect 8996 43296 9002 43308
rect 8996 43268 9720 43296
rect 8996 43256 9002 43268
rect 9214 43188 9220 43240
rect 9272 43228 9278 43240
rect 9582 43228 9588 43240
rect 9272 43200 9588 43228
rect 9272 43188 9278 43200
rect 9582 43188 9588 43200
rect 9640 43188 9646 43240
rect 9692 43237 9720 43268
rect 10410 43256 10416 43308
rect 10468 43296 10474 43308
rect 10505 43299 10563 43305
rect 10505 43296 10517 43299
rect 10468 43268 10517 43296
rect 10468 43256 10474 43268
rect 10505 43265 10517 43268
rect 10551 43265 10563 43299
rect 10505 43259 10563 43265
rect 12342 43256 12348 43308
rect 12400 43256 12406 43308
rect 13722 43256 13728 43308
rect 13780 43256 13786 43308
rect 15105 43299 15163 43305
rect 15105 43265 15117 43299
rect 15151 43296 15163 43299
rect 15378 43296 15384 43308
rect 15151 43268 15384 43296
rect 15151 43265 15163 43268
rect 15105 43259 15163 43265
rect 15378 43256 15384 43268
rect 15436 43256 15442 43308
rect 21634 43256 21640 43308
rect 21692 43296 21698 43308
rect 22373 43299 22431 43305
rect 22373 43296 22385 43299
rect 21692 43268 22385 43296
rect 21692 43256 21698 43268
rect 22373 43265 22385 43268
rect 22419 43265 22431 43299
rect 22373 43259 22431 43265
rect 9677 43231 9735 43237
rect 9677 43197 9689 43231
rect 9723 43197 9735 43231
rect 9677 43191 9735 43197
rect 15197 43231 15255 43237
rect 15197 43197 15209 43231
rect 15243 43197 15255 43231
rect 15197 43191 15255 43197
rect 1857 43163 1915 43169
rect 1857 43129 1869 43163
rect 1903 43160 1915 43163
rect 3970 43160 3976 43172
rect 1903 43132 3976 43160
rect 1903 43129 1915 43132
rect 1857 43123 1915 43129
rect 3970 43120 3976 43132
rect 4028 43120 4034 43172
rect 9125 43163 9183 43169
rect 9125 43129 9137 43163
rect 9171 43160 9183 43163
rect 11146 43160 11152 43172
rect 9171 43132 11152 43160
rect 9171 43129 9183 43132
rect 9125 43123 9183 43129
rect 11146 43120 11152 43132
rect 11204 43120 11210 43172
rect 14734 43120 14740 43172
rect 14792 43160 14798 43172
rect 15212 43160 15240 43191
rect 15654 43188 15660 43240
rect 15712 43228 15718 43240
rect 17218 43228 17224 43240
rect 15712 43200 17224 43228
rect 15712 43188 15718 43200
rect 17218 43188 17224 43200
rect 17276 43228 17282 43240
rect 17589 43231 17647 43237
rect 17589 43228 17601 43231
rect 17276 43200 17601 43228
rect 17276 43188 17282 43200
rect 17589 43197 17601 43200
rect 17635 43197 17647 43231
rect 17589 43191 17647 43197
rect 18322 43188 18328 43240
rect 18380 43188 18386 43240
rect 18601 43231 18659 43237
rect 18601 43197 18613 43231
rect 18647 43228 18659 43231
rect 20622 43228 20628 43240
rect 18647 43200 20628 43228
rect 18647 43197 18659 43200
rect 18601 43191 18659 43197
rect 14792 43132 15240 43160
rect 14792 43120 14798 43132
rect 10778 43052 10784 43104
rect 10836 43092 10842 43104
rect 11057 43095 11115 43101
rect 11057 43092 11069 43095
rect 10836 43064 11069 43092
rect 10836 43052 10842 43064
rect 11057 43061 11069 43064
rect 11103 43092 11115 43095
rect 12158 43092 12164 43104
rect 11103 43064 12164 43092
rect 11103 43061 11115 43064
rect 11057 43055 11115 43061
rect 12158 43052 12164 43064
rect 12216 43052 12222 43104
rect 14642 43052 14648 43104
rect 14700 43052 14706 43104
rect 15378 43052 15384 43104
rect 15436 43092 15442 43104
rect 15657 43095 15715 43101
rect 15657 43092 15669 43095
rect 15436 43064 15669 43092
rect 15436 43052 15442 43064
rect 15657 43061 15669 43064
rect 15703 43061 15715 43095
rect 15657 43055 15715 43061
rect 17034 43052 17040 43104
rect 17092 43052 17098 43104
rect 18340 43092 18368 43188
rect 19720 43172 19748 43200
rect 20622 43188 20628 43200
rect 20680 43188 20686 43240
rect 22646 43188 22652 43240
rect 22704 43188 22710 43240
rect 23474 43188 23480 43240
rect 23532 43228 23538 43240
rect 23569 43231 23627 43237
rect 23569 43228 23581 43231
rect 23532 43200 23581 43228
rect 23532 43188 23538 43200
rect 23569 43197 23581 43200
rect 23615 43197 23627 43231
rect 23569 43191 23627 43197
rect 19702 43120 19708 43172
rect 19760 43120 19766 43172
rect 19242 43092 19248 43104
rect 18340 43064 19248 43092
rect 19242 43052 19248 43064
rect 19300 43052 19306 43104
rect 20441 43095 20499 43101
rect 20441 43061 20453 43095
rect 20487 43092 20499 43095
rect 20530 43092 20536 43104
rect 20487 43064 20536 43092
rect 20487 43061 20499 43064
rect 20441 43055 20499 43061
rect 20530 43052 20536 43064
rect 20588 43092 20594 43104
rect 20898 43092 20904 43104
rect 20588 43064 20904 43092
rect 20588 43052 20594 43064
rect 20898 43052 20904 43064
rect 20956 43092 20962 43104
rect 21361 43095 21419 43101
rect 21361 43092 21373 43095
rect 20956 43064 21373 43092
rect 20956 43052 20962 43064
rect 21361 43061 21373 43064
rect 21407 43061 21419 43095
rect 21361 43055 21419 43061
rect 21634 43052 21640 43104
rect 21692 43052 21698 43104
rect 22005 43095 22063 43101
rect 22005 43061 22017 43095
rect 22051 43092 22063 43095
rect 24946 43092 24952 43104
rect 22051 43064 24952 43092
rect 22051 43061 22063 43064
rect 22005 43055 22063 43061
rect 24946 43052 24952 43064
rect 25004 43052 25010 43104
rect 25317 43095 25375 43101
rect 25317 43061 25329 43095
rect 25363 43092 25375 43095
rect 25498 43092 25504 43104
rect 25363 43064 25504 43092
rect 25363 43061 25375 43064
rect 25317 43055 25375 43061
rect 25498 43052 25504 43064
rect 25556 43052 25562 43104
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 8297 42891 8355 42897
rect 8297 42857 8309 42891
rect 8343 42888 8355 42891
rect 8478 42888 8484 42900
rect 8343 42860 8484 42888
rect 8343 42857 8355 42860
rect 8297 42851 8355 42857
rect 8478 42848 8484 42860
rect 8536 42848 8542 42900
rect 8938 42848 8944 42900
rect 8996 42888 9002 42900
rect 19784 42891 19842 42897
rect 8996 42860 17724 42888
rect 8996 42848 9002 42860
rect 12434 42780 12440 42832
rect 12492 42820 12498 42832
rect 14550 42820 14556 42832
rect 12492 42792 14556 42820
rect 12492 42780 12498 42792
rect 14550 42780 14556 42792
rect 14608 42780 14614 42832
rect 17129 42823 17187 42829
rect 17129 42789 17141 42823
rect 17175 42789 17187 42823
rect 17129 42783 17187 42789
rect 4890 42712 4896 42764
rect 4948 42752 4954 42764
rect 4985 42755 5043 42761
rect 4985 42752 4997 42755
rect 4948 42724 4997 42752
rect 4948 42712 4954 42724
rect 4985 42721 4997 42724
rect 5031 42721 5043 42755
rect 4985 42715 5043 42721
rect 9122 42712 9128 42764
rect 9180 42752 9186 42764
rect 10781 42755 10839 42761
rect 10781 42752 10793 42755
rect 9180 42724 10793 42752
rect 9180 42712 9186 42724
rect 10781 42721 10793 42724
rect 10827 42752 10839 42755
rect 12342 42752 12348 42764
rect 10827 42724 12348 42752
rect 10827 42721 10839 42724
rect 10781 42715 10839 42721
rect 12342 42712 12348 42724
rect 12400 42712 12406 42764
rect 14826 42712 14832 42764
rect 14884 42712 14890 42764
rect 15102 42712 15108 42764
rect 15160 42752 15166 42764
rect 17144 42752 17172 42783
rect 17696 42761 17724 42860
rect 19784 42857 19796 42891
rect 19830 42888 19842 42891
rect 20346 42888 20352 42900
rect 19830 42860 20352 42888
rect 19830 42857 19842 42860
rect 19784 42851 19842 42857
rect 20346 42848 20352 42860
rect 20404 42888 20410 42900
rect 21542 42888 21548 42900
rect 20404 42860 21548 42888
rect 20404 42848 20410 42860
rect 21542 42848 21548 42860
rect 21600 42848 21606 42900
rect 15160 42724 17172 42752
rect 17681 42755 17739 42761
rect 15160 42712 15166 42724
rect 17681 42721 17693 42755
rect 17727 42752 17739 42755
rect 18141 42755 18199 42761
rect 18141 42752 18153 42755
rect 17727 42724 18153 42752
rect 17727 42721 17739 42724
rect 17681 42715 17739 42721
rect 18141 42721 18153 42724
rect 18187 42721 18199 42755
rect 18141 42715 18199 42721
rect 19521 42755 19579 42761
rect 19521 42721 19533 42755
rect 19567 42752 19579 42755
rect 19567 42724 21772 42752
rect 19567 42721 19579 42724
rect 19521 42715 19579 42721
rect 12158 42644 12164 42696
rect 12216 42684 12222 42696
rect 12618 42684 12624 42696
rect 12216 42656 12624 42684
rect 12216 42644 12222 42656
rect 12618 42644 12624 42656
rect 12676 42644 12682 42696
rect 21744 42684 21772 42724
rect 22002 42712 22008 42764
rect 22060 42752 22066 42764
rect 22281 42755 22339 42761
rect 22281 42752 22293 42755
rect 22060 42724 22293 42752
rect 22060 42712 22066 42724
rect 22281 42721 22293 42724
rect 22327 42721 22339 42755
rect 22281 42715 22339 42721
rect 22465 42755 22523 42761
rect 22465 42721 22477 42755
rect 22511 42752 22523 42755
rect 22554 42752 22560 42764
rect 22511 42724 22560 42752
rect 22511 42721 22523 42724
rect 22465 42715 22523 42721
rect 22554 42712 22560 42724
rect 22612 42712 22618 42764
rect 25130 42752 25136 42764
rect 22940 42724 25136 42752
rect 22186 42684 22192 42696
rect 21744 42656 22192 42684
rect 22186 42644 22192 42656
rect 22244 42644 22250 42696
rect 4801 42619 4859 42625
rect 4801 42585 4813 42619
rect 4847 42616 4859 42619
rect 4847 42588 5304 42616
rect 4847 42585 4859 42588
rect 4801 42579 4859 42585
rect 5276 42560 5304 42588
rect 8846 42576 8852 42628
rect 8904 42616 8910 42628
rect 9309 42619 9367 42625
rect 9309 42616 9321 42619
rect 8904 42588 9321 42616
rect 8904 42576 8910 42588
rect 9309 42585 9321 42588
rect 9355 42585 9367 42619
rect 11057 42619 11115 42625
rect 11057 42616 11069 42619
rect 9309 42579 9367 42585
rect 10888 42588 11069 42616
rect 10888 42560 10916 42588
rect 11057 42585 11069 42588
rect 11103 42585 11115 42619
rect 15105 42619 15163 42625
rect 15105 42616 15117 42619
rect 11057 42579 11115 42585
rect 12544 42588 15117 42616
rect 5258 42508 5264 42560
rect 5316 42508 5322 42560
rect 8294 42508 8300 42560
rect 8352 42548 8358 42560
rect 8754 42548 8760 42560
rect 8352 42520 8760 42548
rect 8352 42508 8358 42520
rect 8754 42508 8760 42520
rect 8812 42508 8818 42560
rect 8938 42508 8944 42560
rect 8996 42508 9002 42560
rect 10321 42551 10379 42557
rect 10321 42517 10333 42551
rect 10367 42548 10379 42551
rect 10410 42548 10416 42560
rect 10367 42520 10416 42548
rect 10367 42517 10379 42520
rect 10321 42511 10379 42517
rect 10410 42508 10416 42520
rect 10468 42508 10474 42560
rect 10870 42508 10876 42560
rect 10928 42508 10934 42560
rect 12434 42508 12440 42560
rect 12492 42548 12498 42560
rect 12544 42557 12572 42588
rect 15105 42585 15117 42588
rect 15151 42585 15163 42619
rect 17497 42619 17555 42625
rect 15105 42579 15163 42585
rect 15212 42588 15594 42616
rect 12529 42551 12587 42557
rect 12529 42548 12541 42551
rect 12492 42520 12541 42548
rect 12492 42508 12498 42520
rect 12529 42517 12541 42520
rect 12575 42517 12587 42551
rect 12529 42511 12587 42517
rect 12618 42508 12624 42560
rect 12676 42548 12682 42560
rect 12805 42551 12863 42557
rect 12805 42548 12817 42551
rect 12676 42520 12817 42548
rect 12676 42508 12682 42520
rect 12805 42517 12817 42520
rect 12851 42548 12863 42551
rect 13722 42548 13728 42560
rect 12851 42520 13728 42548
rect 12851 42517 12863 42520
rect 12805 42511 12863 42517
rect 13722 42508 13728 42520
rect 13780 42548 13786 42560
rect 14277 42551 14335 42557
rect 14277 42548 14289 42551
rect 13780 42520 14289 42548
rect 13780 42508 13786 42520
rect 14277 42517 14289 42520
rect 14323 42548 14335 42551
rect 15010 42548 15016 42560
rect 14323 42520 15016 42548
rect 14323 42517 14335 42520
rect 14277 42511 14335 42517
rect 15010 42508 15016 42520
rect 15068 42548 15074 42560
rect 15212 42548 15240 42588
rect 17497 42585 17509 42619
rect 17543 42616 17555 42619
rect 19794 42616 19800 42628
rect 17543 42588 19800 42616
rect 17543 42585 17555 42588
rect 17497 42579 17555 42585
rect 19794 42576 19800 42588
rect 19852 42576 19858 42628
rect 20530 42576 20536 42628
rect 20588 42576 20594 42628
rect 22940 42616 22968 42724
rect 25130 42712 25136 42724
rect 25188 42712 25194 42764
rect 23201 42687 23259 42693
rect 23201 42653 23213 42687
rect 23247 42653 23259 42687
rect 23201 42647 23259 42653
rect 23477 42687 23535 42693
rect 23477 42653 23489 42687
rect 23523 42684 23535 42687
rect 23658 42684 23664 42696
rect 23523 42656 23664 42684
rect 23523 42653 23535 42656
rect 23477 42647 23535 42653
rect 21100 42588 22968 42616
rect 23216 42616 23244 42647
rect 23658 42644 23664 42656
rect 23716 42644 23722 42696
rect 23750 42644 23756 42696
rect 23808 42684 23814 42696
rect 24854 42684 24860 42696
rect 23808 42656 24860 42684
rect 23808 42644 23814 42656
rect 24854 42644 24860 42656
rect 24912 42644 24918 42696
rect 23216 42588 24532 42616
rect 15068 42520 15240 42548
rect 16577 42551 16635 42557
rect 15068 42508 15074 42520
rect 16577 42517 16589 42551
rect 16623 42548 16635 42551
rect 16758 42548 16764 42560
rect 16623 42520 16764 42548
rect 16623 42517 16635 42520
rect 16577 42511 16635 42517
rect 16758 42508 16764 42520
rect 16816 42508 16822 42560
rect 17589 42551 17647 42557
rect 17589 42517 17601 42551
rect 17635 42548 17647 42551
rect 19150 42548 19156 42560
rect 17635 42520 19156 42548
rect 17635 42517 17647 42520
rect 17589 42511 17647 42517
rect 19150 42508 19156 42520
rect 19208 42548 19214 42560
rect 21100 42548 21128 42588
rect 19208 42520 21128 42548
rect 19208 42508 19214 42520
rect 21266 42508 21272 42560
rect 21324 42508 21330 42560
rect 21818 42508 21824 42560
rect 21876 42508 21882 42560
rect 22186 42508 22192 42560
rect 22244 42508 22250 42560
rect 24504 42557 24532 42588
rect 24578 42576 24584 42628
rect 24636 42616 24642 42628
rect 25317 42619 25375 42625
rect 25317 42616 25329 42619
rect 24636 42588 25329 42616
rect 24636 42576 24642 42588
rect 25317 42585 25329 42588
rect 25363 42585 25375 42619
rect 25317 42579 25375 42585
rect 24489 42551 24547 42557
rect 24489 42517 24501 42551
rect 24535 42548 24547 42551
rect 24854 42548 24860 42560
rect 24535 42520 24860 42548
rect 24535 42517 24547 42520
rect 24489 42511 24547 42517
rect 24854 42508 24860 42520
rect 24912 42508 24918 42560
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 4338 42304 4344 42356
rect 4396 42304 4402 42356
rect 5074 42304 5080 42356
rect 5132 42304 5138 42356
rect 6733 42347 6791 42353
rect 6733 42344 6745 42347
rect 5184 42316 6745 42344
rect 4154 42236 4160 42288
rect 4212 42276 4218 42288
rect 5184 42276 5212 42316
rect 6733 42313 6745 42316
rect 6779 42313 6791 42347
rect 8478 42344 8484 42356
rect 6733 42307 6791 42313
rect 7576 42316 8484 42344
rect 6641 42279 6699 42285
rect 6641 42276 6653 42279
rect 4212 42248 5212 42276
rect 6564 42248 6653 42276
rect 4212 42236 4218 42248
rect 3881 42211 3939 42217
rect 3881 42177 3893 42211
rect 3927 42208 3939 42211
rect 4246 42208 4252 42220
rect 3927 42180 4252 42208
rect 3927 42177 3939 42180
rect 3881 42171 3939 42177
rect 4246 42168 4252 42180
rect 4304 42168 4310 42220
rect 4985 42211 5043 42217
rect 4985 42177 4997 42211
rect 5031 42208 5043 42211
rect 5031 42180 5580 42208
rect 5031 42177 5043 42180
rect 4985 42171 5043 42177
rect 5552 42013 5580 42180
rect 6564 42140 6592 42248
rect 6641 42245 6653 42248
rect 6687 42245 6699 42279
rect 7576 42276 7604 42316
rect 8478 42304 8484 42316
rect 8536 42344 8542 42356
rect 10226 42344 10232 42356
rect 8536 42316 10232 42344
rect 8536 42304 8542 42316
rect 10226 42304 10232 42316
rect 10284 42304 10290 42356
rect 11790 42304 11796 42356
rect 11848 42304 11854 42356
rect 12989 42347 13047 42353
rect 12989 42313 13001 42347
rect 13035 42344 13047 42347
rect 13446 42344 13452 42356
rect 13035 42316 13452 42344
rect 13035 42313 13047 42316
rect 12989 42307 13047 42313
rect 13446 42304 13452 42316
rect 13504 42304 13510 42356
rect 15194 42304 15200 42356
rect 15252 42344 15258 42356
rect 15381 42347 15439 42353
rect 15381 42344 15393 42347
rect 15252 42316 15393 42344
rect 15252 42304 15258 42316
rect 15381 42313 15393 42316
rect 15427 42313 15439 42347
rect 15381 42307 15439 42313
rect 15841 42347 15899 42353
rect 15841 42313 15853 42347
rect 15887 42344 15899 42347
rect 16853 42347 16911 42353
rect 16853 42344 16865 42347
rect 15887 42316 16865 42344
rect 15887 42313 15899 42316
rect 15841 42307 15899 42313
rect 16853 42313 16865 42316
rect 16899 42313 16911 42347
rect 16853 42307 16911 42313
rect 17221 42347 17279 42353
rect 17221 42313 17233 42347
rect 17267 42344 17279 42347
rect 19610 42344 19616 42356
rect 17267 42316 19616 42344
rect 17267 42313 17279 42316
rect 17221 42307 17279 42313
rect 19610 42304 19616 42316
rect 19668 42344 19674 42356
rect 19668 42316 20668 42344
rect 19668 42304 19674 42316
rect 12253 42279 12311 42285
rect 6641 42239 6699 42245
rect 7484 42248 7604 42276
rect 9048 42248 10272 42276
rect 6730 42168 6736 42220
rect 6788 42208 6794 42220
rect 7484 42217 7512 42248
rect 7469 42211 7527 42217
rect 7469 42208 7481 42211
rect 6788 42180 7481 42208
rect 6788 42168 6794 42180
rect 7469 42177 7481 42180
rect 7515 42177 7527 42211
rect 7469 42171 7527 42177
rect 8846 42168 8852 42220
rect 8904 42168 8910 42220
rect 9048 42208 9076 42248
rect 8956 42180 9076 42208
rect 10045 42211 10103 42217
rect 6564 42112 6914 42140
rect 5537 42007 5595 42013
rect 5537 41973 5549 42007
rect 5583 42004 5595 42007
rect 6270 42004 6276 42016
rect 5583 41976 6276 42004
rect 5583 41973 5595 41976
rect 5537 41967 5595 41973
rect 6270 41964 6276 41976
rect 6328 41964 6334 42016
rect 6886 42004 6914 42112
rect 7742 42100 7748 42152
rect 7800 42140 7806 42152
rect 8956 42140 8984 42180
rect 10045 42177 10057 42211
rect 10091 42177 10103 42211
rect 10045 42171 10103 42177
rect 7800 42112 8984 42140
rect 7800 42100 7806 42112
rect 10060 42072 10088 42171
rect 10134 42100 10140 42152
rect 10192 42100 10198 42152
rect 10244 42149 10272 42248
rect 12253 42245 12265 42279
rect 12299 42276 12311 42279
rect 15102 42276 15108 42288
rect 12299 42248 15108 42276
rect 12299 42245 12311 42248
rect 12253 42239 12311 42245
rect 15102 42236 15108 42248
rect 15160 42236 15166 42288
rect 20640 42276 20668 42316
rect 20714 42304 20720 42356
rect 20772 42304 20778 42356
rect 20898 42304 20904 42356
rect 20956 42344 20962 42356
rect 21269 42347 21327 42353
rect 21269 42344 21281 42347
rect 20956 42316 21281 42344
rect 20956 42304 20962 42316
rect 21269 42313 21281 42316
rect 21315 42313 21327 42347
rect 21269 42307 21327 42313
rect 23382 42304 23388 42356
rect 23440 42344 23446 42356
rect 25225 42347 25283 42353
rect 25225 42344 25237 42347
rect 23440 42316 25237 42344
rect 23440 42304 23446 42316
rect 25225 42313 25237 42316
rect 25271 42313 25283 42347
rect 25225 42307 25283 42313
rect 23750 42276 23756 42288
rect 16040 42248 17448 42276
rect 20640 42248 23756 42276
rect 11146 42168 11152 42220
rect 11204 42208 11210 42220
rect 12161 42211 12219 42217
rect 12161 42208 12173 42211
rect 11204 42180 12173 42208
rect 11204 42168 11210 42180
rect 12161 42177 12173 42180
rect 12207 42177 12219 42211
rect 12161 42171 12219 42177
rect 13357 42211 13415 42217
rect 13357 42177 13369 42211
rect 13403 42208 13415 42211
rect 14185 42211 14243 42217
rect 14185 42208 14197 42211
rect 13403 42180 14197 42208
rect 13403 42177 13415 42180
rect 13357 42171 13415 42177
rect 14185 42177 14197 42180
rect 14231 42177 14243 42211
rect 14185 42171 14243 42177
rect 15746 42168 15752 42220
rect 15804 42168 15810 42220
rect 10229 42143 10287 42149
rect 10229 42109 10241 42143
rect 10275 42109 10287 42143
rect 10229 42103 10287 42109
rect 12434 42100 12440 42152
rect 12492 42100 12498 42152
rect 12526 42100 12532 42152
rect 12584 42140 12590 42152
rect 13449 42143 13507 42149
rect 13449 42140 13461 42143
rect 12584 42112 13461 42140
rect 12584 42100 12590 42112
rect 13449 42109 13461 42112
rect 13495 42109 13507 42143
rect 13449 42103 13507 42109
rect 13633 42143 13691 42149
rect 13633 42109 13645 42143
rect 13679 42109 13691 42143
rect 13633 42103 13691 42109
rect 15933 42143 15991 42149
rect 15933 42109 15945 42143
rect 15979 42109 15991 42143
rect 15933 42103 15991 42109
rect 9048 42044 10088 42072
rect 13648 42072 13676 42103
rect 14182 42072 14188 42084
rect 13648 42044 14188 42072
rect 7190 42004 7196 42016
rect 6886 41976 7196 42004
rect 7190 41964 7196 41976
rect 7248 41964 7254 42016
rect 7558 41964 7564 42016
rect 7616 42004 7622 42016
rect 9048 42004 9076 42044
rect 14182 42032 14188 42044
rect 14240 42072 14246 42084
rect 15948 42072 15976 42103
rect 14240 42044 15976 42072
rect 14240 42032 14246 42044
rect 7616 41976 9076 42004
rect 7616 41964 7622 41976
rect 9214 41964 9220 42016
rect 9272 41964 9278 42016
rect 9306 41964 9312 42016
rect 9364 42004 9370 42016
rect 9677 42007 9735 42013
rect 9677 42004 9689 42007
rect 9364 41976 9689 42004
rect 9364 41964 9370 41976
rect 9677 41973 9689 41976
rect 9723 41973 9735 42007
rect 9677 41967 9735 41973
rect 10778 41964 10784 42016
rect 10836 41964 10842 42016
rect 13446 41964 13452 42016
rect 13504 42004 13510 42016
rect 13630 42004 13636 42016
rect 13504 41976 13636 42004
rect 13504 41964 13510 41976
rect 13630 41964 13636 41976
rect 13688 42004 13694 42016
rect 16040 42004 16068 42248
rect 17420 42149 17448 42248
rect 23750 42236 23756 42248
rect 23808 42236 23814 42288
rect 24486 42236 24492 42288
rect 24544 42236 24550 42288
rect 18877 42211 18935 42217
rect 18877 42177 18889 42211
rect 18923 42177 18935 42211
rect 18877 42171 18935 42177
rect 17313 42143 17371 42149
rect 17313 42140 17325 42143
rect 16546 42112 17325 42140
rect 13688 41976 16068 42004
rect 13688 41964 13694 41976
rect 16390 41964 16396 42016
rect 16448 42004 16454 42016
rect 16546 42004 16574 42112
rect 17313 42109 17325 42112
rect 17359 42109 17371 42143
rect 17313 42103 17371 42109
rect 17405 42143 17463 42149
rect 17405 42109 17417 42143
rect 17451 42109 17463 42143
rect 17405 42103 17463 42109
rect 18892 42072 18920 42171
rect 20622 42168 20628 42220
rect 20680 42168 20686 42220
rect 22005 42211 22063 42217
rect 22005 42208 22017 42211
rect 21560 42180 22017 42208
rect 19242 42100 19248 42152
rect 19300 42140 19306 42152
rect 19613 42143 19671 42149
rect 19613 42140 19625 42143
rect 19300 42112 19625 42140
rect 19300 42100 19306 42112
rect 19613 42109 19625 42112
rect 19659 42109 19671 42143
rect 19613 42103 19671 42109
rect 19978 42100 19984 42152
rect 20036 42140 20042 42152
rect 20809 42143 20867 42149
rect 20809 42140 20821 42143
rect 20036 42112 20821 42140
rect 20036 42100 20042 42112
rect 20809 42109 20821 42112
rect 20855 42140 20867 42143
rect 21266 42140 21272 42152
rect 20855 42112 21272 42140
rect 20855 42109 20867 42112
rect 20809 42103 20867 42109
rect 21266 42100 21272 42112
rect 21324 42100 21330 42152
rect 21560 42081 21588 42180
rect 22005 42177 22017 42180
rect 22051 42177 22063 42211
rect 22005 42171 22063 42177
rect 22278 42100 22284 42152
rect 22336 42140 22342 42152
rect 22830 42140 22836 42152
rect 22336 42112 22836 42140
rect 22336 42100 22342 42112
rect 22830 42100 22836 42112
rect 22888 42140 22894 42152
rect 23474 42140 23480 42152
rect 22888 42112 23480 42140
rect 22888 42100 22894 42112
rect 23474 42100 23480 42112
rect 23532 42100 23538 42152
rect 23753 42143 23811 42149
rect 23753 42109 23765 42143
rect 23799 42140 23811 42143
rect 25498 42140 25504 42152
rect 23799 42112 25504 42140
rect 23799 42109 23811 42112
rect 23753 42103 23811 42109
rect 25498 42100 25504 42112
rect 25556 42100 25562 42152
rect 21545 42075 21603 42081
rect 21545 42072 21557 42075
rect 18524 42044 21557 42072
rect 16448 41976 16574 42004
rect 16448 41964 16454 41976
rect 18322 41964 18328 42016
rect 18380 42004 18386 42016
rect 18524 42013 18552 42044
rect 21545 42041 21557 42044
rect 21591 42041 21603 42075
rect 21545 42035 21603 42041
rect 18509 42007 18567 42013
rect 18509 42004 18521 42007
rect 18380 41976 18521 42004
rect 18380 41964 18386 41976
rect 18509 41973 18521 41976
rect 18555 41973 18567 42007
rect 18509 41967 18567 41973
rect 20254 41964 20260 42016
rect 20312 41964 20318 42016
rect 24854 41964 24860 42016
rect 24912 42004 24918 42016
rect 25038 42004 25044 42016
rect 24912 41976 25044 42004
rect 24912 41964 24918 41976
rect 25038 41964 25044 41976
rect 25096 41964 25102 42016
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 5166 41760 5172 41812
rect 5224 41760 5230 41812
rect 7653 41803 7711 41809
rect 7653 41769 7665 41803
rect 7699 41800 7711 41803
rect 7742 41800 7748 41812
rect 7699 41772 7748 41800
rect 7699 41769 7711 41772
rect 7653 41763 7711 41769
rect 7742 41760 7748 41772
rect 7800 41760 7806 41812
rect 8021 41803 8079 41809
rect 8021 41769 8033 41803
rect 8067 41800 8079 41803
rect 8294 41800 8300 41812
rect 8067 41772 8300 41800
rect 8067 41769 8079 41772
rect 8021 41763 8079 41769
rect 5905 41667 5963 41673
rect 5905 41633 5917 41667
rect 5951 41664 5963 41667
rect 6178 41664 6184 41676
rect 5951 41636 6184 41664
rect 5951 41633 5963 41636
rect 5905 41627 5963 41633
rect 6178 41624 6184 41636
rect 6236 41664 6242 41676
rect 6730 41664 6736 41676
rect 6236 41636 6736 41664
rect 6236 41624 6242 41636
rect 6730 41624 6736 41636
rect 6788 41624 6794 41676
rect 8036 41596 8064 41763
rect 8294 41760 8300 41772
rect 8352 41800 8358 41812
rect 8846 41800 8852 41812
rect 8352 41772 8852 41800
rect 8352 41760 8358 41772
rect 8846 41760 8852 41772
rect 8904 41760 8910 41812
rect 10689 41803 10747 41809
rect 10689 41769 10701 41803
rect 10735 41800 10747 41803
rect 11054 41800 11060 41812
rect 10735 41772 11060 41800
rect 10735 41769 10747 41772
rect 10689 41763 10747 41769
rect 11054 41760 11060 41772
rect 11112 41760 11118 41812
rect 14458 41760 14464 41812
rect 14516 41800 14522 41812
rect 16390 41800 16396 41812
rect 14516 41772 16396 41800
rect 14516 41760 14522 41772
rect 16390 41760 16396 41772
rect 16448 41760 16454 41812
rect 17310 41760 17316 41812
rect 17368 41800 17374 41812
rect 17368 41772 21128 41800
rect 17368 41760 17374 41772
rect 9214 41692 9220 41744
rect 9272 41732 9278 41744
rect 10870 41732 10876 41744
rect 9272 41704 10876 41732
rect 9272 41692 9278 41704
rect 10870 41692 10876 41704
rect 10928 41692 10934 41744
rect 15746 41692 15752 41744
rect 15804 41732 15810 41744
rect 19334 41732 19340 41744
rect 15804 41704 19340 41732
rect 15804 41692 15810 41704
rect 19334 41692 19340 41704
rect 19392 41692 19398 41744
rect 21100 41732 21128 41772
rect 21174 41760 21180 41812
rect 21232 41760 21238 41812
rect 23198 41800 23204 41812
rect 21284 41772 23204 41800
rect 21284 41732 21312 41772
rect 23198 41760 23204 41772
rect 23256 41800 23262 41812
rect 25314 41800 25320 41812
rect 23256 41772 25320 41800
rect 23256 41760 23262 41772
rect 25314 41760 25320 41772
rect 25372 41760 25378 41812
rect 21100 41704 21312 41732
rect 21637 41735 21695 41741
rect 21637 41701 21649 41735
rect 21683 41732 21695 41735
rect 22554 41732 22560 41744
rect 21683 41704 22560 41732
rect 21683 41701 21695 41704
rect 21637 41695 21695 41701
rect 22554 41692 22560 41704
rect 22612 41692 22618 41744
rect 22833 41735 22891 41741
rect 22833 41701 22845 41735
rect 22879 41732 22891 41735
rect 25038 41732 25044 41744
rect 22879 41704 25044 41732
rect 22879 41701 22891 41704
rect 22833 41695 22891 41701
rect 25038 41692 25044 41704
rect 25096 41692 25102 41744
rect 10137 41667 10195 41673
rect 10137 41633 10149 41667
rect 10183 41664 10195 41667
rect 10226 41664 10232 41676
rect 10183 41636 10232 41664
rect 10183 41633 10195 41636
rect 10137 41627 10195 41633
rect 10226 41624 10232 41636
rect 10284 41624 10290 41676
rect 10686 41624 10692 41676
rect 10744 41664 10750 41676
rect 11241 41667 11299 41673
rect 11241 41664 11253 41667
rect 10744 41636 11253 41664
rect 10744 41624 10750 41636
rect 11241 41633 11253 41636
rect 11287 41633 11299 41667
rect 11241 41627 11299 41633
rect 12342 41624 12348 41676
rect 12400 41664 12406 41676
rect 12713 41667 12771 41673
rect 12713 41664 12725 41667
rect 12400 41636 12725 41664
rect 12400 41624 12406 41636
rect 12713 41633 12725 41636
rect 12759 41664 12771 41667
rect 12802 41664 12808 41676
rect 12759 41636 12808 41664
rect 12759 41633 12771 41636
rect 12713 41627 12771 41633
rect 12802 41624 12808 41636
rect 12860 41664 12866 41676
rect 13630 41664 13636 41676
rect 12860 41636 13636 41664
rect 12860 41624 12866 41636
rect 13630 41624 13636 41636
rect 13688 41624 13694 41676
rect 15194 41624 15200 41676
rect 15252 41664 15258 41676
rect 16114 41664 16120 41676
rect 15252 41636 16120 41664
rect 15252 41624 15258 41636
rect 16114 41624 16120 41636
rect 16172 41664 16178 41676
rect 16761 41667 16819 41673
rect 16761 41664 16773 41667
rect 16172 41636 16773 41664
rect 16172 41624 16178 41636
rect 16761 41633 16773 41636
rect 16807 41633 16819 41667
rect 16761 41627 16819 41633
rect 18506 41624 18512 41676
rect 18564 41664 18570 41676
rect 18601 41667 18659 41673
rect 18601 41664 18613 41667
rect 18564 41636 18613 41664
rect 18564 41624 18570 41636
rect 18601 41633 18613 41636
rect 18647 41633 18659 41667
rect 18601 41627 18659 41633
rect 18785 41667 18843 41673
rect 18785 41633 18797 41667
rect 18831 41664 18843 41667
rect 18966 41664 18972 41676
rect 18831 41636 18972 41664
rect 18831 41633 18843 41636
rect 18785 41627 18843 41633
rect 18966 41624 18972 41636
rect 19024 41624 19030 41676
rect 19242 41624 19248 41676
rect 19300 41664 19306 41676
rect 19429 41667 19487 41673
rect 19429 41664 19441 41667
rect 19300 41636 19441 41664
rect 19300 41624 19306 41636
rect 19429 41633 19441 41636
rect 19475 41633 19487 41667
rect 20898 41664 20904 41676
rect 19429 41627 19487 41633
rect 20824 41636 20904 41664
rect 7314 41568 8064 41596
rect 10318 41556 10324 41608
rect 10376 41596 10382 41608
rect 11882 41596 11888 41608
rect 10376 41568 11888 41596
rect 10376 41556 10382 41568
rect 11882 41556 11888 41568
rect 11940 41556 11946 41608
rect 16666 41556 16672 41608
rect 16724 41556 16730 41608
rect 17494 41556 17500 41608
rect 17552 41596 17558 41608
rect 17552 41568 19472 41596
rect 20824 41582 20852 41636
rect 20898 41624 20904 41636
rect 20956 41624 20962 41676
rect 22281 41667 22339 41673
rect 22281 41633 22293 41667
rect 22327 41664 22339 41667
rect 22462 41664 22468 41676
rect 22327 41636 22468 41664
rect 22327 41633 22339 41636
rect 22281 41627 22339 41633
rect 22462 41624 22468 41636
rect 22520 41624 22526 41676
rect 23290 41624 23296 41676
rect 23348 41624 23354 41676
rect 23385 41667 23443 41673
rect 23385 41633 23397 41667
rect 23431 41664 23443 41667
rect 23474 41664 23480 41676
rect 23431 41636 23480 41664
rect 23431 41633 23443 41636
rect 23385 41627 23443 41633
rect 23474 41624 23480 41636
rect 23532 41624 23538 41676
rect 23566 41624 23572 41676
rect 23624 41664 23630 41676
rect 25682 41664 25688 41676
rect 23624 41636 25688 41664
rect 23624 41624 23630 41636
rect 25682 41624 25688 41636
rect 25740 41624 25746 41676
rect 24673 41599 24731 41605
rect 17552 41556 17558 41568
rect 5077 41531 5135 41537
rect 5077 41497 5089 41531
rect 5123 41528 5135 41531
rect 6181 41531 6239 41537
rect 5123 41500 5672 41528
rect 5123 41497 5135 41500
rect 5077 41491 5135 41497
rect 5644 41469 5672 41500
rect 6181 41497 6193 41531
rect 6227 41497 6239 41531
rect 6181 41491 6239 41497
rect 9309 41531 9367 41537
rect 9309 41497 9321 41531
rect 9355 41528 9367 41531
rect 10410 41528 10416 41540
rect 9355 41500 10416 41528
rect 9355 41497 9367 41500
rect 9309 41491 9367 41497
rect 5629 41463 5687 41469
rect 5629 41429 5641 41463
rect 5675 41460 5687 41463
rect 5718 41460 5724 41472
rect 5675 41432 5724 41460
rect 5675 41429 5687 41432
rect 5629 41423 5687 41429
rect 5718 41420 5724 41432
rect 5776 41420 5782 41472
rect 6196 41460 6224 41491
rect 10410 41488 10416 41500
rect 10468 41528 10474 41540
rect 10778 41528 10784 41540
rect 10468 41500 10784 41528
rect 10468 41488 10474 41500
rect 10778 41488 10784 41500
rect 10836 41528 10842 41540
rect 11977 41531 12035 41537
rect 11977 41528 11989 41531
rect 10836 41500 11989 41528
rect 10836 41488 10842 41500
rect 11977 41497 11989 41500
rect 12023 41528 12035 41531
rect 13265 41531 13323 41537
rect 13265 41528 13277 41531
rect 12023 41500 13277 41528
rect 12023 41497 12035 41500
rect 11977 41491 12035 41497
rect 13265 41497 13277 41500
rect 13311 41528 13323 41531
rect 18322 41528 18328 41540
rect 13311 41500 18328 41528
rect 13311 41497 13323 41500
rect 13265 41491 13323 41497
rect 18322 41488 18328 41500
rect 18380 41488 18386 41540
rect 19444 41528 19472 41568
rect 24673 41565 24685 41599
rect 24719 41596 24731 41599
rect 25314 41596 25320 41608
rect 24719 41568 25320 41596
rect 24719 41565 24731 41568
rect 24673 41559 24731 41565
rect 25314 41556 25320 41568
rect 25372 41556 25378 41608
rect 19705 41531 19763 41537
rect 19705 41528 19717 41531
rect 19444 41500 19717 41528
rect 19705 41497 19717 41500
rect 19751 41528 19763 41531
rect 19978 41528 19984 41540
rect 19751 41500 19984 41528
rect 19751 41497 19763 41500
rect 19705 41491 19763 41497
rect 19978 41488 19984 41500
rect 20036 41488 20042 41540
rect 21082 41488 21088 41540
rect 21140 41528 21146 41540
rect 22097 41531 22155 41537
rect 22097 41528 22109 41531
rect 21140 41500 22109 41528
rect 21140 41488 21146 41500
rect 22097 41497 22109 41500
rect 22143 41497 22155 41531
rect 22097 41491 22155 41497
rect 22278 41488 22284 41540
rect 22336 41528 22342 41540
rect 23201 41531 23259 41537
rect 23201 41528 23213 41531
rect 22336 41500 23213 41528
rect 22336 41488 22342 41500
rect 23201 41497 23213 41500
rect 23247 41497 23259 41531
rect 23201 41491 23259 41497
rect 24489 41531 24547 41537
rect 24489 41497 24501 41531
rect 24535 41528 24547 41531
rect 24535 41500 25360 41528
rect 24535 41497 24547 41500
rect 24489 41491 24547 41497
rect 25332 41472 25360 41500
rect 7006 41460 7012 41472
rect 6196 41432 7012 41460
rect 7006 41420 7012 41432
rect 7064 41420 7070 41472
rect 11054 41420 11060 41472
rect 11112 41420 11118 41472
rect 11149 41463 11207 41469
rect 11149 41429 11161 41463
rect 11195 41460 11207 41463
rect 14182 41460 14188 41472
rect 11195 41432 14188 41460
rect 11195 41429 11207 41432
rect 11149 41423 11207 41429
rect 14182 41420 14188 41432
rect 14240 41420 14246 41472
rect 16209 41463 16267 41469
rect 16209 41429 16221 41463
rect 16255 41460 16267 41463
rect 16482 41460 16488 41472
rect 16255 41432 16488 41460
rect 16255 41429 16267 41432
rect 16209 41423 16267 41429
rect 16482 41420 16488 41432
rect 16540 41420 16546 41472
rect 16577 41463 16635 41469
rect 16577 41429 16589 41463
rect 16623 41460 16635 41463
rect 17310 41460 17316 41472
rect 16623 41432 17316 41460
rect 16623 41429 16635 41432
rect 16577 41423 16635 41429
rect 17310 41420 17316 41432
rect 17368 41420 17374 41472
rect 18141 41463 18199 41469
rect 18141 41429 18153 41463
rect 18187 41460 18199 41463
rect 18414 41460 18420 41472
rect 18187 41432 18420 41460
rect 18187 41429 18199 41432
rect 18141 41423 18199 41429
rect 18414 41420 18420 41432
rect 18472 41420 18478 41472
rect 18509 41463 18567 41469
rect 18509 41429 18521 41463
rect 18555 41460 18567 41463
rect 18874 41460 18880 41472
rect 18555 41432 18880 41460
rect 18555 41429 18567 41432
rect 18509 41423 18567 41429
rect 18874 41420 18880 41432
rect 18932 41420 18938 41472
rect 22002 41420 22008 41472
rect 22060 41420 22066 41472
rect 24578 41420 24584 41472
rect 24636 41460 24642 41472
rect 24857 41463 24915 41469
rect 24857 41460 24869 41463
rect 24636 41432 24869 41460
rect 24636 41420 24642 41432
rect 24857 41429 24869 41432
rect 24903 41429 24915 41463
rect 24857 41423 24915 41429
rect 25130 41420 25136 41472
rect 25188 41420 25194 41472
rect 25314 41420 25320 41472
rect 25372 41420 25378 41472
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 3326 41216 3332 41268
rect 3384 41216 3390 41268
rect 11698 41216 11704 41268
rect 11756 41216 11762 41268
rect 12161 41259 12219 41265
rect 12161 41225 12173 41259
rect 12207 41256 12219 41259
rect 14918 41256 14924 41268
rect 12207 41228 14924 41256
rect 12207 41225 12219 41228
rect 12161 41219 12219 41225
rect 14918 41216 14924 41228
rect 14976 41216 14982 41268
rect 19242 41256 19248 41268
rect 16868 41228 19248 41256
rect 9122 41188 9128 41200
rect 8956 41160 9128 41188
rect 1302 41080 1308 41132
rect 1360 41120 1366 41132
rect 1765 41123 1823 41129
rect 1765 41120 1777 41123
rect 1360 41092 1777 41120
rect 1360 41080 1366 41092
rect 1765 41089 1777 41092
rect 1811 41120 1823 41123
rect 2041 41123 2099 41129
rect 2041 41120 2053 41123
rect 1811 41092 2053 41120
rect 1811 41089 1823 41092
rect 1765 41083 1823 41089
rect 2041 41089 2053 41092
rect 2087 41089 2099 41123
rect 2041 41083 2099 41089
rect 3237 41123 3295 41129
rect 3237 41089 3249 41123
rect 3283 41120 3295 41123
rect 3697 41123 3755 41129
rect 3697 41120 3709 41123
rect 3283 41092 3709 41120
rect 3283 41089 3295 41092
rect 3237 41083 3295 41089
rect 3697 41089 3709 41092
rect 3743 41120 3755 41123
rect 4614 41120 4620 41132
rect 3743 41092 4620 41120
rect 3743 41089 3755 41092
rect 3697 41083 3755 41089
rect 4614 41080 4620 41092
rect 4672 41080 4678 41132
rect 8956 41129 8984 41160
rect 9122 41148 9128 41160
rect 9180 41148 9186 41200
rect 8941 41123 8999 41129
rect 8941 41089 8953 41123
rect 8987 41089 8999 41123
rect 10350 41092 11100 41120
rect 8941 41083 8999 41089
rect 9217 41055 9275 41061
rect 9217 41021 9229 41055
rect 9263 41052 9275 41055
rect 10870 41052 10876 41064
rect 9263 41024 10876 41052
rect 9263 41021 9275 41024
rect 9217 41015 9275 41021
rect 10870 41012 10876 41024
rect 10928 41012 10934 41064
rect 1578 40876 1584 40928
rect 1636 40876 1642 40928
rect 9950 40876 9956 40928
rect 10008 40916 10014 40928
rect 10686 40916 10692 40928
rect 10008 40888 10692 40916
rect 10008 40876 10014 40888
rect 10686 40876 10692 40888
rect 10744 40876 10750 40928
rect 11072 40925 11100 41092
rect 12066 41080 12072 41132
rect 12124 41080 12130 41132
rect 13630 41080 13636 41132
rect 13688 41080 13694 41132
rect 15010 41080 15016 41132
rect 15068 41120 15074 41132
rect 16868 41129 16896 41228
rect 19242 41216 19248 41228
rect 19300 41216 19306 41268
rect 19797 41259 19855 41265
rect 19797 41225 19809 41259
rect 19843 41256 19855 41259
rect 20162 41256 20168 41268
rect 19843 41228 20168 41256
rect 19843 41225 19855 41228
rect 19797 41219 19855 41225
rect 20162 41216 20168 41228
rect 20220 41216 20226 41268
rect 21082 41216 21088 41268
rect 21140 41256 21146 41268
rect 21542 41256 21548 41268
rect 21140 41228 21548 41256
rect 21140 41216 21146 41228
rect 21542 41216 21548 41228
rect 21600 41216 21606 41268
rect 22002 41216 22008 41268
rect 22060 41216 22066 41268
rect 23474 41216 23480 41268
rect 23532 41256 23538 41268
rect 24673 41259 24731 41265
rect 24673 41256 24685 41259
rect 23532 41228 24685 41256
rect 23532 41216 23538 41228
rect 24673 41225 24685 41228
rect 24719 41225 24731 41259
rect 24673 41219 24731 41225
rect 18414 41188 18420 41200
rect 18354 41160 18420 41188
rect 18414 41148 18420 41160
rect 18472 41188 18478 41200
rect 18877 41191 18935 41197
rect 18877 41188 18889 41191
rect 18472 41160 18889 41188
rect 18472 41148 18478 41160
rect 18877 41157 18889 41160
rect 18923 41157 18935 41191
rect 18877 41151 18935 41157
rect 19886 41148 19892 41200
rect 19944 41148 19950 41200
rect 21008 41160 22094 41188
rect 16853 41123 16911 41129
rect 15068 41092 15792 41120
rect 15068 41080 15074 41092
rect 12250 41012 12256 41064
rect 12308 41012 12314 41064
rect 13909 41055 13967 41061
rect 13909 41021 13921 41055
rect 13955 41052 13967 41055
rect 13998 41052 14004 41064
rect 13955 41024 14004 41052
rect 13955 41021 13967 41024
rect 13909 41015 13967 41021
rect 13998 41012 14004 41024
rect 14056 41052 14062 41064
rect 15194 41052 15200 41064
rect 14056 41024 15200 41052
rect 14056 41012 14062 41024
rect 15194 41012 15200 41024
rect 15252 41012 15258 41064
rect 11057 40919 11115 40925
rect 11057 40885 11069 40919
rect 11103 40916 11115 40919
rect 11330 40916 11336 40928
rect 11103 40888 11336 40916
rect 11103 40885 11115 40888
rect 11057 40879 11115 40885
rect 11330 40876 11336 40888
rect 11388 40916 11394 40928
rect 12250 40916 12256 40928
rect 11388 40888 12256 40916
rect 11388 40876 11394 40888
rect 12250 40876 12256 40888
rect 12308 40916 12314 40928
rect 12618 40916 12624 40928
rect 12308 40888 12624 40916
rect 12308 40876 12314 40888
rect 12618 40876 12624 40888
rect 12676 40876 12682 40928
rect 15381 40919 15439 40925
rect 15381 40885 15393 40919
rect 15427 40916 15439 40919
rect 15562 40916 15568 40928
rect 15427 40888 15568 40916
rect 15427 40885 15439 40888
rect 15381 40879 15439 40885
rect 15562 40876 15568 40888
rect 15620 40876 15626 40928
rect 15764 40925 15792 41092
rect 16853 41089 16865 41123
rect 16899 41089 16911 41123
rect 16853 41083 16911 41089
rect 18598 41080 18604 41132
rect 18656 41120 18662 41132
rect 21008 41120 21036 41160
rect 18656 41092 21036 41120
rect 18656 41080 18662 41092
rect 21082 41080 21088 41132
rect 21140 41080 21146 41132
rect 16758 41012 16764 41064
rect 16816 41052 16822 41064
rect 17129 41055 17187 41061
rect 17129 41052 17141 41055
rect 16816 41024 17141 41052
rect 16816 41012 16822 41024
rect 17129 41021 17141 41024
rect 17175 41052 17187 41055
rect 17175 41024 18460 41052
rect 17175 41021 17187 41024
rect 17129 41015 17187 41021
rect 18432 40984 18460 41024
rect 19702 41012 19708 41064
rect 19760 41052 19766 41064
rect 19978 41052 19984 41064
rect 19760 41024 19984 41052
rect 19760 41012 19766 41024
rect 19978 41012 19984 41024
rect 20036 41012 20042 41064
rect 20714 41012 20720 41064
rect 20772 41052 20778 41064
rect 20990 41052 20996 41064
rect 20772 41024 20996 41052
rect 20772 41012 20778 41024
rect 20990 41012 20996 41024
rect 21048 41052 21054 41064
rect 21177 41055 21235 41061
rect 21177 41052 21189 41055
rect 21048 41024 21189 41052
rect 21048 41012 21054 41024
rect 21177 41021 21189 41024
rect 21223 41021 21235 41055
rect 21177 41015 21235 41021
rect 21269 41055 21327 41061
rect 21269 41021 21281 41055
rect 21315 41021 21327 41055
rect 21269 41015 21327 41021
rect 21284 40984 21312 41015
rect 18432 40956 21312 40984
rect 22066 40984 22094 41160
rect 22370 41148 22376 41200
rect 22428 41188 22434 41200
rect 23201 41191 23259 41197
rect 23201 41188 23213 41191
rect 22428 41160 23213 41188
rect 22428 41148 22434 41160
rect 23201 41157 23213 41160
rect 23247 41157 23259 41191
rect 24486 41188 24492 41200
rect 24426 41160 24492 41188
rect 23201 41151 23259 41157
rect 24486 41148 24492 41160
rect 24544 41148 24550 41200
rect 25314 41080 25320 41132
rect 25372 41080 25378 41132
rect 22830 41012 22836 41064
rect 22888 41052 22894 41064
rect 22925 41055 22983 41061
rect 22925 41052 22937 41055
rect 22888 41024 22937 41052
rect 22888 41012 22894 41024
rect 22925 41021 22937 41024
rect 22971 41021 22983 41055
rect 23658 41052 23664 41064
rect 22925 41015 22983 41021
rect 23032 41024 23664 41052
rect 23032 40984 23060 41024
rect 23658 41012 23664 41024
rect 23716 41012 23722 41064
rect 22066 40956 23060 40984
rect 15749 40919 15807 40925
rect 15749 40885 15761 40919
rect 15795 40916 15807 40919
rect 18414 40916 18420 40928
rect 15795 40888 18420 40916
rect 15795 40885 15807 40888
rect 15749 40879 15807 40885
rect 18414 40876 18420 40888
rect 18472 40876 18478 40928
rect 18601 40919 18659 40925
rect 18601 40885 18613 40919
rect 18647 40916 18659 40919
rect 18690 40916 18696 40928
rect 18647 40888 18696 40916
rect 18647 40885 18659 40888
rect 18601 40879 18659 40885
rect 18690 40876 18696 40888
rect 18748 40876 18754 40928
rect 18874 40876 18880 40928
rect 18932 40916 18938 40928
rect 19061 40919 19119 40925
rect 19061 40916 19073 40919
rect 18932 40888 19073 40916
rect 18932 40876 18938 40888
rect 19061 40885 19073 40888
rect 19107 40885 19119 40919
rect 19061 40879 19119 40885
rect 19426 40876 19432 40928
rect 19484 40876 19490 40928
rect 20717 40919 20775 40925
rect 20717 40885 20729 40919
rect 20763 40916 20775 40919
rect 20898 40916 20904 40928
rect 20763 40888 20904 40916
rect 20763 40885 20775 40888
rect 20717 40879 20775 40885
rect 20898 40876 20904 40888
rect 20956 40876 20962 40928
rect 21082 40876 21088 40928
rect 21140 40916 21146 40928
rect 25133 40919 25191 40925
rect 25133 40916 25145 40919
rect 21140 40888 25145 40916
rect 21140 40876 21146 40888
rect 25133 40885 25145 40888
rect 25179 40885 25191 40919
rect 25133 40879 25191 40885
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 8294 40672 8300 40724
rect 8352 40672 8358 40724
rect 9490 40672 9496 40724
rect 9548 40712 9554 40724
rect 9548 40684 11928 40712
rect 9548 40672 9554 40684
rect 9217 40647 9275 40653
rect 9217 40613 9229 40647
rect 9263 40644 9275 40647
rect 10226 40644 10232 40656
rect 9263 40616 10232 40644
rect 9263 40613 9275 40616
rect 9217 40607 9275 40613
rect 10226 40604 10232 40616
rect 10284 40604 10290 40656
rect 10689 40647 10747 40653
rect 10689 40613 10701 40647
rect 10735 40644 10747 40647
rect 11330 40644 11336 40656
rect 10735 40616 11336 40644
rect 10735 40613 10747 40616
rect 10689 40607 10747 40613
rect 11330 40604 11336 40616
rect 11388 40604 11394 40656
rect 6457 40579 6515 40585
rect 6457 40545 6469 40579
rect 6503 40576 6515 40579
rect 6546 40576 6552 40588
rect 6503 40548 6552 40576
rect 6503 40545 6515 40548
rect 6457 40539 6515 40545
rect 6546 40536 6552 40548
rect 6604 40576 6610 40588
rect 6604 40548 8432 40576
rect 6604 40536 6610 40548
rect 6178 40468 6184 40520
rect 6236 40468 6242 40520
rect 8404 40508 8432 40548
rect 9398 40536 9404 40588
rect 9456 40576 9462 40588
rect 9582 40576 9588 40588
rect 9456 40548 9588 40576
rect 9456 40536 9462 40548
rect 9582 40536 9588 40548
rect 9640 40536 9646 40588
rect 9674 40536 9680 40588
rect 9732 40576 9738 40588
rect 11900 40585 11928 40684
rect 14826 40672 14832 40724
rect 14884 40712 14890 40724
rect 18598 40712 18604 40724
rect 14884 40684 18604 40712
rect 14884 40672 14890 40684
rect 18598 40672 18604 40684
rect 18656 40672 18662 40724
rect 20901 40715 20959 40721
rect 20901 40681 20913 40715
rect 20947 40712 20959 40715
rect 22186 40712 22192 40724
rect 20947 40684 22192 40712
rect 20947 40681 20959 40684
rect 20901 40675 20959 40681
rect 22186 40672 22192 40684
rect 22244 40672 22250 40724
rect 24854 40712 24860 40724
rect 22296 40684 24860 40712
rect 12621 40647 12679 40653
rect 12621 40613 12633 40647
rect 12667 40644 12679 40647
rect 13354 40644 13360 40656
rect 12667 40616 13360 40644
rect 12667 40613 12679 40616
rect 12621 40607 12679 40613
rect 13354 40604 13360 40616
rect 13412 40604 13418 40656
rect 13725 40647 13783 40653
rect 13725 40613 13737 40647
rect 13771 40644 13783 40647
rect 15838 40644 15844 40656
rect 13771 40616 15844 40644
rect 13771 40613 13783 40616
rect 13725 40607 13783 40613
rect 9769 40579 9827 40585
rect 9769 40576 9781 40579
rect 9732 40548 9781 40576
rect 9732 40536 9738 40548
rect 9769 40545 9781 40548
rect 9815 40545 9827 40579
rect 9769 40539 9827 40545
rect 11885 40579 11943 40585
rect 11885 40545 11897 40579
rect 11931 40545 11943 40579
rect 11885 40539 11943 40545
rect 11977 40579 12035 40585
rect 11977 40545 11989 40579
rect 12023 40545 12035 40579
rect 11977 40539 12035 40545
rect 13265 40579 13323 40585
rect 13265 40545 13277 40579
rect 13311 40576 13323 40579
rect 13630 40576 13636 40588
rect 13311 40548 13636 40576
rect 13311 40545 13323 40548
rect 13265 40539 13323 40545
rect 11992 40508 12020 40539
rect 13630 40536 13636 40548
rect 13688 40536 13694 40588
rect 8404 40480 12020 40508
rect 12710 40468 12716 40520
rect 12768 40508 12774 40520
rect 12989 40511 13047 40517
rect 12989 40508 13001 40511
rect 12768 40480 13001 40508
rect 12768 40468 12774 40480
rect 12989 40477 13001 40480
rect 13035 40477 13047 40511
rect 12989 40471 13047 40477
rect 13081 40511 13139 40517
rect 13081 40477 13093 40511
rect 13127 40508 13139 40511
rect 13740 40508 13768 40607
rect 15838 40604 15844 40616
rect 15896 40604 15902 40656
rect 16942 40604 16948 40656
rect 17000 40644 17006 40656
rect 17000 40616 17264 40644
rect 17000 40604 17006 40616
rect 15470 40536 15476 40588
rect 15528 40576 15534 40588
rect 15746 40576 15752 40588
rect 15528 40548 15752 40576
rect 15528 40536 15534 40548
rect 15746 40536 15752 40548
rect 15804 40536 15810 40588
rect 17034 40536 17040 40588
rect 17092 40576 17098 40588
rect 17236 40585 17264 40616
rect 19794 40604 19800 40656
rect 19852 40644 19858 40656
rect 20530 40644 20536 40656
rect 19852 40616 20536 40644
rect 19852 40604 19858 40616
rect 20530 40604 20536 40616
rect 20588 40604 20594 40656
rect 22002 40604 22008 40656
rect 22060 40644 22066 40656
rect 22097 40647 22155 40653
rect 22097 40644 22109 40647
rect 22060 40616 22109 40644
rect 22060 40604 22066 40616
rect 22097 40613 22109 40616
rect 22143 40644 22155 40647
rect 22296 40644 22324 40684
rect 24854 40672 24860 40684
rect 24912 40672 24918 40724
rect 22143 40616 22324 40644
rect 22143 40613 22155 40616
rect 22097 40607 22155 40613
rect 22462 40604 22468 40656
rect 22520 40604 22526 40656
rect 22738 40604 22744 40656
rect 22796 40644 22802 40656
rect 22796 40616 23060 40644
rect 22796 40604 22802 40616
rect 17129 40579 17187 40585
rect 17129 40576 17141 40579
rect 17092 40548 17141 40576
rect 17092 40536 17098 40548
rect 17129 40545 17141 40548
rect 17175 40545 17187 40579
rect 17129 40539 17187 40545
rect 17221 40579 17279 40585
rect 17221 40545 17233 40579
rect 17267 40545 17279 40579
rect 17221 40539 17279 40545
rect 18874 40536 18880 40588
rect 18932 40576 18938 40588
rect 21358 40576 21364 40588
rect 18932 40548 21364 40576
rect 18932 40536 18938 40548
rect 21358 40536 21364 40548
rect 21416 40536 21422 40588
rect 21450 40536 21456 40588
rect 21508 40536 21514 40588
rect 23032 40585 23060 40616
rect 23106 40604 23112 40656
rect 23164 40644 23170 40656
rect 23842 40644 23848 40656
rect 23164 40616 23848 40644
rect 23164 40604 23170 40616
rect 23842 40604 23848 40616
rect 23900 40604 23906 40656
rect 21545 40579 21603 40585
rect 21545 40545 21557 40579
rect 21591 40545 21603 40579
rect 21545 40539 21603 40545
rect 23017 40579 23075 40585
rect 23017 40545 23029 40579
rect 23063 40545 23075 40579
rect 25406 40576 25412 40588
rect 23017 40539 23075 40545
rect 23308 40548 25412 40576
rect 13127 40480 13768 40508
rect 15565 40511 15623 40517
rect 13127 40477 13139 40480
rect 13081 40471 13139 40477
rect 15565 40477 15577 40511
rect 15611 40508 15623 40511
rect 21468 40508 21496 40536
rect 15611 40480 21496 40508
rect 15611 40477 15623 40480
rect 15565 40471 15623 40477
rect 8294 40440 8300 40452
rect 7682 40412 8300 40440
rect 8294 40400 8300 40412
rect 8352 40440 8358 40452
rect 9214 40440 9220 40452
rect 8352 40412 9220 40440
rect 8352 40400 8358 40412
rect 9214 40400 9220 40412
rect 9272 40400 9278 40452
rect 9582 40400 9588 40452
rect 9640 40400 9646 40452
rect 11333 40443 11391 40449
rect 11333 40409 11345 40443
rect 11379 40440 11391 40443
rect 11793 40443 11851 40449
rect 11793 40440 11805 40443
rect 11379 40412 11805 40440
rect 11379 40409 11391 40412
rect 11333 40403 11391 40409
rect 11793 40409 11805 40412
rect 11839 40440 11851 40443
rect 11839 40412 12020 40440
rect 11839 40409 11851 40412
rect 11793 40403 11851 40409
rect 7098 40332 7104 40384
rect 7156 40372 7162 40384
rect 7742 40372 7748 40384
rect 7156 40344 7748 40372
rect 7156 40332 7162 40344
rect 7742 40332 7748 40344
rect 7800 40372 7806 40384
rect 7929 40375 7987 40381
rect 7929 40372 7941 40375
rect 7800 40344 7941 40372
rect 7800 40332 7806 40344
rect 7929 40341 7941 40344
rect 7975 40341 7987 40375
rect 7929 40335 7987 40341
rect 9398 40332 9404 40384
rect 9456 40372 9462 40384
rect 9677 40375 9735 40381
rect 9677 40372 9689 40375
rect 9456 40344 9689 40372
rect 9456 40332 9462 40344
rect 9677 40341 9689 40344
rect 9723 40341 9735 40375
rect 9677 40335 9735 40341
rect 11422 40332 11428 40384
rect 11480 40332 11486 40384
rect 11992 40372 12020 40412
rect 12434 40400 12440 40452
rect 12492 40440 12498 40452
rect 15657 40443 15715 40449
rect 15657 40440 15669 40443
rect 12492 40412 15669 40440
rect 12492 40400 12498 40412
rect 15657 40409 15669 40412
rect 15703 40409 15715 40443
rect 17678 40440 17684 40452
rect 15657 40403 15715 40409
rect 16684 40412 17684 40440
rect 14826 40372 14832 40384
rect 11992 40344 14832 40372
rect 14826 40332 14832 40344
rect 14884 40332 14890 40384
rect 15194 40332 15200 40384
rect 15252 40332 15258 40384
rect 16684 40381 16712 40412
rect 17678 40400 17684 40412
rect 17736 40400 17742 40452
rect 20162 40400 20168 40452
rect 20220 40440 20226 40452
rect 20349 40443 20407 40449
rect 20349 40440 20361 40443
rect 20220 40412 20361 40440
rect 20220 40400 20226 40412
rect 20349 40409 20361 40412
rect 20395 40440 20407 40443
rect 20395 40412 21404 40440
rect 20395 40409 20407 40412
rect 20349 40403 20407 40409
rect 16669 40375 16727 40381
rect 16669 40341 16681 40375
rect 16715 40341 16727 40375
rect 16669 40335 16727 40341
rect 17034 40332 17040 40384
rect 17092 40332 17098 40384
rect 17310 40332 17316 40384
rect 17368 40372 17374 40384
rect 18874 40372 18880 40384
rect 17368 40344 18880 40372
rect 17368 40332 17374 40344
rect 18874 40332 18880 40344
rect 18932 40332 18938 40384
rect 20990 40332 20996 40384
rect 21048 40372 21054 40384
rect 21269 40375 21327 40381
rect 21269 40372 21281 40375
rect 21048 40344 21281 40372
rect 21048 40332 21054 40344
rect 21269 40341 21281 40344
rect 21315 40341 21327 40375
rect 21376 40372 21404 40412
rect 21450 40400 21456 40452
rect 21508 40440 21514 40452
rect 21560 40440 21588 40539
rect 23308 40520 23336 40548
rect 25406 40536 25412 40548
rect 25464 40536 25470 40588
rect 22554 40468 22560 40520
rect 22612 40508 22618 40520
rect 22833 40511 22891 40517
rect 22833 40508 22845 40511
rect 22612 40480 22845 40508
rect 22612 40468 22618 40480
rect 22833 40477 22845 40480
rect 22879 40477 22891 40511
rect 22833 40471 22891 40477
rect 22922 40468 22928 40520
rect 22980 40468 22986 40520
rect 23290 40468 23296 40520
rect 23348 40468 23354 40520
rect 24026 40468 24032 40520
rect 24084 40508 24090 40520
rect 24397 40511 24455 40517
rect 24397 40508 24409 40511
rect 24084 40480 24409 40508
rect 24084 40468 24090 40480
rect 24397 40477 24409 40480
rect 24443 40508 24455 40511
rect 24486 40508 24492 40520
rect 24443 40480 24492 40508
rect 24443 40477 24455 40480
rect 24397 40471 24455 40477
rect 24486 40468 24492 40480
rect 24544 40468 24550 40520
rect 24673 40511 24731 40517
rect 24673 40477 24685 40511
rect 24719 40508 24731 40511
rect 24762 40508 24768 40520
rect 24719 40480 24768 40508
rect 24719 40477 24731 40480
rect 24673 40471 24731 40477
rect 24762 40468 24768 40480
rect 24820 40508 24826 40520
rect 25317 40511 25375 40517
rect 25317 40508 25329 40511
rect 24820 40480 25329 40508
rect 24820 40468 24826 40480
rect 25317 40477 25329 40480
rect 25363 40477 25375 40511
rect 25317 40471 25375 40477
rect 21508 40412 21588 40440
rect 21508 40400 21514 40412
rect 21634 40400 21640 40452
rect 21692 40440 21698 40452
rect 22005 40443 22063 40449
rect 22005 40440 22017 40443
rect 21692 40412 22017 40440
rect 21692 40400 21698 40412
rect 22005 40409 22017 40412
rect 22051 40440 22063 40443
rect 22186 40440 22192 40452
rect 22051 40412 22192 40440
rect 22051 40409 22063 40412
rect 22005 40403 22063 40409
rect 22186 40400 22192 40412
rect 22244 40440 22250 40452
rect 23566 40440 23572 40452
rect 22244 40412 23572 40440
rect 22244 40400 22250 40412
rect 23566 40400 23572 40412
rect 23624 40400 23630 40452
rect 24857 40443 24915 40449
rect 24857 40409 24869 40443
rect 24903 40440 24915 40443
rect 24903 40412 25360 40440
rect 24903 40409 24915 40412
rect 24857 40403 24915 40409
rect 25332 40384 25360 40412
rect 23290 40372 23296 40384
rect 21376 40344 23296 40372
rect 21269 40335 21327 40341
rect 23290 40332 23296 40344
rect 23348 40332 23354 40384
rect 24026 40332 24032 40384
rect 24084 40332 24090 40384
rect 24210 40332 24216 40384
rect 24268 40332 24274 40384
rect 24578 40332 24584 40384
rect 24636 40372 24642 40384
rect 25133 40375 25191 40381
rect 25133 40372 25145 40375
rect 24636 40344 25145 40372
rect 24636 40332 24642 40344
rect 25133 40341 25145 40344
rect 25179 40341 25191 40375
rect 25133 40335 25191 40341
rect 25314 40332 25320 40384
rect 25372 40332 25378 40384
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 7285 40171 7343 40177
rect 7285 40137 7297 40171
rect 7331 40168 7343 40171
rect 8662 40168 8668 40180
rect 7331 40140 8668 40168
rect 7331 40137 7343 40140
rect 7285 40131 7343 40137
rect 8662 40128 8668 40140
rect 8720 40128 8726 40180
rect 9582 40128 9588 40180
rect 9640 40168 9646 40180
rect 9640 40140 10548 40168
rect 9640 40128 9646 40140
rect 7653 40103 7711 40109
rect 7653 40069 7665 40103
rect 7699 40100 7711 40103
rect 8754 40100 8760 40112
rect 7699 40072 8760 40100
rect 7699 40069 7711 40072
rect 7653 40063 7711 40069
rect 8754 40060 8760 40072
rect 8812 40060 8818 40112
rect 9214 40060 9220 40112
rect 9272 40060 9278 40112
rect 10520 40109 10548 40140
rect 14292 40140 14504 40168
rect 10505 40103 10563 40109
rect 10505 40069 10517 40103
rect 10551 40069 10563 40103
rect 10505 40063 10563 40069
rect 10962 40060 10968 40112
rect 11020 40060 11026 40112
rect 8478 39992 8484 40044
rect 8536 39992 8542 40044
rect 10980 40032 11008 40060
rect 14292 40044 14320 40140
rect 14476 40100 14504 40140
rect 15010 40128 15016 40180
rect 15068 40128 15074 40180
rect 15102 40128 15108 40180
rect 15160 40168 15166 40180
rect 15565 40171 15623 40177
rect 15565 40168 15577 40171
rect 15160 40140 15577 40168
rect 15160 40128 15166 40140
rect 15565 40137 15577 40140
rect 15611 40137 15623 40171
rect 15565 40131 15623 40137
rect 19797 40171 19855 40177
rect 19797 40137 19809 40171
rect 19843 40168 19855 40171
rect 20622 40168 20628 40180
rect 19843 40140 20628 40168
rect 19843 40137 19855 40140
rect 19797 40131 19855 40137
rect 20622 40128 20628 40140
rect 20680 40128 20686 40180
rect 21450 40128 21456 40180
rect 21508 40168 21514 40180
rect 22094 40168 22100 40180
rect 21508 40140 22100 40168
rect 21508 40128 21514 40140
rect 22094 40128 22100 40140
rect 22152 40168 22158 40180
rect 25225 40171 25283 40177
rect 25225 40168 25237 40171
rect 22152 40140 25237 40168
rect 22152 40128 22158 40140
rect 25225 40137 25237 40140
rect 25271 40137 25283 40171
rect 25225 40131 25283 40137
rect 15028 40100 15056 40128
rect 14398 40072 15056 40100
rect 15838 40060 15844 40112
rect 15896 40100 15902 40112
rect 15933 40103 15991 40109
rect 15933 40100 15945 40103
rect 15896 40072 15945 40100
rect 15896 40060 15902 40072
rect 15933 40069 15945 40072
rect 15979 40069 15991 40103
rect 15933 40063 15991 40069
rect 16942 40060 16948 40112
rect 17000 40100 17006 40112
rect 18601 40103 18659 40109
rect 18601 40100 18613 40103
rect 17000 40072 18613 40100
rect 17000 40060 17006 40072
rect 18601 40069 18613 40072
rect 18647 40069 18659 40103
rect 18601 40063 18659 40069
rect 20165 40103 20223 40109
rect 20165 40069 20177 40103
rect 20211 40069 20223 40103
rect 20165 40063 20223 40069
rect 12710 40032 12716 40044
rect 10980 40004 12716 40032
rect 12710 39992 12716 40004
rect 12768 39992 12774 40044
rect 12802 39992 12808 40044
rect 12860 40032 12866 40044
rect 12897 40035 12955 40041
rect 12897 40032 12909 40035
rect 12860 40004 12909 40032
rect 12860 39992 12866 40004
rect 12897 40001 12909 40004
rect 12943 40001 12955 40035
rect 12897 39995 12955 40001
rect 14274 39992 14280 40044
rect 14332 39992 14338 40044
rect 17126 39992 17132 40044
rect 17184 40032 17190 40044
rect 20180 40032 20208 40063
rect 20990 40060 20996 40112
rect 21048 40100 21054 40112
rect 22002 40100 22008 40112
rect 21048 40072 22008 40100
rect 21048 40060 21054 40072
rect 22002 40060 22008 40072
rect 22060 40100 22066 40112
rect 22281 40103 22339 40109
rect 22281 40100 22293 40103
rect 22060 40072 22293 40100
rect 22060 40060 22066 40072
rect 22281 40069 22293 40072
rect 22327 40069 22339 40103
rect 22281 40063 22339 40069
rect 22830 40060 22836 40112
rect 22888 40100 22894 40112
rect 22888 40072 23428 40100
rect 22888 40060 22894 40072
rect 21085 40035 21143 40041
rect 21085 40032 21097 40035
rect 17184 40004 21097 40032
rect 17184 39992 17190 40004
rect 21085 40001 21097 40004
rect 21131 40032 21143 40035
rect 23400 40032 23428 40072
rect 24026 40060 24032 40112
rect 24084 40100 24090 40112
rect 24084 40072 24242 40100
rect 24084 40060 24090 40072
rect 23477 40035 23535 40041
rect 23477 40032 23489 40035
rect 21131 40004 22094 40032
rect 23400 40004 23489 40032
rect 21131 40001 21143 40004
rect 21085 39995 21143 40001
rect 7742 39924 7748 39976
rect 7800 39924 7806 39976
rect 7834 39924 7840 39976
rect 7892 39924 7898 39976
rect 8757 39967 8815 39973
rect 8757 39933 8769 39967
rect 8803 39964 8815 39967
rect 9950 39964 9956 39976
rect 8803 39936 9956 39964
rect 8803 39933 8815 39936
rect 8757 39927 8815 39933
rect 9950 39924 9956 39936
rect 10008 39924 10014 39976
rect 10962 39924 10968 39976
rect 11020 39924 11026 39976
rect 13173 39967 13231 39973
rect 13173 39933 13185 39967
rect 13219 39964 13231 39967
rect 15562 39964 15568 39976
rect 13219 39936 15568 39964
rect 13219 39933 13231 39936
rect 13173 39927 13231 39933
rect 15562 39924 15568 39936
rect 15620 39924 15626 39976
rect 16022 39924 16028 39976
rect 16080 39924 16086 39976
rect 16117 39967 16175 39973
rect 16117 39933 16129 39967
rect 16163 39933 16175 39967
rect 16117 39927 16175 39933
rect 16132 39896 16160 39927
rect 18506 39924 18512 39976
rect 18564 39964 18570 39976
rect 18693 39967 18751 39973
rect 18693 39964 18705 39967
rect 18564 39936 18705 39964
rect 18564 39924 18570 39936
rect 18693 39933 18705 39936
rect 18739 39933 18751 39967
rect 18693 39927 18751 39933
rect 18782 39924 18788 39976
rect 18840 39924 18846 39976
rect 19518 39924 19524 39976
rect 19576 39964 19582 39976
rect 19794 39964 19800 39976
rect 19576 39936 19800 39964
rect 19576 39924 19582 39936
rect 19794 39924 19800 39936
rect 19852 39964 19858 39976
rect 20257 39967 20315 39973
rect 20257 39964 20269 39967
rect 19852 39936 20269 39964
rect 19852 39924 19858 39936
rect 20257 39933 20269 39936
rect 20303 39933 20315 39967
rect 20257 39927 20315 39933
rect 14292 39868 16160 39896
rect 20272 39896 20300 39927
rect 20346 39924 20352 39976
rect 20404 39924 20410 39976
rect 22066 39964 22094 40004
rect 23477 40001 23489 40004
rect 23523 40001 23535 40035
rect 23477 39995 23535 40001
rect 22554 39964 22560 39976
rect 22066 39936 22560 39964
rect 22554 39924 22560 39936
rect 22612 39924 22618 39976
rect 23753 39967 23811 39973
rect 23753 39933 23765 39967
rect 23799 39964 23811 39967
rect 24486 39964 24492 39976
rect 23799 39936 24492 39964
rect 23799 39933 23811 39936
rect 23753 39927 23811 39933
rect 24486 39924 24492 39936
rect 24544 39924 24550 39976
rect 20809 39899 20867 39905
rect 20809 39896 20821 39899
rect 20272 39868 20821 39896
rect 10778 39788 10784 39840
rect 10836 39828 10842 39840
rect 14292 39828 14320 39868
rect 20809 39865 20821 39868
rect 20855 39896 20867 39899
rect 20855 39868 22094 39896
rect 20855 39865 20867 39868
rect 20809 39859 20867 39865
rect 10836 39800 14320 39828
rect 10836 39788 10842 39800
rect 14550 39788 14556 39840
rect 14608 39828 14614 39840
rect 14645 39831 14703 39837
rect 14645 39828 14657 39831
rect 14608 39800 14657 39828
rect 14608 39788 14614 39800
rect 14645 39797 14657 39800
rect 14691 39828 14703 39831
rect 14734 39828 14740 39840
rect 14691 39800 14740 39828
rect 14691 39797 14703 39800
rect 14645 39791 14703 39797
rect 14734 39788 14740 39800
rect 14792 39788 14798 39840
rect 18233 39831 18291 39837
rect 18233 39797 18245 39831
rect 18279 39828 18291 39831
rect 19242 39828 19248 39840
rect 18279 39800 19248 39828
rect 18279 39797 18291 39800
rect 18233 39791 18291 39797
rect 19242 39788 19248 39800
rect 19300 39788 19306 39840
rect 22066 39828 22094 39868
rect 23750 39828 23756 39840
rect 22066 39800 23756 39828
rect 23750 39788 23756 39800
rect 23808 39788 23814 39840
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 6546 39584 6552 39636
rect 6604 39624 6610 39636
rect 6641 39627 6699 39633
rect 6641 39624 6653 39627
rect 6604 39596 6653 39624
rect 6604 39584 6610 39596
rect 6641 39593 6653 39596
rect 6687 39593 6699 39627
rect 6641 39587 6699 39593
rect 7742 39584 7748 39636
rect 7800 39624 7806 39636
rect 9769 39627 9827 39633
rect 9769 39624 9781 39627
rect 7800 39596 9781 39624
rect 7800 39584 7806 39596
rect 9769 39593 9781 39596
rect 9815 39593 9827 39627
rect 9769 39587 9827 39593
rect 10870 39584 10876 39636
rect 10928 39624 10934 39636
rect 12894 39624 12900 39636
rect 10928 39596 12900 39624
rect 10928 39584 10934 39596
rect 12894 39584 12900 39596
rect 12952 39584 12958 39636
rect 13078 39584 13084 39636
rect 13136 39624 13142 39636
rect 14274 39624 14280 39636
rect 13136 39596 14280 39624
rect 13136 39584 13142 39596
rect 14274 39584 14280 39596
rect 14332 39584 14338 39636
rect 14369 39627 14427 39633
rect 14369 39593 14381 39627
rect 14415 39624 14427 39627
rect 17034 39624 17040 39636
rect 14415 39596 17040 39624
rect 14415 39593 14427 39596
rect 14369 39587 14427 39593
rect 17034 39584 17040 39596
rect 17092 39584 17098 39636
rect 21269 39627 21327 39633
rect 21269 39593 21281 39627
rect 21315 39624 21327 39627
rect 22278 39624 22284 39636
rect 21315 39596 22284 39624
rect 21315 39593 21327 39596
rect 21269 39587 21327 39593
rect 22278 39584 22284 39596
rect 22336 39584 22342 39636
rect 25130 39624 25136 39636
rect 22388 39596 25136 39624
rect 6730 39516 6736 39568
rect 6788 39556 6794 39568
rect 8570 39556 8576 39568
rect 6788 39528 8576 39556
rect 6788 39516 6794 39528
rect 8570 39516 8576 39528
rect 8628 39516 8634 39568
rect 12710 39516 12716 39568
rect 12768 39556 12774 39568
rect 15565 39559 15623 39565
rect 15565 39556 15577 39559
rect 12768 39528 15577 39556
rect 12768 39516 12774 39528
rect 15565 39525 15577 39528
rect 15611 39525 15623 39559
rect 15565 39519 15623 39525
rect 16022 39516 16028 39568
rect 16080 39556 16086 39568
rect 22388 39556 22416 39596
rect 25130 39584 25136 39596
rect 25188 39584 25194 39636
rect 16080 39528 22416 39556
rect 22649 39559 22707 39565
rect 16080 39516 16086 39528
rect 22649 39525 22661 39559
rect 22695 39556 22707 39559
rect 22695 39528 24992 39556
rect 22695 39525 22707 39528
rect 22649 39519 22707 39525
rect 4893 39491 4951 39497
rect 4893 39457 4905 39491
rect 4939 39488 4951 39491
rect 6178 39488 6184 39500
rect 4939 39460 6184 39488
rect 4939 39457 4951 39460
rect 4893 39451 4951 39457
rect 6178 39448 6184 39460
rect 6236 39448 6242 39500
rect 10226 39448 10232 39500
rect 10284 39448 10290 39500
rect 10321 39491 10379 39497
rect 10321 39457 10333 39491
rect 10367 39457 10379 39491
rect 10321 39451 10379 39457
rect 10965 39491 11023 39497
rect 10965 39457 10977 39491
rect 11011 39488 11023 39491
rect 12618 39488 12624 39500
rect 11011 39460 12624 39488
rect 11011 39457 11023 39460
rect 10965 39451 11023 39457
rect 8570 39380 8576 39432
rect 8628 39420 8634 39432
rect 10336 39420 10364 39451
rect 12618 39448 12624 39460
rect 12676 39488 12682 39500
rect 12802 39488 12808 39500
rect 12676 39460 12808 39488
rect 12676 39448 12682 39460
rect 12802 39448 12808 39460
rect 12860 39448 12866 39500
rect 15013 39491 15071 39497
rect 15013 39457 15025 39491
rect 15059 39488 15071 39491
rect 15654 39488 15660 39500
rect 15059 39460 15660 39488
rect 15059 39457 15071 39460
rect 15013 39451 15071 39457
rect 15654 39448 15660 39460
rect 15712 39448 15718 39500
rect 16209 39491 16267 39497
rect 16209 39457 16221 39491
rect 16255 39488 16267 39491
rect 17862 39488 17868 39500
rect 16255 39460 17868 39488
rect 16255 39457 16267 39460
rect 16209 39451 16267 39457
rect 17862 39448 17868 39460
rect 17920 39448 17926 39500
rect 18598 39448 18604 39500
rect 18656 39488 18662 39500
rect 18782 39488 18788 39500
rect 18656 39460 18788 39488
rect 18656 39448 18662 39460
rect 18782 39448 18788 39460
rect 18840 39448 18846 39500
rect 19426 39448 19432 39500
rect 19484 39488 19490 39500
rect 19889 39491 19947 39497
rect 19889 39488 19901 39491
rect 19484 39460 19901 39488
rect 19484 39448 19490 39460
rect 19889 39457 19901 39460
rect 19935 39457 19947 39491
rect 19889 39451 19947 39457
rect 20070 39448 20076 39500
rect 20128 39448 20134 39500
rect 21358 39448 21364 39500
rect 21416 39488 21422 39500
rect 21821 39491 21879 39497
rect 21821 39488 21833 39491
rect 21416 39460 21833 39488
rect 21416 39448 21422 39460
rect 21821 39457 21833 39460
rect 21867 39488 21879 39491
rect 22370 39488 22376 39500
rect 21867 39460 22376 39488
rect 21867 39457 21879 39460
rect 21821 39451 21879 39457
rect 22370 39448 22376 39460
rect 22428 39448 22434 39500
rect 22554 39448 22560 39500
rect 22612 39488 22618 39500
rect 23293 39491 23351 39497
rect 22612 39460 23244 39488
rect 22612 39448 22618 39460
rect 8628 39392 10364 39420
rect 8628 39380 8634 39392
rect 12250 39380 12256 39432
rect 12308 39420 12314 39432
rect 13078 39420 13084 39432
rect 12308 39392 13084 39420
rect 12308 39380 12314 39392
rect 13078 39380 13084 39392
rect 13136 39380 13142 39432
rect 18432 39392 19932 39420
rect 5169 39355 5227 39361
rect 5169 39321 5181 39355
rect 5215 39321 5227 39355
rect 11241 39355 11299 39361
rect 6394 39324 7052 39352
rect 5169 39315 5227 39321
rect 5184 39284 5212 39315
rect 5810 39284 5816 39296
rect 5184 39256 5816 39284
rect 5810 39244 5816 39256
rect 5868 39244 5874 39296
rect 7024 39293 7052 39324
rect 11241 39321 11253 39355
rect 11287 39352 11299 39355
rect 11514 39352 11520 39364
rect 11287 39324 11520 39352
rect 11287 39321 11299 39324
rect 11241 39315 11299 39321
rect 11514 39312 11520 39324
rect 11572 39312 11578 39364
rect 14829 39355 14887 39361
rect 14829 39352 14841 39355
rect 13832 39324 14841 39352
rect 13832 39296 13860 39324
rect 14829 39321 14841 39324
rect 14875 39321 14887 39355
rect 14829 39315 14887 39321
rect 15010 39312 15016 39364
rect 15068 39352 15074 39364
rect 18432 39352 18460 39392
rect 15068 39324 18460 39352
rect 15068 39312 15074 39324
rect 18598 39312 18604 39364
rect 18656 39352 18662 39364
rect 19797 39355 19855 39361
rect 19797 39352 19809 39355
rect 18656 39324 19809 39352
rect 18656 39312 18662 39324
rect 19797 39321 19809 39324
rect 19843 39321 19855 39355
rect 19797 39315 19855 39321
rect 7009 39287 7067 39293
rect 7009 39253 7021 39287
rect 7055 39284 7067 39287
rect 7374 39284 7380 39296
rect 7055 39256 7380 39284
rect 7055 39253 7067 39256
rect 7009 39247 7067 39253
rect 7374 39244 7380 39256
rect 7432 39244 7438 39296
rect 8294 39244 8300 39296
rect 8352 39284 8358 39296
rect 9125 39287 9183 39293
rect 9125 39284 9137 39287
rect 8352 39256 9137 39284
rect 8352 39244 8358 39256
rect 9125 39253 9137 39256
rect 9171 39253 9183 39287
rect 9125 39247 9183 39253
rect 10137 39287 10195 39293
rect 10137 39253 10149 39287
rect 10183 39284 10195 39287
rect 12250 39284 12256 39296
rect 10183 39256 12256 39284
rect 10183 39253 10195 39256
rect 10137 39247 10195 39253
rect 12250 39244 12256 39256
rect 12308 39244 12314 39296
rect 12710 39244 12716 39296
rect 12768 39244 12774 39296
rect 13814 39244 13820 39296
rect 13872 39244 13878 39296
rect 14734 39244 14740 39296
rect 14792 39244 14798 39296
rect 15378 39244 15384 39296
rect 15436 39284 15442 39296
rect 15933 39287 15991 39293
rect 15933 39284 15945 39287
rect 15436 39256 15945 39284
rect 15436 39244 15442 39256
rect 15933 39253 15945 39256
rect 15979 39253 15991 39287
rect 15933 39247 15991 39253
rect 16022 39244 16028 39296
rect 16080 39244 16086 39296
rect 18414 39244 18420 39296
rect 18472 39284 18478 39296
rect 18785 39287 18843 39293
rect 18785 39284 18797 39287
rect 18472 39256 18797 39284
rect 18472 39244 18478 39256
rect 18785 39253 18797 39256
rect 18831 39253 18843 39287
rect 18785 39247 18843 39253
rect 19429 39287 19487 39293
rect 19429 39253 19441 39287
rect 19475 39284 19487 39287
rect 19518 39284 19524 39296
rect 19475 39256 19524 39284
rect 19475 39253 19487 39256
rect 19429 39247 19487 39253
rect 19518 39244 19524 39256
rect 19576 39244 19582 39296
rect 19904 39284 19932 39392
rect 20346 39380 20352 39432
rect 20404 39420 20410 39432
rect 23109 39423 23167 39429
rect 23109 39420 23121 39423
rect 20404 39392 23121 39420
rect 20404 39380 20410 39392
rect 23109 39389 23121 39392
rect 23155 39389 23167 39423
rect 23216 39420 23244 39460
rect 23293 39457 23305 39491
rect 23339 39488 23351 39491
rect 23474 39488 23480 39500
rect 23339 39460 23480 39488
rect 23339 39457 23351 39460
rect 23293 39451 23351 39457
rect 23474 39448 23480 39460
rect 23532 39448 23538 39500
rect 23566 39420 23572 39432
rect 23216 39392 23572 39420
rect 23109 39383 23167 39389
rect 23566 39380 23572 39392
rect 23624 39380 23630 39432
rect 24964 39429 24992 39528
rect 25038 39448 25044 39500
rect 25096 39448 25102 39500
rect 25225 39491 25283 39497
rect 25225 39457 25237 39491
rect 25271 39488 25283 39491
rect 25498 39488 25504 39500
rect 25271 39460 25504 39488
rect 25271 39457 25283 39460
rect 25225 39451 25283 39457
rect 25498 39448 25504 39460
rect 25556 39448 25562 39500
rect 24949 39423 25007 39429
rect 24949 39389 24961 39423
rect 24995 39389 25007 39423
rect 24949 39383 25007 39389
rect 20438 39312 20444 39364
rect 20496 39312 20502 39364
rect 21729 39355 21787 39361
rect 21729 39321 21741 39355
rect 21775 39352 21787 39355
rect 22186 39352 22192 39364
rect 21775 39324 22192 39352
rect 21775 39321 21787 39324
rect 21729 39315 21787 39321
rect 22186 39312 22192 39324
rect 22244 39352 22250 39364
rect 22281 39355 22339 39361
rect 22281 39352 22293 39355
rect 22244 39324 22293 39352
rect 22244 39312 22250 39324
rect 22281 39321 22293 39324
rect 22327 39321 22339 39355
rect 22281 39315 22339 39321
rect 23017 39355 23075 39361
rect 23017 39321 23029 39355
rect 23063 39352 23075 39355
rect 23845 39355 23903 39361
rect 23845 39352 23857 39355
rect 23063 39324 23857 39352
rect 23063 39321 23075 39324
rect 23017 39315 23075 39321
rect 23845 39321 23857 39324
rect 23891 39321 23903 39355
rect 23845 39315 23903 39321
rect 20990 39284 20996 39296
rect 19904 39256 20996 39284
rect 20990 39244 20996 39256
rect 21048 39284 21054 39296
rect 21637 39287 21695 39293
rect 21637 39284 21649 39287
rect 21048 39256 21649 39284
rect 21048 39244 21054 39256
rect 21637 39253 21649 39256
rect 21683 39253 21695 39287
rect 21637 39247 21695 39253
rect 24578 39244 24584 39296
rect 24636 39244 24642 39296
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 7374 39040 7380 39092
rect 7432 39080 7438 39092
rect 8757 39083 8815 39089
rect 8757 39080 8769 39083
rect 7432 39052 8769 39080
rect 7432 39040 7438 39052
rect 8757 39049 8769 39052
rect 8803 39080 8815 39083
rect 9214 39080 9220 39092
rect 8803 39052 9220 39080
rect 8803 39049 8815 39052
rect 8757 39043 8815 39049
rect 9214 39040 9220 39052
rect 9272 39040 9278 39092
rect 9490 39040 9496 39092
rect 9548 39040 9554 39092
rect 10781 39083 10839 39089
rect 10781 39049 10793 39083
rect 10827 39080 10839 39083
rect 10962 39080 10968 39092
rect 10827 39052 10968 39080
rect 10827 39049 10839 39052
rect 10781 39043 10839 39049
rect 10962 39040 10968 39052
rect 11020 39040 11026 39092
rect 12250 39040 12256 39092
rect 12308 39080 12314 39092
rect 14277 39083 14335 39089
rect 12308 39052 14228 39080
rect 12308 39040 12314 39052
rect 8662 38972 8668 39024
rect 8720 39012 8726 39024
rect 10873 39015 10931 39021
rect 10873 39012 10885 39015
rect 8720 38984 10885 39012
rect 8720 38972 8726 38984
rect 10873 38981 10885 38984
rect 10919 39012 10931 39015
rect 11517 39015 11575 39021
rect 11517 39012 11529 39015
rect 10919 38984 11529 39012
rect 10919 38981 10931 38984
rect 10873 38975 10931 38981
rect 11517 38981 11529 38984
rect 11563 39012 11575 39015
rect 11974 39012 11980 39024
rect 11563 38984 11980 39012
rect 11563 38981 11575 38984
rect 11517 38975 11575 38981
rect 11974 38972 11980 38984
rect 12032 38972 12038 39024
rect 12618 39012 12624 39024
rect 12084 38984 12624 39012
rect 10778 38904 10784 38956
rect 10836 38944 10842 38956
rect 12084 38953 12112 38984
rect 12618 38972 12624 38984
rect 12676 38972 12682 39024
rect 14200 39012 14228 39052
rect 14277 39049 14289 39083
rect 14323 39080 14335 39083
rect 14734 39080 14740 39092
rect 14323 39052 14740 39080
rect 14323 39049 14335 39052
rect 14277 39043 14335 39049
rect 14734 39040 14740 39052
rect 14792 39040 14798 39092
rect 15289 39083 15347 39089
rect 15289 39049 15301 39083
rect 15335 39080 15347 39083
rect 15930 39080 15936 39092
rect 15335 39052 15936 39080
rect 15335 39049 15347 39052
rect 15289 39043 15347 39049
rect 15930 39040 15936 39052
rect 15988 39040 15994 39092
rect 16022 39040 16028 39092
rect 16080 39080 16086 39092
rect 19153 39083 19211 39089
rect 19153 39080 19165 39083
rect 16080 39052 19165 39080
rect 16080 39040 16086 39052
rect 19153 39049 19165 39052
rect 19199 39049 19211 39083
rect 19153 39043 19211 39049
rect 20714 39040 20720 39092
rect 20772 39040 20778 39092
rect 24489 39083 24547 39089
rect 24489 39080 24501 39083
rect 22066 39052 24501 39080
rect 17770 39012 17776 39024
rect 14200 38984 17776 39012
rect 17770 38972 17776 38984
rect 17828 38972 17834 39024
rect 19613 39015 19671 39021
rect 19613 38981 19625 39015
rect 19659 39012 19671 39015
rect 20898 39012 20904 39024
rect 19659 38984 20904 39012
rect 19659 38981 19671 38984
rect 19613 38975 19671 38981
rect 20898 38972 20904 38984
rect 20956 38972 20962 39024
rect 12069 38947 12127 38953
rect 10836 38916 11008 38944
rect 10836 38904 10842 38916
rect 8573 38879 8631 38885
rect 8573 38845 8585 38879
rect 8619 38876 8631 38879
rect 8846 38876 8852 38888
rect 8619 38848 8852 38876
rect 8619 38845 8631 38848
rect 8573 38839 8631 38845
rect 8846 38836 8852 38848
rect 8904 38876 8910 38888
rect 9582 38876 9588 38888
rect 8904 38848 9588 38876
rect 8904 38836 8910 38848
rect 9582 38836 9588 38848
rect 9640 38836 9646 38888
rect 10980 38885 11008 38916
rect 12069 38913 12081 38947
rect 12115 38913 12127 38947
rect 14274 38944 14280 38956
rect 13478 38916 14280 38944
rect 12069 38907 12127 38913
rect 14274 38904 14280 38916
rect 14332 38904 14338 38956
rect 18325 38947 18383 38953
rect 18325 38913 18337 38947
rect 18371 38944 18383 38947
rect 19150 38944 19156 38956
rect 18371 38916 19156 38944
rect 18371 38913 18383 38916
rect 18325 38907 18383 38913
rect 19150 38904 19156 38916
rect 19208 38904 19214 38956
rect 19521 38947 19579 38953
rect 19521 38913 19533 38947
rect 19567 38944 19579 38947
rect 19567 38916 19840 38944
rect 19567 38913 19579 38916
rect 19521 38907 19579 38913
rect 9677 38879 9735 38885
rect 9677 38845 9689 38879
rect 9723 38845 9735 38879
rect 9677 38839 9735 38845
rect 10965 38879 11023 38885
rect 10965 38845 10977 38879
rect 11011 38845 11023 38879
rect 10965 38839 11023 38845
rect 12345 38879 12403 38885
rect 12345 38845 12357 38879
rect 12391 38876 12403 38879
rect 14550 38876 14556 38888
rect 12391 38848 14556 38876
rect 12391 38845 12403 38848
rect 12345 38839 12403 38845
rect 8478 38768 8484 38820
rect 8536 38808 8542 38820
rect 9692 38808 9720 38839
rect 14550 38836 14556 38848
rect 14608 38836 14614 38888
rect 15381 38879 15439 38885
rect 15381 38845 15393 38879
rect 15427 38845 15439 38879
rect 15381 38839 15439 38845
rect 15565 38879 15623 38885
rect 15565 38845 15577 38879
rect 15611 38876 15623 38879
rect 15654 38876 15660 38888
rect 15611 38848 15660 38876
rect 15611 38845 15623 38848
rect 15565 38839 15623 38845
rect 8536 38780 9720 38808
rect 10413 38811 10471 38817
rect 8536 38768 8542 38780
rect 10413 38777 10425 38811
rect 10459 38808 10471 38811
rect 11146 38808 11152 38820
rect 10459 38780 11152 38808
rect 10459 38777 10471 38780
rect 10413 38771 10471 38777
rect 11146 38768 11152 38780
rect 11204 38768 11210 38820
rect 14921 38811 14979 38817
rect 14921 38808 14933 38811
rect 13648 38780 14933 38808
rect 9122 38700 9128 38752
rect 9180 38700 9186 38752
rect 11698 38700 11704 38752
rect 11756 38740 11762 38752
rect 13648 38740 13676 38780
rect 14921 38777 14933 38780
rect 14967 38777 14979 38811
rect 15396 38808 15424 38839
rect 15654 38836 15660 38848
rect 15712 38876 15718 38888
rect 16114 38876 16120 38888
rect 15712 38848 16120 38876
rect 15712 38836 15718 38848
rect 16114 38836 16120 38848
rect 16172 38836 16178 38888
rect 16850 38836 16856 38888
rect 16908 38836 16914 38888
rect 18414 38836 18420 38888
rect 18472 38836 18478 38888
rect 18601 38879 18659 38885
rect 18601 38845 18613 38879
rect 18647 38845 18659 38879
rect 19705 38879 19763 38885
rect 19705 38876 19717 38879
rect 18601 38839 18659 38845
rect 19260 38848 19717 38876
rect 18616 38808 18644 38839
rect 19150 38808 19156 38820
rect 15396 38780 16068 38808
rect 18616 38780 19156 38808
rect 14921 38771 14979 38777
rect 15488 38752 15516 38780
rect 16040 38752 16068 38780
rect 19150 38768 19156 38780
rect 19208 38768 19214 38820
rect 11756 38712 13676 38740
rect 13817 38743 13875 38749
rect 11756 38700 11762 38712
rect 13817 38709 13829 38743
rect 13863 38740 13875 38743
rect 13906 38740 13912 38752
rect 13863 38712 13912 38740
rect 13863 38709 13875 38712
rect 13817 38703 13875 38709
rect 13906 38700 13912 38712
rect 13964 38700 13970 38752
rect 15470 38700 15476 38752
rect 15528 38700 15534 38752
rect 16022 38700 16028 38752
rect 16080 38700 16086 38752
rect 16206 38700 16212 38752
rect 16264 38740 16270 38752
rect 17957 38743 18015 38749
rect 17957 38740 17969 38743
rect 16264 38712 17969 38740
rect 16264 38700 16270 38712
rect 17957 38709 17969 38712
rect 18003 38709 18015 38743
rect 17957 38703 18015 38709
rect 18230 38700 18236 38752
rect 18288 38740 18294 38752
rect 18690 38740 18696 38752
rect 18288 38712 18696 38740
rect 18288 38700 18294 38712
rect 18690 38700 18696 38712
rect 18748 38740 18754 38752
rect 19260 38740 19288 38848
rect 19705 38845 19717 38848
rect 19751 38845 19763 38879
rect 19705 38839 19763 38845
rect 19812 38808 19840 38916
rect 19886 38904 19892 38956
rect 19944 38944 19950 38956
rect 22066 38944 22094 39052
rect 24489 39049 24501 39052
rect 24535 39049 24547 39083
rect 24489 39043 24547 39049
rect 23750 38972 23756 39024
rect 23808 39012 23814 39024
rect 24121 39015 24179 39021
rect 24121 39012 24133 39015
rect 23808 38984 24133 39012
rect 23808 38972 23814 38984
rect 24121 38981 24133 38984
rect 24167 39012 24179 39015
rect 25774 39012 25780 39024
rect 24167 38984 25780 39012
rect 24167 38981 24179 38984
rect 24121 38975 24179 38981
rect 25774 38972 25780 38984
rect 25832 38972 25838 39024
rect 24026 38944 24032 38956
rect 19944 38916 22094 38944
rect 23506 38916 24032 38944
rect 19944 38904 19950 38916
rect 24026 38904 24032 38916
rect 24084 38904 24090 38956
rect 24210 38904 24216 38956
rect 24268 38944 24274 38956
rect 24673 38947 24731 38953
rect 24673 38944 24685 38947
rect 24268 38916 24685 38944
rect 24268 38904 24274 38916
rect 24673 38913 24685 38916
rect 24719 38944 24731 38947
rect 24854 38944 24860 38956
rect 24719 38916 24860 38944
rect 24719 38913 24731 38916
rect 24673 38907 24731 38913
rect 24854 38904 24860 38916
rect 24912 38904 24918 38956
rect 25314 38904 25320 38956
rect 25372 38904 25378 38956
rect 20438 38836 20444 38888
rect 20496 38876 20502 38888
rect 20809 38879 20867 38885
rect 20809 38876 20821 38879
rect 20496 38848 20821 38876
rect 20496 38836 20502 38848
rect 20809 38845 20821 38848
rect 20855 38845 20867 38879
rect 20809 38839 20867 38845
rect 20898 38836 20904 38888
rect 20956 38836 20962 38888
rect 22094 38836 22100 38888
rect 22152 38836 22158 38888
rect 22373 38879 22431 38885
rect 22373 38845 22385 38879
rect 22419 38876 22431 38879
rect 23382 38876 23388 38888
rect 22419 38848 23388 38876
rect 22419 38845 22431 38848
rect 22373 38839 22431 38845
rect 23382 38836 23388 38848
rect 23440 38836 23446 38888
rect 21726 38808 21732 38820
rect 19812 38780 21732 38808
rect 21726 38768 21732 38780
rect 21784 38768 21790 38820
rect 23566 38768 23572 38820
rect 23624 38808 23630 38820
rect 25866 38808 25872 38820
rect 23624 38780 25872 38808
rect 23624 38768 23630 38780
rect 25866 38768 25872 38780
rect 25924 38768 25930 38820
rect 18748 38712 19288 38740
rect 20349 38743 20407 38749
rect 18748 38700 18754 38712
rect 20349 38709 20361 38743
rect 20395 38740 20407 38743
rect 21266 38740 21272 38752
rect 20395 38712 21272 38740
rect 20395 38709 20407 38712
rect 20349 38703 20407 38709
rect 21266 38700 21272 38712
rect 21324 38700 21330 38752
rect 23658 38700 23664 38752
rect 23716 38740 23722 38752
rect 23845 38743 23903 38749
rect 23845 38740 23857 38743
rect 23716 38712 23857 38740
rect 23716 38700 23722 38712
rect 23845 38709 23857 38712
rect 23891 38709 23903 38743
rect 23845 38703 23903 38709
rect 25130 38700 25136 38752
rect 25188 38700 25194 38752
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 7558 38496 7564 38548
rect 7616 38536 7622 38548
rect 7837 38539 7895 38545
rect 7837 38536 7849 38539
rect 7616 38508 7849 38536
rect 7616 38496 7622 38508
rect 7837 38505 7849 38508
rect 7883 38505 7895 38539
rect 7837 38499 7895 38505
rect 10413 38539 10471 38545
rect 10413 38505 10425 38539
rect 10459 38536 10471 38539
rect 11054 38536 11060 38548
rect 10459 38508 11060 38536
rect 10459 38505 10471 38508
rect 10413 38499 10471 38505
rect 11054 38496 11060 38508
rect 11112 38496 11118 38548
rect 14182 38496 14188 38548
rect 14240 38536 14246 38548
rect 14277 38539 14335 38545
rect 14277 38536 14289 38539
rect 14240 38508 14289 38536
rect 14240 38496 14246 38508
rect 14277 38505 14289 38508
rect 14323 38505 14335 38539
rect 14277 38499 14335 38505
rect 14826 38496 14832 38548
rect 14884 38536 14890 38548
rect 14884 38508 16068 38536
rect 14884 38496 14890 38508
rect 7650 38428 7656 38480
rect 7708 38468 7714 38480
rect 7708 38440 9904 38468
rect 7708 38428 7714 38440
rect 5445 38403 5503 38409
rect 5445 38369 5457 38403
rect 5491 38400 5503 38403
rect 6454 38400 6460 38412
rect 5491 38372 6460 38400
rect 5491 38369 5503 38372
rect 5445 38363 5503 38369
rect 6454 38360 6460 38372
rect 6512 38360 6518 38412
rect 6914 38360 6920 38412
rect 6972 38400 6978 38412
rect 7193 38403 7251 38409
rect 7193 38400 7205 38403
rect 6972 38372 7205 38400
rect 6972 38360 6978 38372
rect 7193 38369 7205 38372
rect 7239 38400 7251 38403
rect 7834 38400 7840 38412
rect 7239 38372 7840 38400
rect 7239 38369 7251 38372
rect 7193 38363 7251 38369
rect 7834 38360 7840 38372
rect 7892 38360 7898 38412
rect 8496 38409 8524 38440
rect 8481 38403 8539 38409
rect 8481 38369 8493 38403
rect 8527 38369 8539 38403
rect 8481 38363 8539 38369
rect 9122 38360 9128 38412
rect 9180 38400 9186 38412
rect 9677 38403 9735 38409
rect 9677 38400 9689 38403
rect 9180 38372 9689 38400
rect 9180 38360 9186 38372
rect 9677 38369 9689 38372
rect 9723 38369 9735 38403
rect 9677 38363 9735 38369
rect 9769 38403 9827 38409
rect 9769 38369 9781 38403
rect 9815 38369 9827 38403
rect 9769 38363 9827 38369
rect 1302 38292 1308 38344
rect 1360 38332 1366 38344
rect 1765 38335 1823 38341
rect 1765 38332 1777 38335
rect 1360 38304 1777 38332
rect 1360 38292 1366 38304
rect 1765 38301 1777 38304
rect 1811 38332 1823 38335
rect 2041 38335 2099 38341
rect 2041 38332 2053 38335
rect 1811 38304 2053 38332
rect 1811 38301 1823 38304
rect 1765 38295 1823 38301
rect 2041 38301 2053 38304
rect 2087 38301 2099 38335
rect 7374 38332 7380 38344
rect 6854 38304 7380 38332
rect 2041 38295 2099 38301
rect 7374 38292 7380 38304
rect 7432 38292 7438 38344
rect 8205 38335 8263 38341
rect 8205 38301 8217 38335
rect 8251 38332 8263 38335
rect 8294 38332 8300 38344
rect 8251 38304 8300 38332
rect 8251 38301 8263 38304
rect 8205 38295 8263 38301
rect 8294 38292 8300 38304
rect 8352 38292 8358 38344
rect 9214 38292 9220 38344
rect 9272 38332 9278 38344
rect 9784 38332 9812 38363
rect 9272 38304 9812 38332
rect 9876 38332 9904 38440
rect 10134 38428 10140 38480
rect 10192 38468 10198 38480
rect 11885 38471 11943 38477
rect 11885 38468 11897 38471
rect 10192 38440 11897 38468
rect 10192 38428 10198 38440
rect 11885 38437 11897 38440
rect 11931 38437 11943 38471
rect 11885 38431 11943 38437
rect 10870 38360 10876 38412
rect 10928 38400 10934 38412
rect 10965 38403 11023 38409
rect 10965 38400 10977 38403
rect 10928 38372 10977 38400
rect 10928 38360 10934 38372
rect 10965 38369 10977 38372
rect 11011 38369 11023 38403
rect 10965 38363 11023 38369
rect 11422 38360 11428 38412
rect 11480 38400 11486 38412
rect 12345 38403 12403 38409
rect 12345 38400 12357 38403
rect 11480 38372 12357 38400
rect 11480 38360 11486 38372
rect 12345 38369 12357 38372
rect 12391 38369 12403 38403
rect 12345 38363 12403 38369
rect 12437 38403 12495 38409
rect 12437 38369 12449 38403
rect 12483 38369 12495 38403
rect 12437 38363 12495 38369
rect 12452 38332 12480 38363
rect 12710 38360 12716 38412
rect 12768 38400 12774 38412
rect 14829 38403 14887 38409
rect 14829 38400 14841 38403
rect 12768 38372 14841 38400
rect 12768 38360 12774 38372
rect 14829 38369 14841 38372
rect 14875 38369 14887 38403
rect 16040 38400 16068 38508
rect 16574 38496 16580 38548
rect 16632 38536 16638 38548
rect 16632 38508 17264 38536
rect 16632 38496 16638 38508
rect 17236 38468 17264 38508
rect 17770 38496 17776 38548
rect 17828 38536 17834 38548
rect 18141 38539 18199 38545
rect 18141 38536 18153 38539
rect 17828 38508 18153 38536
rect 17828 38496 17834 38508
rect 18141 38505 18153 38508
rect 18187 38505 18199 38539
rect 19150 38536 19156 38548
rect 18141 38499 18199 38505
rect 18248 38508 18736 38536
rect 18248 38468 18276 38508
rect 17236 38440 18276 38468
rect 18598 38428 18604 38480
rect 18656 38428 18662 38480
rect 16209 38403 16267 38409
rect 16209 38400 16221 38403
rect 16040 38372 16221 38400
rect 14829 38363 14887 38369
rect 16209 38369 16221 38372
rect 16255 38400 16267 38403
rect 18230 38400 18236 38412
rect 16255 38372 18236 38400
rect 16255 38369 16267 38372
rect 16209 38363 16267 38369
rect 18230 38360 18236 38372
rect 18288 38360 18294 38412
rect 18616 38400 18644 38428
rect 18708 38409 18736 38508
rect 18892 38508 19156 38536
rect 18892 38480 18920 38508
rect 19150 38496 19156 38508
rect 19208 38496 19214 38548
rect 19334 38496 19340 38548
rect 19392 38536 19398 38548
rect 19429 38539 19487 38545
rect 19429 38536 19441 38539
rect 19392 38508 19441 38536
rect 19392 38496 19398 38508
rect 19429 38505 19441 38508
rect 19475 38505 19487 38539
rect 19429 38499 19487 38505
rect 20162 38496 20168 38548
rect 20220 38536 20226 38548
rect 21450 38536 21456 38548
rect 20220 38508 21456 38536
rect 20220 38496 20226 38508
rect 21450 38496 21456 38508
rect 21508 38496 21514 38548
rect 21634 38496 21640 38548
rect 21692 38536 21698 38548
rect 25590 38536 25596 38548
rect 21692 38508 25596 38536
rect 21692 38496 21698 38508
rect 25590 38496 25596 38508
rect 25648 38496 25654 38548
rect 18874 38428 18880 38480
rect 18932 38428 18938 38480
rect 22370 38428 22376 38480
rect 22428 38468 22434 38480
rect 22830 38468 22836 38480
rect 22428 38440 22836 38468
rect 22428 38428 22434 38440
rect 22830 38428 22836 38440
rect 22888 38428 22894 38480
rect 23382 38428 23388 38480
rect 23440 38468 23446 38480
rect 23440 38440 23796 38468
rect 23440 38428 23446 38440
rect 18340 38372 18644 38400
rect 18693 38403 18751 38409
rect 9876 38304 12480 38332
rect 13909 38335 13967 38341
rect 9272 38292 9278 38304
rect 13909 38301 13921 38335
rect 13955 38332 13967 38335
rect 14274 38332 14280 38344
rect 13955 38304 14280 38332
rect 13955 38301 13967 38304
rect 13909 38295 13967 38301
rect 14274 38292 14280 38304
rect 14332 38292 14338 38344
rect 14737 38335 14795 38341
rect 14737 38301 14749 38335
rect 14783 38332 14795 38335
rect 15194 38332 15200 38344
rect 14783 38304 15200 38332
rect 14783 38301 14795 38304
rect 14737 38295 14795 38301
rect 15194 38292 15200 38304
rect 15252 38292 15258 38344
rect 15930 38292 15936 38344
rect 15988 38292 15994 38344
rect 17770 38292 17776 38344
rect 17828 38332 17834 38344
rect 18340 38332 18368 38372
rect 18693 38369 18705 38403
rect 18739 38369 18751 38403
rect 18693 38363 18751 38369
rect 19426 38360 19432 38412
rect 19484 38400 19490 38412
rect 19981 38403 20039 38409
rect 19981 38400 19993 38403
rect 19484 38372 19993 38400
rect 19484 38360 19490 38372
rect 19981 38369 19993 38372
rect 20027 38369 20039 38403
rect 19981 38363 20039 38369
rect 20254 38360 20260 38412
rect 20312 38400 20318 38412
rect 21085 38403 21143 38409
rect 21085 38400 21097 38403
rect 20312 38372 21097 38400
rect 20312 38360 20318 38372
rect 21085 38369 21097 38372
rect 21131 38369 21143 38403
rect 21085 38363 21143 38369
rect 21174 38360 21180 38412
rect 21232 38360 21238 38412
rect 21910 38360 21916 38412
rect 21968 38400 21974 38412
rect 22465 38403 22523 38409
rect 22465 38400 22477 38403
rect 21968 38372 22477 38400
rect 21968 38360 21974 38372
rect 22465 38369 22477 38372
rect 22511 38369 22523 38403
rect 22465 38363 22523 38369
rect 22554 38360 22560 38412
rect 22612 38400 22618 38412
rect 23658 38400 23664 38412
rect 22612 38372 23664 38400
rect 22612 38360 22618 38372
rect 23658 38360 23664 38372
rect 23716 38360 23722 38412
rect 23768 38409 23796 38440
rect 23753 38403 23811 38409
rect 23753 38369 23765 38403
rect 23799 38369 23811 38403
rect 23753 38363 23811 38369
rect 23842 38360 23848 38412
rect 23900 38400 23906 38412
rect 25133 38403 25191 38409
rect 25133 38400 25145 38403
rect 23900 38372 25145 38400
rect 23900 38360 23906 38372
rect 25133 38369 25145 38372
rect 25179 38369 25191 38403
rect 25133 38363 25191 38369
rect 21634 38332 21640 38344
rect 17828 38304 18368 38332
rect 19812 38304 21640 38332
rect 17828 38292 17834 38304
rect 5721 38267 5779 38273
rect 5721 38233 5733 38267
rect 5767 38233 5779 38267
rect 8570 38264 8576 38276
rect 5721 38227 5779 38233
rect 7392 38236 8576 38264
rect 1581 38199 1639 38205
rect 1581 38165 1593 38199
rect 1627 38196 1639 38199
rect 4062 38196 4068 38208
rect 1627 38168 4068 38196
rect 1627 38165 1639 38168
rect 1581 38159 1639 38165
rect 4062 38156 4068 38168
rect 4120 38156 4126 38208
rect 5736 38196 5764 38227
rect 7392 38196 7420 38236
rect 8570 38224 8576 38236
rect 8628 38224 8634 38276
rect 9585 38267 9643 38273
rect 9585 38233 9597 38267
rect 9631 38264 9643 38267
rect 16298 38264 16304 38276
rect 9631 38236 16304 38264
rect 9631 38233 9643 38236
rect 9585 38227 9643 38233
rect 16298 38224 16304 38236
rect 16356 38224 16362 38276
rect 18414 38264 18420 38276
rect 17434 38236 18420 38264
rect 18414 38224 18420 38236
rect 18472 38224 18478 38276
rect 18601 38267 18659 38273
rect 18601 38233 18613 38267
rect 18647 38264 18659 38267
rect 19812 38264 19840 38304
rect 21634 38292 21640 38304
rect 21692 38292 21698 38344
rect 23934 38332 23940 38344
rect 22066 38304 23940 38332
rect 18647 38236 19840 38264
rect 18647 38233 18659 38236
rect 18601 38227 18659 38233
rect 19886 38224 19892 38276
rect 19944 38224 19950 38276
rect 20438 38224 20444 38276
rect 20496 38264 20502 38276
rect 22066 38264 22094 38304
rect 23934 38292 23940 38304
rect 23992 38292 23998 38344
rect 24946 38292 24952 38344
rect 25004 38332 25010 38344
rect 25041 38335 25099 38341
rect 25041 38332 25053 38335
rect 25004 38304 25053 38332
rect 25004 38292 25010 38304
rect 25041 38301 25053 38304
rect 25087 38301 25099 38335
rect 25041 38295 25099 38301
rect 20496 38236 22094 38264
rect 22373 38267 22431 38273
rect 20496 38224 20502 38236
rect 22373 38233 22385 38267
rect 22419 38264 22431 38267
rect 22419 38236 23244 38264
rect 22419 38233 22431 38236
rect 22373 38227 22431 38233
rect 5736 38168 7420 38196
rect 7561 38199 7619 38205
rect 7561 38165 7573 38199
rect 7607 38196 7619 38199
rect 8202 38196 8208 38208
rect 7607 38168 8208 38196
rect 7607 38165 7619 38168
rect 7561 38159 7619 38165
rect 8202 38156 8208 38168
rect 8260 38196 8266 38208
rect 8297 38199 8355 38205
rect 8297 38196 8309 38199
rect 8260 38168 8309 38196
rect 8260 38156 8266 38168
rect 8297 38165 8309 38168
rect 8343 38165 8355 38199
rect 8297 38159 8355 38165
rect 8386 38156 8392 38208
rect 8444 38196 8450 38208
rect 9217 38199 9275 38205
rect 9217 38196 9229 38199
rect 8444 38168 9229 38196
rect 8444 38156 8450 38168
rect 9217 38165 9229 38168
rect 9263 38165 9275 38199
rect 9217 38159 9275 38165
rect 10778 38156 10784 38208
rect 10836 38156 10842 38208
rect 10870 38156 10876 38208
rect 10928 38156 10934 38208
rect 12250 38156 12256 38208
rect 12308 38156 12314 38208
rect 14645 38199 14703 38205
rect 14645 38165 14657 38199
rect 14691 38196 14703 38199
rect 17218 38196 17224 38208
rect 14691 38168 17224 38196
rect 14691 38165 14703 38168
rect 14645 38159 14703 38165
rect 17218 38156 17224 38168
rect 17276 38156 17282 38208
rect 17681 38199 17739 38205
rect 17681 38165 17693 38199
rect 17727 38196 17739 38199
rect 17862 38196 17868 38208
rect 17727 38168 17868 38196
rect 17727 38165 17739 38168
rect 17681 38159 17739 38165
rect 17862 38156 17868 38168
rect 17920 38156 17926 38208
rect 18506 38156 18512 38208
rect 18564 38156 18570 38208
rect 19334 38156 19340 38208
rect 19392 38196 19398 38208
rect 19797 38199 19855 38205
rect 19797 38196 19809 38199
rect 19392 38168 19809 38196
rect 19392 38156 19398 38168
rect 19797 38165 19809 38168
rect 19843 38165 19855 38199
rect 19797 38159 19855 38165
rect 20622 38156 20628 38208
rect 20680 38156 20686 38208
rect 20990 38156 20996 38208
rect 21048 38156 21054 38208
rect 22005 38199 22063 38205
rect 22005 38165 22017 38199
rect 22051 38196 22063 38199
rect 22278 38196 22284 38208
rect 22051 38168 22284 38196
rect 22051 38165 22063 38168
rect 22005 38159 22063 38165
rect 22278 38156 22284 38168
rect 22336 38156 22342 38208
rect 23216 38205 23244 38236
rect 23474 38224 23480 38276
rect 23532 38264 23538 38276
rect 24302 38264 24308 38276
rect 23532 38236 24308 38264
rect 23532 38224 23538 38236
rect 24302 38224 24308 38236
rect 24360 38224 24366 38276
rect 23201 38199 23259 38205
rect 23201 38165 23213 38199
rect 23247 38165 23259 38199
rect 23201 38159 23259 38165
rect 23566 38156 23572 38208
rect 23624 38156 23630 38208
rect 23658 38156 23664 38208
rect 23716 38156 23722 38208
rect 23750 38156 23756 38208
rect 23808 38196 23814 38208
rect 24581 38199 24639 38205
rect 24581 38196 24593 38199
rect 23808 38168 24593 38196
rect 23808 38156 23814 38168
rect 24581 38165 24593 38168
rect 24627 38165 24639 38199
rect 24581 38159 24639 38165
rect 24670 38156 24676 38208
rect 24728 38196 24734 38208
rect 24949 38199 25007 38205
rect 24949 38196 24961 38199
rect 24728 38168 24961 38196
rect 24728 38156 24734 38168
rect 24949 38165 24961 38168
rect 24995 38165 25007 38199
rect 24949 38159 25007 38165
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 5261 37995 5319 38001
rect 5261 37961 5273 37995
rect 5307 37992 5319 37995
rect 5350 37992 5356 38004
rect 5307 37964 5356 37992
rect 5307 37961 5319 37964
rect 5261 37955 5319 37961
rect 5350 37952 5356 37964
rect 5408 37952 5414 38004
rect 5721 37995 5779 38001
rect 5721 37961 5733 37995
rect 5767 37992 5779 37995
rect 7834 37992 7840 38004
rect 5767 37964 7840 37992
rect 5767 37961 5779 37964
rect 5721 37955 5779 37961
rect 7834 37952 7840 37964
rect 7892 37952 7898 38004
rect 8938 37952 8944 38004
rect 8996 37992 9002 38004
rect 9033 37995 9091 38001
rect 9033 37992 9045 37995
rect 8996 37964 9045 37992
rect 8996 37952 9002 37964
rect 9033 37961 9045 37964
rect 9079 37961 9091 37995
rect 9033 37955 9091 37961
rect 6825 37927 6883 37933
rect 6825 37893 6837 37927
rect 6871 37924 6883 37927
rect 6914 37924 6920 37936
rect 6871 37896 6920 37924
rect 6871 37893 6883 37896
rect 6825 37887 6883 37893
rect 6914 37884 6920 37896
rect 6972 37884 6978 37936
rect 7374 37884 7380 37936
rect 7432 37884 7438 37936
rect 9048 37924 9076 37955
rect 10778 37952 10784 38004
rect 10836 37992 10842 38004
rect 11701 37995 11759 38001
rect 11701 37992 11713 37995
rect 10836 37964 11713 37992
rect 10836 37952 10842 37964
rect 11701 37961 11713 37964
rect 11747 37961 11759 37995
rect 11701 37955 11759 37961
rect 12434 37952 12440 38004
rect 12492 37992 12498 38004
rect 12805 37995 12863 38001
rect 12805 37992 12817 37995
rect 12492 37964 12817 37992
rect 12492 37952 12498 37964
rect 12805 37961 12817 37964
rect 12851 37961 12863 37995
rect 14093 37995 14151 38001
rect 14093 37992 14105 37995
rect 12805 37955 12863 37961
rect 12912 37964 14105 37992
rect 12912 37924 12940 37964
rect 14093 37961 14105 37964
rect 14139 37992 14151 37995
rect 15470 37992 15476 38004
rect 14139 37964 15476 37992
rect 14139 37961 14151 37964
rect 14093 37955 14151 37961
rect 15470 37952 15476 37964
rect 15528 37952 15534 38004
rect 16390 37952 16396 38004
rect 16448 37952 16454 38004
rect 16850 37952 16856 38004
rect 16908 37992 16914 38004
rect 17221 37995 17279 38001
rect 17221 37992 17233 37995
rect 16908 37964 17233 37992
rect 16908 37952 16914 37964
rect 17221 37961 17233 37964
rect 17267 37961 17279 37995
rect 17221 37955 17279 37961
rect 17957 37995 18015 38001
rect 17957 37961 17969 37995
rect 18003 37992 18015 37995
rect 18414 37992 18420 38004
rect 18003 37964 18420 37992
rect 18003 37961 18015 37964
rect 17957 37955 18015 37961
rect 18414 37952 18420 37964
rect 18472 37952 18478 38004
rect 18969 37995 19027 38001
rect 18969 37961 18981 37995
rect 19015 37992 19027 37995
rect 19429 37995 19487 38001
rect 19015 37964 19334 37992
rect 19015 37961 19027 37964
rect 18969 37955 19027 37961
rect 9048 37896 10548 37924
rect 4982 37816 4988 37868
rect 5040 37856 5046 37868
rect 5629 37859 5687 37865
rect 5629 37856 5641 37859
rect 5040 37828 5641 37856
rect 5040 37816 5046 37828
rect 5629 37825 5641 37828
rect 5675 37825 5687 37859
rect 5629 37819 5687 37825
rect 9401 37859 9459 37865
rect 9401 37825 9413 37859
rect 9447 37856 9459 37859
rect 10413 37859 10471 37865
rect 10413 37856 10425 37859
rect 9447 37828 10425 37856
rect 9447 37825 9459 37828
rect 9401 37819 9459 37825
rect 10413 37825 10425 37828
rect 10459 37825 10471 37859
rect 10520 37856 10548 37896
rect 12728 37896 12940 37924
rect 16408 37924 16436 37952
rect 17313 37927 17371 37933
rect 17313 37924 17325 37927
rect 16408 37896 17325 37924
rect 12728 37865 12756 37896
rect 17313 37893 17325 37896
rect 17359 37893 17371 37927
rect 17313 37887 17371 37893
rect 18598 37884 18604 37936
rect 18656 37924 18662 37936
rect 18874 37924 18880 37936
rect 18656 37896 18880 37924
rect 18656 37884 18662 37896
rect 18874 37884 18880 37896
rect 18932 37884 18938 37936
rect 19306 37924 19334 37964
rect 19429 37961 19441 37995
rect 19475 37992 19487 37995
rect 19702 37992 19708 38004
rect 19475 37964 19708 37992
rect 19475 37961 19487 37964
rect 19429 37955 19487 37961
rect 19702 37952 19708 37964
rect 19760 37952 19766 38004
rect 20257 37995 20315 38001
rect 20257 37961 20269 37995
rect 20303 37992 20315 37995
rect 20346 37992 20352 38004
rect 20303 37964 20352 37992
rect 20303 37961 20315 37964
rect 20257 37955 20315 37961
rect 20346 37952 20352 37964
rect 20404 37952 20410 38004
rect 22005 37995 22063 38001
rect 22005 37961 22017 37995
rect 22051 37992 22063 37995
rect 24670 37992 24676 38004
rect 22051 37964 24676 37992
rect 22051 37961 22063 37964
rect 22005 37955 22063 37961
rect 24670 37952 24676 37964
rect 24728 37952 24734 38004
rect 21361 37927 21419 37933
rect 21361 37924 21373 37927
rect 19306 37896 19564 37924
rect 12713 37859 12771 37865
rect 10520 37828 10640 37856
rect 10413 37819 10471 37825
rect 5810 37748 5816 37800
rect 5868 37748 5874 37800
rect 6546 37748 6552 37800
rect 6604 37748 6610 37800
rect 8478 37748 8484 37800
rect 8536 37788 8542 37800
rect 8573 37791 8631 37797
rect 8573 37788 8585 37791
rect 8536 37760 8585 37788
rect 8536 37748 8542 37760
rect 8573 37757 8585 37760
rect 8619 37757 8631 37791
rect 9950 37788 9956 37800
rect 8573 37751 8631 37757
rect 8864 37760 9956 37788
rect 6638 37612 6644 37664
rect 6696 37652 6702 37664
rect 8864 37661 8892 37760
rect 9950 37748 9956 37760
rect 10008 37788 10014 37800
rect 10612 37797 10640 37828
rect 12713 37825 12725 37859
rect 12759 37825 12771 37859
rect 14369 37859 14427 37865
rect 12713 37819 12771 37825
rect 12912 37828 14320 37856
rect 10505 37791 10563 37797
rect 10505 37788 10517 37791
rect 10008 37760 10517 37788
rect 10008 37748 10014 37760
rect 10505 37757 10517 37760
rect 10551 37757 10563 37791
rect 10505 37751 10563 37757
rect 10597 37791 10655 37797
rect 10597 37757 10609 37791
rect 10643 37788 10655 37791
rect 12912 37788 12940 37828
rect 10643 37760 12940 37788
rect 12989 37791 13047 37797
rect 10643 37757 10655 37760
rect 10597 37751 10655 37757
rect 12989 37757 13001 37791
rect 13035 37788 13047 37791
rect 13446 37788 13452 37800
rect 13035 37760 13452 37788
rect 13035 37757 13047 37760
rect 12989 37751 13047 37757
rect 13446 37748 13452 37760
rect 13504 37748 13510 37800
rect 13538 37748 13544 37800
rect 13596 37748 13602 37800
rect 14292 37788 14320 37828
rect 14369 37825 14381 37859
rect 14415 37856 14427 37859
rect 15381 37859 15439 37865
rect 15381 37856 15393 37859
rect 14415 37828 15393 37856
rect 14415 37825 14427 37828
rect 14369 37819 14427 37825
rect 15381 37825 15393 37828
rect 15427 37825 15439 37859
rect 15381 37819 15439 37825
rect 15473 37859 15531 37865
rect 15473 37825 15485 37859
rect 15519 37856 15531 37859
rect 15838 37856 15844 37868
rect 15519 37828 15844 37856
rect 15519 37825 15531 37828
rect 15473 37819 15531 37825
rect 15838 37816 15844 37828
rect 15896 37856 15902 37868
rect 16114 37856 16120 37868
rect 15896 37828 16120 37856
rect 15896 37816 15902 37828
rect 16114 37816 16120 37828
rect 16172 37816 16178 37868
rect 18690 37816 18696 37868
rect 18748 37856 18754 37868
rect 19337 37859 19395 37865
rect 19337 37856 19349 37859
rect 18748 37828 19349 37856
rect 18748 37816 18754 37828
rect 19337 37825 19349 37828
rect 19383 37825 19395 37859
rect 19337 37819 19395 37825
rect 15194 37788 15200 37800
rect 14292 37760 15200 37788
rect 15194 37748 15200 37760
rect 15252 37748 15258 37800
rect 15654 37748 15660 37800
rect 15712 37748 15718 37800
rect 16022 37748 16028 37800
rect 16080 37788 16086 37800
rect 17497 37791 17555 37797
rect 16080 37760 17448 37788
rect 16080 37748 16086 37760
rect 10045 37723 10103 37729
rect 10045 37689 10057 37723
rect 10091 37720 10103 37723
rect 12066 37720 12072 37732
rect 10091 37692 12072 37720
rect 10091 37689 10103 37692
rect 10045 37683 10103 37689
rect 12066 37680 12072 37692
rect 12124 37680 12130 37732
rect 12158 37680 12164 37732
rect 12216 37720 12222 37732
rect 16758 37720 16764 37732
rect 12216 37692 16764 37720
rect 12216 37680 12222 37692
rect 16758 37680 16764 37692
rect 16816 37680 16822 37732
rect 16853 37723 16911 37729
rect 16853 37689 16865 37723
rect 16899 37720 16911 37723
rect 16942 37720 16948 37732
rect 16899 37692 16948 37720
rect 16899 37689 16911 37692
rect 16853 37683 16911 37689
rect 16942 37680 16948 37692
rect 17000 37680 17006 37732
rect 17420 37720 17448 37760
rect 17497 37757 17509 37791
rect 17543 37788 17555 37791
rect 17586 37788 17592 37800
rect 17543 37760 17592 37788
rect 17543 37757 17555 37760
rect 17497 37751 17555 37757
rect 17586 37748 17592 37760
rect 17644 37748 17650 37800
rect 18322 37720 18328 37732
rect 17420 37692 18328 37720
rect 18322 37680 18328 37692
rect 18380 37720 18386 37732
rect 18874 37720 18880 37732
rect 18380 37692 18880 37720
rect 18380 37680 18386 37692
rect 18874 37680 18880 37692
rect 18932 37680 18938 37732
rect 19536 37720 19564 37896
rect 20640 37896 21373 37924
rect 20162 37856 20168 37868
rect 19628 37828 20168 37856
rect 19628 37797 19656 37828
rect 20162 37816 20168 37828
rect 20220 37816 20226 37868
rect 20254 37816 20260 37868
rect 20312 37856 20318 37868
rect 20640 37865 20668 37896
rect 21361 37893 21373 37896
rect 21407 37893 21419 37927
rect 23474 37924 23480 37936
rect 21361 37887 21419 37893
rect 22066 37896 23480 37924
rect 20625 37859 20683 37865
rect 20625 37856 20637 37859
rect 20312 37828 20637 37856
rect 20312 37816 20318 37828
rect 20625 37825 20637 37828
rect 20671 37825 20683 37859
rect 21545 37859 21603 37865
rect 21545 37856 21557 37859
rect 20625 37819 20683 37825
rect 20732 37828 21557 37856
rect 19613 37791 19671 37797
rect 19613 37757 19625 37791
rect 19659 37757 19671 37791
rect 19613 37751 19671 37757
rect 19702 37748 19708 37800
rect 19760 37788 19766 37800
rect 20438 37788 20444 37800
rect 19760 37760 20444 37788
rect 19760 37748 19766 37760
rect 20438 37748 20444 37760
rect 20496 37788 20502 37800
rect 20732 37797 20760 37828
rect 21545 37825 21557 37828
rect 21591 37856 21603 37859
rect 22066 37856 22094 37896
rect 23474 37884 23480 37896
rect 23532 37884 23538 37936
rect 23842 37884 23848 37936
rect 23900 37884 23906 37936
rect 24302 37884 24308 37936
rect 24360 37884 24366 37936
rect 21591 37828 22094 37856
rect 21591 37825 21603 37828
rect 21545 37819 21603 37825
rect 22370 37816 22376 37868
rect 22428 37816 22434 37868
rect 22465 37859 22523 37865
rect 22465 37825 22477 37859
rect 22511 37856 22523 37859
rect 22738 37856 22744 37868
rect 22511 37828 22744 37856
rect 22511 37825 22523 37828
rect 22465 37819 22523 37825
rect 22738 37816 22744 37828
rect 22796 37856 22802 37868
rect 23109 37859 23167 37865
rect 23109 37856 23121 37859
rect 22796 37828 23121 37856
rect 22796 37816 22802 37828
rect 23109 37825 23121 37828
rect 23155 37856 23167 37859
rect 23290 37856 23296 37868
rect 23155 37828 23296 37856
rect 23155 37825 23167 37828
rect 23109 37819 23167 37825
rect 23290 37816 23296 37828
rect 23348 37816 23354 37868
rect 20717 37791 20775 37797
rect 20717 37788 20729 37791
rect 20496 37760 20729 37788
rect 20496 37748 20502 37760
rect 20717 37757 20729 37760
rect 20763 37757 20775 37791
rect 20717 37751 20775 37757
rect 20901 37791 20959 37797
rect 20901 37757 20913 37791
rect 20947 37788 20959 37791
rect 21358 37788 21364 37800
rect 20947 37760 21364 37788
rect 20947 37757 20959 37760
rect 20901 37751 20959 37757
rect 21358 37748 21364 37760
rect 21416 37748 21422 37800
rect 22557 37791 22615 37797
rect 22557 37757 22569 37791
rect 22603 37757 22615 37791
rect 22557 37751 22615 37757
rect 21542 37720 21548 37732
rect 19536 37692 21548 37720
rect 21542 37680 21548 37692
rect 21600 37680 21606 37732
rect 22572 37720 22600 37751
rect 22830 37748 22836 37800
rect 22888 37788 22894 37800
rect 23201 37791 23259 37797
rect 23201 37788 23213 37791
rect 22888 37760 23213 37788
rect 22888 37748 22894 37760
rect 23201 37757 23213 37760
rect 23247 37757 23259 37791
rect 23201 37751 23259 37757
rect 23569 37791 23627 37797
rect 23569 37757 23581 37791
rect 23615 37757 23627 37791
rect 23569 37751 23627 37757
rect 22646 37720 22652 37732
rect 22572 37692 22652 37720
rect 22646 37680 22652 37692
rect 22704 37680 22710 37732
rect 23584 37720 23612 37751
rect 24486 37748 24492 37800
rect 24544 37788 24550 37800
rect 25317 37791 25375 37797
rect 25317 37788 25329 37791
rect 24544 37760 25329 37788
rect 24544 37748 24550 37760
rect 25317 37757 25329 37760
rect 25363 37757 25375 37791
rect 25317 37751 25375 37757
rect 22848 37692 23612 37720
rect 22848 37664 22876 37692
rect 8849 37655 8907 37661
rect 8849 37652 8861 37655
rect 6696 37624 8861 37652
rect 6696 37612 6702 37624
rect 8849 37621 8861 37624
rect 8895 37621 8907 37655
rect 8849 37615 8907 37621
rect 10134 37612 10140 37664
rect 10192 37652 10198 37664
rect 12345 37655 12403 37661
rect 12345 37652 12357 37655
rect 10192 37624 12357 37652
rect 10192 37612 10198 37624
rect 12345 37621 12357 37624
rect 12391 37621 12403 37655
rect 12345 37615 12403 37621
rect 12802 37612 12808 37664
rect 12860 37652 12866 37664
rect 15013 37655 15071 37661
rect 15013 37652 15025 37655
rect 12860 37624 15025 37652
rect 12860 37612 12866 37624
rect 15013 37621 15025 37624
rect 15059 37621 15071 37655
rect 15013 37615 15071 37621
rect 15470 37612 15476 37664
rect 15528 37652 15534 37664
rect 20346 37652 20352 37664
rect 15528 37624 20352 37652
rect 15528 37612 15534 37624
rect 20346 37612 20352 37624
rect 20404 37612 20410 37664
rect 22830 37612 22836 37664
rect 22888 37612 22894 37664
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 8570 37408 8576 37460
rect 8628 37408 8634 37460
rect 10410 37408 10416 37460
rect 10468 37408 10474 37460
rect 13998 37448 14004 37460
rect 13464 37420 14004 37448
rect 8478 37340 8484 37392
rect 8536 37380 8542 37392
rect 12158 37380 12164 37392
rect 8536 37352 12164 37380
rect 8536 37340 8542 37352
rect 12158 37340 12164 37352
rect 12216 37340 12222 37392
rect 7101 37315 7159 37321
rect 7101 37281 7113 37315
rect 7147 37312 7159 37315
rect 8294 37312 8300 37324
rect 7147 37284 8300 37312
rect 7147 37281 7159 37284
rect 7101 37275 7159 37281
rect 8294 37272 8300 37284
rect 8352 37312 8358 37324
rect 9490 37312 9496 37324
rect 8352 37284 9496 37312
rect 8352 37272 8358 37284
rect 9490 37272 9496 37284
rect 9548 37272 9554 37324
rect 11238 37272 11244 37324
rect 11296 37312 11302 37324
rect 11793 37315 11851 37321
rect 11793 37312 11805 37315
rect 11296 37284 11805 37312
rect 11296 37272 11302 37284
rect 11793 37281 11805 37284
rect 11839 37281 11851 37315
rect 11793 37275 11851 37281
rect 11974 37272 11980 37324
rect 12032 37312 12038 37324
rect 13464 37321 13492 37420
rect 13998 37408 14004 37420
rect 14056 37408 14062 37460
rect 14366 37408 14372 37460
rect 14424 37408 14430 37460
rect 15562 37408 15568 37460
rect 15620 37448 15626 37460
rect 15620 37420 15700 37448
rect 15620 37408 15626 37420
rect 14458 37340 14464 37392
rect 14516 37380 14522 37392
rect 14645 37383 14703 37389
rect 14645 37380 14657 37383
rect 14516 37352 14657 37380
rect 14516 37340 14522 37352
rect 14645 37349 14657 37352
rect 14691 37380 14703 37383
rect 15672 37380 15700 37420
rect 16298 37408 16304 37460
rect 16356 37448 16362 37460
rect 17313 37451 17371 37457
rect 17313 37448 17325 37451
rect 16356 37420 17325 37448
rect 16356 37408 16362 37420
rect 17313 37417 17325 37420
rect 17359 37417 17371 37451
rect 17313 37411 17371 37417
rect 18506 37408 18512 37460
rect 18564 37448 18570 37460
rect 20714 37448 20720 37460
rect 18564 37420 20720 37448
rect 18564 37408 18570 37420
rect 20714 37408 20720 37420
rect 20772 37408 20778 37460
rect 23566 37408 23572 37460
rect 23624 37448 23630 37460
rect 23937 37451 23995 37457
rect 23937 37448 23949 37451
rect 23624 37420 23949 37448
rect 23624 37408 23630 37420
rect 23937 37417 23949 37420
rect 23983 37417 23995 37451
rect 23937 37411 23995 37417
rect 14691 37352 15608 37380
rect 15672 37352 16712 37380
rect 14691 37349 14703 37352
rect 14645 37343 14703 37349
rect 15120 37324 15148 37352
rect 15580 37324 15608 37352
rect 12437 37315 12495 37321
rect 12437 37312 12449 37315
rect 12032 37284 12449 37312
rect 12032 37272 12038 37284
rect 12437 37281 12449 37284
rect 12483 37312 12495 37315
rect 13357 37315 13415 37321
rect 13357 37312 13369 37315
rect 12483 37284 13369 37312
rect 12483 37281 12495 37284
rect 12437 37275 12495 37281
rect 13357 37281 13369 37284
rect 13403 37281 13415 37315
rect 13357 37275 13415 37281
rect 13449 37315 13507 37321
rect 13449 37281 13461 37315
rect 13495 37281 13507 37315
rect 15010 37312 15016 37324
rect 13449 37275 13507 37281
rect 14200 37284 15016 37312
rect 6546 37204 6552 37256
rect 6604 37244 6610 37256
rect 6825 37247 6883 37253
rect 6825 37244 6837 37247
rect 6604 37216 6837 37244
rect 6604 37204 6610 37216
rect 6825 37213 6837 37216
rect 6871 37213 6883 37247
rect 6825 37207 6883 37213
rect 9125 37247 9183 37253
rect 9125 37213 9137 37247
rect 9171 37244 9183 37247
rect 10410 37244 10416 37256
rect 9171 37216 10416 37244
rect 9171 37213 9183 37216
rect 9125 37207 9183 37213
rect 6840 37108 6868 37207
rect 10410 37204 10416 37216
rect 10468 37204 10474 37256
rect 11698 37204 11704 37256
rect 11756 37204 11762 37256
rect 13265 37247 13323 37253
rect 13265 37213 13277 37247
rect 13311 37244 13323 37247
rect 13538 37244 13544 37256
rect 13311 37216 13544 37244
rect 13311 37213 13323 37216
rect 13265 37207 13323 37213
rect 13538 37204 13544 37216
rect 13596 37204 13602 37256
rect 14200 37188 14228 37284
rect 15010 37272 15016 37284
rect 15068 37272 15074 37324
rect 15102 37272 15108 37324
rect 15160 37272 15166 37324
rect 15194 37272 15200 37324
rect 15252 37312 15258 37324
rect 15473 37315 15531 37321
rect 15473 37312 15485 37315
rect 15252 37284 15485 37312
rect 15252 37272 15258 37284
rect 15473 37281 15485 37284
rect 15519 37281 15531 37315
rect 15473 37275 15531 37281
rect 15562 37272 15568 37324
rect 15620 37272 15626 37324
rect 16390 37272 16396 37324
rect 16448 37312 16454 37324
rect 16684 37321 16712 37352
rect 17034 37340 17040 37392
rect 17092 37380 17098 37392
rect 17770 37380 17776 37392
rect 17092 37352 17776 37380
rect 17092 37340 17098 37352
rect 17770 37340 17776 37352
rect 17828 37340 17834 37392
rect 18874 37340 18880 37392
rect 18932 37380 18938 37392
rect 18969 37383 19027 37389
rect 18969 37380 18981 37383
rect 18932 37352 18981 37380
rect 18932 37340 18938 37352
rect 18969 37349 18981 37352
rect 19015 37349 19027 37383
rect 18969 37343 19027 37349
rect 23845 37383 23903 37389
rect 23845 37349 23857 37383
rect 23891 37380 23903 37383
rect 24026 37380 24032 37392
rect 23891 37352 24032 37380
rect 23891 37349 23903 37352
rect 23845 37343 23903 37349
rect 16577 37315 16635 37321
rect 16577 37312 16589 37315
rect 16448 37284 16589 37312
rect 16448 37272 16454 37284
rect 16577 37281 16589 37284
rect 16623 37281 16635 37315
rect 16577 37275 16635 37281
rect 16669 37315 16727 37321
rect 16669 37281 16681 37315
rect 16715 37281 16727 37315
rect 16669 37275 16727 37281
rect 16758 37272 16764 37324
rect 16816 37312 16822 37324
rect 17865 37315 17923 37321
rect 17865 37312 17877 37315
rect 16816 37284 17877 37312
rect 16816 37272 16822 37284
rect 17865 37281 17877 37284
rect 17911 37281 17923 37315
rect 18984 37312 19012 37343
rect 24026 37340 24032 37352
rect 24084 37380 24090 37392
rect 24210 37380 24216 37392
rect 24084 37352 24216 37380
rect 24084 37340 24090 37352
rect 24210 37340 24216 37352
rect 24268 37380 24274 37392
rect 24673 37383 24731 37389
rect 24673 37380 24685 37383
rect 24268 37352 24685 37380
rect 24268 37340 24274 37352
rect 24673 37349 24685 37352
rect 24719 37349 24731 37383
rect 24673 37343 24731 37349
rect 18984 37284 19472 37312
rect 17865 37275 17923 37281
rect 14734 37204 14740 37256
rect 14792 37244 14798 37256
rect 16485 37247 16543 37253
rect 16485 37244 16497 37247
rect 14792 37216 16497 37244
rect 14792 37204 14798 37216
rect 16485 37213 16497 37216
rect 16531 37213 16543 37247
rect 16485 37207 16543 37213
rect 17770 37204 17776 37256
rect 17828 37204 17834 37256
rect 19444 37253 19472 37284
rect 20438 37272 20444 37324
rect 20496 37312 20502 37324
rect 20625 37315 20683 37321
rect 20625 37312 20637 37315
rect 20496 37284 20637 37312
rect 20496 37272 20502 37284
rect 20625 37281 20637 37284
rect 20671 37281 20683 37315
rect 20625 37275 20683 37281
rect 24581 37315 24639 37321
rect 24581 37281 24593 37315
rect 24627 37312 24639 37315
rect 24627 37284 25360 37312
rect 24627 37281 24639 37284
rect 24581 37275 24639 37281
rect 25332 37256 25360 37284
rect 19429 37247 19487 37253
rect 19429 37213 19441 37247
rect 19475 37244 19487 37247
rect 21085 37247 21143 37253
rect 21085 37244 21097 37247
rect 19475 37216 21097 37244
rect 19475 37213 19487 37216
rect 19429 37207 19487 37213
rect 21085 37213 21097 37216
rect 21131 37244 21143 37247
rect 21453 37247 21511 37253
rect 21453 37244 21465 37247
rect 21131 37216 21465 37244
rect 21131 37213 21143 37216
rect 21085 37207 21143 37213
rect 21453 37213 21465 37216
rect 21499 37213 21511 37247
rect 21453 37207 21511 37213
rect 22094 37204 22100 37256
rect 22152 37244 22158 37256
rect 22189 37247 22247 37253
rect 22189 37244 22201 37247
rect 22152 37216 22201 37244
rect 22152 37204 22158 37216
rect 22189 37213 22201 37216
rect 22235 37213 22247 37247
rect 22189 37207 22247 37213
rect 22296 37216 25176 37244
rect 7374 37136 7380 37188
rect 7432 37176 7438 37188
rect 9861 37179 9919 37185
rect 9861 37176 9873 37179
rect 7432 37148 7590 37176
rect 8404 37148 9873 37176
rect 7432 37136 7438 37148
rect 8404 37108 8432 37148
rect 9861 37145 9873 37148
rect 9907 37145 9919 37179
rect 9861 37139 9919 37145
rect 11609 37179 11667 37185
rect 11609 37145 11621 37179
rect 11655 37176 11667 37179
rect 12802 37176 12808 37188
rect 11655 37148 12808 37176
rect 11655 37145 11667 37148
rect 11609 37139 11667 37145
rect 12802 37136 12808 37148
rect 12860 37136 12866 37188
rect 14182 37136 14188 37188
rect 14240 37136 14246 37188
rect 17681 37179 17739 37185
rect 17681 37145 17693 37179
rect 17727 37176 17739 37179
rect 20070 37176 20076 37188
rect 17727 37148 20076 37176
rect 17727 37145 17739 37148
rect 17681 37139 17739 37145
rect 20070 37136 20076 37148
rect 20128 37136 20134 37188
rect 20162 37136 20168 37188
rect 20220 37136 20226 37188
rect 20714 37136 20720 37188
rect 20772 37176 20778 37188
rect 22296 37176 22324 37216
rect 20772 37148 22324 37176
rect 24213 37179 24271 37185
rect 20772 37136 20778 37148
rect 24213 37145 24225 37179
rect 24259 37176 24271 37179
rect 24670 37176 24676 37188
rect 24259 37148 24676 37176
rect 24259 37145 24271 37148
rect 24213 37139 24271 37145
rect 24670 37136 24676 37148
rect 24728 37136 24734 37188
rect 6840 37080 8432 37108
rect 10502 37068 10508 37120
rect 10560 37108 10566 37120
rect 11241 37111 11299 37117
rect 11241 37108 11253 37111
rect 10560 37080 11253 37108
rect 10560 37068 10566 37080
rect 11241 37077 11253 37080
rect 11287 37077 11299 37111
rect 11241 37071 11299 37077
rect 12621 37111 12679 37117
rect 12621 37077 12633 37111
rect 12667 37108 12679 37111
rect 12710 37108 12716 37120
rect 12667 37080 12716 37108
rect 12667 37077 12679 37080
rect 12621 37071 12679 37077
rect 12710 37068 12716 37080
rect 12768 37068 12774 37120
rect 12897 37111 12955 37117
rect 12897 37077 12909 37111
rect 12943 37108 12955 37111
rect 14734 37108 14740 37120
rect 12943 37080 14740 37108
rect 12943 37077 12955 37080
rect 12897 37071 12955 37077
rect 14734 37068 14740 37080
rect 14792 37068 14798 37120
rect 14918 37068 14924 37120
rect 14976 37068 14982 37120
rect 15102 37068 15108 37120
rect 15160 37108 15166 37120
rect 15289 37111 15347 37117
rect 15289 37108 15301 37111
rect 15160 37080 15301 37108
rect 15160 37068 15166 37080
rect 15289 37077 15301 37080
rect 15335 37077 15347 37111
rect 15289 37071 15347 37077
rect 15381 37111 15439 37117
rect 15381 37077 15393 37111
rect 15427 37108 15439 37111
rect 15838 37108 15844 37120
rect 15427 37080 15844 37108
rect 15427 37077 15439 37080
rect 15381 37071 15439 37077
rect 15838 37068 15844 37080
rect 15896 37068 15902 37120
rect 16117 37111 16175 37117
rect 16117 37077 16129 37111
rect 16163 37108 16175 37111
rect 16298 37108 16304 37120
rect 16163 37080 16304 37108
rect 16163 37077 16175 37080
rect 16117 37071 16175 37077
rect 16298 37068 16304 37080
rect 16356 37068 16362 37120
rect 18506 37068 18512 37120
rect 18564 37068 18570 37120
rect 25148 37117 25176 37216
rect 25314 37204 25320 37256
rect 25372 37204 25378 37256
rect 25133 37111 25191 37117
rect 25133 37077 25145 37111
rect 25179 37077 25191 37111
rect 25133 37071 25191 37077
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 5534 36904 5540 36916
rect 4080 36876 5540 36904
rect 4080 36836 4108 36876
rect 5534 36864 5540 36876
rect 5592 36904 5598 36916
rect 6546 36904 6552 36916
rect 5592 36876 6552 36904
rect 5592 36864 5598 36876
rect 6546 36864 6552 36876
rect 6604 36864 6610 36916
rect 7466 36864 7472 36916
rect 7524 36864 7530 36916
rect 7929 36907 7987 36913
rect 7929 36873 7941 36907
rect 7975 36904 7987 36907
rect 8386 36904 8392 36916
rect 7975 36876 8392 36904
rect 7975 36873 7987 36876
rect 7929 36867 7987 36873
rect 8386 36864 8392 36876
rect 8444 36864 8450 36916
rect 9030 36864 9036 36916
rect 9088 36864 9094 36916
rect 9398 36864 9404 36916
rect 9456 36904 9462 36916
rect 11609 36907 11667 36913
rect 9456 36876 10548 36904
rect 9456 36864 9462 36876
rect 6089 36839 6147 36845
rect 6089 36836 6101 36839
rect 3988 36808 4108 36836
rect 5474 36808 6101 36836
rect 3988 36777 4016 36808
rect 6089 36805 6101 36808
rect 6135 36836 6147 36839
rect 6914 36836 6920 36848
rect 6135 36808 6920 36836
rect 6135 36805 6147 36808
rect 6089 36799 6147 36805
rect 6914 36796 6920 36808
rect 6972 36836 6978 36848
rect 7374 36836 7380 36848
rect 6972 36808 7380 36836
rect 6972 36796 6978 36808
rect 7374 36796 7380 36808
rect 7432 36836 7438 36848
rect 8662 36836 8668 36848
rect 7432 36808 8668 36836
rect 7432 36796 7438 36808
rect 8662 36796 8668 36808
rect 8720 36796 8726 36848
rect 10229 36839 10287 36845
rect 10229 36805 10241 36839
rect 10275 36836 10287 36839
rect 10410 36836 10416 36848
rect 10275 36808 10416 36836
rect 10275 36805 10287 36808
rect 10229 36799 10287 36805
rect 10410 36796 10416 36808
rect 10468 36796 10474 36848
rect 10520 36836 10548 36876
rect 11609 36873 11621 36907
rect 11655 36904 11667 36907
rect 16022 36904 16028 36916
rect 11655 36876 16028 36904
rect 11655 36873 11667 36876
rect 11609 36867 11667 36873
rect 16022 36864 16028 36876
rect 16080 36864 16086 36916
rect 17034 36864 17040 36916
rect 17092 36864 17098 36916
rect 17405 36907 17463 36913
rect 17405 36873 17417 36907
rect 17451 36904 17463 36907
rect 18506 36904 18512 36916
rect 17451 36876 18512 36904
rect 17451 36873 17463 36876
rect 17405 36867 17463 36873
rect 18506 36864 18512 36876
rect 18564 36864 18570 36916
rect 19610 36864 19616 36916
rect 19668 36904 19674 36916
rect 20441 36907 20499 36913
rect 20441 36904 20453 36907
rect 19668 36876 20453 36904
rect 19668 36864 19674 36876
rect 20441 36873 20453 36876
rect 20487 36873 20499 36907
rect 20441 36867 20499 36873
rect 23842 36864 23848 36916
rect 23900 36904 23906 36916
rect 24581 36907 24639 36913
rect 24581 36904 24593 36907
rect 23900 36876 24593 36904
rect 23900 36864 23906 36876
rect 24581 36873 24593 36876
rect 24627 36873 24639 36907
rect 24581 36867 24639 36873
rect 12621 36839 12679 36845
rect 12621 36836 12633 36839
rect 10520 36808 12633 36836
rect 12621 36805 12633 36808
rect 12667 36805 12679 36839
rect 12621 36799 12679 36805
rect 13817 36839 13875 36845
rect 13817 36805 13829 36839
rect 13863 36836 13875 36839
rect 14642 36836 14648 36848
rect 13863 36808 14648 36836
rect 13863 36805 13875 36808
rect 13817 36799 13875 36805
rect 14642 36796 14648 36808
rect 14700 36796 14706 36848
rect 15194 36796 15200 36848
rect 15252 36836 15258 36848
rect 15565 36839 15623 36845
rect 15565 36836 15577 36839
rect 15252 36808 15577 36836
rect 15252 36796 15258 36808
rect 15565 36805 15577 36808
rect 15611 36805 15623 36839
rect 15565 36799 15623 36805
rect 15838 36796 15844 36848
rect 15896 36836 15902 36848
rect 17770 36836 17776 36848
rect 15896 36808 17776 36836
rect 15896 36796 15902 36808
rect 17770 36796 17776 36808
rect 17828 36796 17834 36848
rect 19886 36796 19892 36848
rect 19944 36836 19950 36848
rect 20349 36839 20407 36845
rect 20349 36836 20361 36839
rect 19944 36808 20361 36836
rect 19944 36796 19950 36808
rect 20349 36805 20361 36808
rect 20395 36805 20407 36839
rect 20349 36799 20407 36805
rect 22646 36796 22652 36848
rect 22704 36836 22710 36848
rect 23109 36839 23167 36845
rect 23109 36836 23121 36839
rect 22704 36808 23121 36836
rect 22704 36796 22710 36808
rect 23109 36805 23121 36808
rect 23155 36836 23167 36839
rect 23382 36836 23388 36848
rect 23155 36808 23388 36836
rect 23155 36805 23167 36808
rect 23109 36799 23167 36805
rect 23382 36796 23388 36808
rect 23440 36796 23446 36848
rect 3973 36771 4031 36777
rect 3973 36737 3985 36771
rect 4019 36737 4031 36771
rect 3973 36731 4031 36737
rect 7837 36771 7895 36777
rect 7837 36737 7849 36771
rect 7883 36768 7895 36771
rect 9122 36768 9128 36780
rect 7883 36740 9128 36768
rect 7883 36737 7895 36740
rect 7837 36731 7895 36737
rect 9122 36728 9128 36740
rect 9180 36728 9186 36780
rect 9306 36728 9312 36780
rect 9364 36768 9370 36780
rect 9401 36771 9459 36777
rect 9401 36768 9413 36771
rect 9364 36740 9413 36768
rect 9364 36728 9370 36740
rect 9401 36737 9413 36740
rect 9447 36737 9459 36771
rect 9401 36731 9459 36737
rect 9493 36771 9551 36777
rect 9493 36737 9505 36771
rect 9539 36768 9551 36771
rect 10594 36768 10600 36780
rect 9539 36740 10600 36768
rect 9539 36737 9551 36740
rect 9493 36731 9551 36737
rect 10594 36728 10600 36740
rect 10652 36728 10658 36780
rect 12069 36771 12127 36777
rect 12069 36737 12081 36771
rect 12115 36768 12127 36771
rect 12529 36771 12587 36777
rect 12529 36768 12541 36771
rect 12115 36740 12541 36768
rect 12115 36737 12127 36740
rect 12069 36731 12127 36737
rect 12529 36737 12541 36740
rect 12575 36768 12587 36771
rect 12710 36768 12716 36780
rect 12575 36740 12716 36768
rect 12575 36737 12587 36740
rect 12529 36731 12587 36737
rect 12710 36728 12716 36740
rect 12768 36728 12774 36780
rect 13446 36728 13452 36780
rect 13504 36768 13510 36780
rect 13725 36771 13783 36777
rect 13725 36768 13737 36771
rect 13504 36740 13737 36768
rect 13504 36728 13510 36740
rect 13725 36737 13737 36740
rect 13771 36768 13783 36771
rect 14182 36768 14188 36780
rect 13771 36740 14188 36768
rect 13771 36737 13783 36740
rect 13725 36731 13783 36737
rect 14182 36728 14188 36740
rect 14240 36728 14246 36780
rect 14921 36771 14979 36777
rect 14921 36737 14933 36771
rect 14967 36768 14979 36771
rect 14967 36740 15884 36768
rect 14967 36737 14979 36740
rect 14921 36731 14979 36737
rect 15856 36712 15884 36740
rect 16758 36728 16764 36780
rect 16816 36768 16822 36780
rect 17497 36771 17555 36777
rect 17497 36768 17509 36771
rect 16816 36740 17509 36768
rect 16816 36728 16822 36740
rect 17497 36737 17509 36740
rect 17543 36737 17555 36771
rect 19978 36768 19984 36780
rect 17497 36731 17555 36737
rect 17696 36740 19984 36768
rect 4249 36703 4307 36709
rect 4249 36669 4261 36703
rect 4295 36700 4307 36703
rect 5442 36700 5448 36712
rect 4295 36672 5448 36700
rect 4295 36669 4307 36672
rect 4249 36663 4307 36669
rect 5442 36660 5448 36672
rect 5500 36700 5506 36712
rect 5721 36703 5779 36709
rect 5500 36672 5672 36700
rect 5500 36660 5506 36672
rect 5644 36632 5672 36672
rect 5721 36669 5733 36703
rect 5767 36700 5779 36703
rect 5810 36700 5816 36712
rect 5767 36672 5816 36700
rect 5767 36669 5779 36672
rect 5721 36663 5779 36669
rect 5810 36660 5816 36672
rect 5868 36660 5874 36712
rect 5994 36660 6000 36712
rect 6052 36700 6058 36712
rect 8021 36703 8079 36709
rect 8021 36700 8033 36703
rect 6052 36672 8033 36700
rect 6052 36660 6058 36672
rect 8021 36669 8033 36672
rect 8067 36669 8079 36703
rect 8021 36663 8079 36669
rect 9582 36660 9588 36712
rect 9640 36660 9646 36712
rect 10962 36660 10968 36712
rect 11020 36660 11026 36712
rect 12802 36660 12808 36712
rect 12860 36660 12866 36712
rect 13906 36660 13912 36712
rect 13964 36660 13970 36712
rect 14366 36660 14372 36712
rect 14424 36700 14430 36712
rect 15013 36703 15071 36709
rect 15013 36700 15025 36703
rect 14424 36672 15025 36700
rect 14424 36660 14430 36672
rect 15013 36669 15025 36672
rect 15059 36669 15071 36703
rect 15013 36663 15071 36669
rect 15102 36660 15108 36712
rect 15160 36660 15166 36712
rect 15838 36660 15844 36712
rect 15896 36660 15902 36712
rect 17696 36709 17724 36740
rect 19978 36728 19984 36740
rect 20036 36728 20042 36780
rect 22094 36728 22100 36780
rect 22152 36768 22158 36780
rect 22830 36768 22836 36780
rect 22152 36740 22836 36768
rect 22152 36728 22158 36740
rect 22830 36728 22836 36740
rect 22888 36728 22894 36780
rect 24210 36728 24216 36780
rect 24268 36728 24274 36780
rect 24670 36728 24676 36780
rect 24728 36768 24734 36780
rect 25314 36768 25320 36780
rect 24728 36740 25320 36768
rect 24728 36728 24734 36740
rect 25314 36728 25320 36740
rect 25372 36728 25378 36780
rect 17681 36703 17739 36709
rect 17681 36669 17693 36703
rect 17727 36669 17739 36703
rect 17681 36663 17739 36669
rect 18874 36660 18880 36712
rect 18932 36700 18938 36712
rect 20533 36703 20591 36709
rect 20533 36700 20545 36703
rect 18932 36672 20545 36700
rect 18932 36660 18938 36672
rect 20533 36669 20545 36672
rect 20579 36669 20591 36703
rect 20533 36663 20591 36669
rect 21910 36660 21916 36712
rect 21968 36700 21974 36712
rect 24762 36700 24768 36712
rect 21968 36672 24768 36700
rect 21968 36660 21974 36672
rect 24762 36660 24768 36672
rect 24820 36660 24826 36712
rect 7650 36632 7656 36644
rect 5644 36604 7656 36632
rect 7650 36592 7656 36604
rect 7708 36592 7714 36644
rect 11974 36592 11980 36644
rect 12032 36632 12038 36644
rect 13924 36632 13952 36660
rect 12032 36604 13952 36632
rect 12032 36592 12038 36604
rect 18966 36592 18972 36644
rect 19024 36632 19030 36644
rect 21928 36632 21956 36660
rect 19024 36604 21956 36632
rect 19024 36592 19030 36604
rect 10778 36524 10784 36576
rect 10836 36564 10842 36576
rect 12161 36567 12219 36573
rect 12161 36564 12173 36567
rect 10836 36536 12173 36564
rect 10836 36524 10842 36536
rect 12161 36533 12173 36536
rect 12207 36533 12219 36567
rect 12161 36527 12219 36533
rect 13357 36567 13415 36573
rect 13357 36533 13369 36567
rect 13403 36564 13415 36567
rect 14458 36564 14464 36576
rect 13403 36536 14464 36564
rect 13403 36533 13415 36536
rect 13357 36527 13415 36533
rect 14458 36524 14464 36536
rect 14516 36524 14522 36576
rect 14550 36524 14556 36576
rect 14608 36524 14614 36576
rect 15838 36524 15844 36576
rect 15896 36524 15902 36576
rect 17218 36524 17224 36576
rect 17276 36564 17282 36576
rect 19981 36567 20039 36573
rect 19981 36564 19993 36567
rect 17276 36536 19993 36564
rect 17276 36524 17282 36536
rect 19981 36533 19993 36536
rect 20027 36533 20039 36567
rect 19981 36527 20039 36533
rect 20070 36524 20076 36576
rect 20128 36564 20134 36576
rect 25133 36567 25191 36573
rect 25133 36564 25145 36567
rect 20128 36536 25145 36564
rect 20128 36524 20134 36536
rect 25133 36533 25145 36536
rect 25179 36533 25191 36567
rect 25133 36527 25191 36533
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 7006 36320 7012 36372
rect 7064 36360 7070 36372
rect 7653 36363 7711 36369
rect 7653 36360 7665 36363
rect 7064 36332 7665 36360
rect 7064 36320 7070 36332
rect 7653 36329 7665 36332
rect 7699 36329 7711 36363
rect 7653 36323 7711 36329
rect 7834 36320 7840 36372
rect 7892 36360 7898 36372
rect 9125 36363 9183 36369
rect 9125 36360 9137 36363
rect 7892 36332 9137 36360
rect 7892 36320 7898 36332
rect 9125 36329 9137 36332
rect 9171 36329 9183 36363
rect 9125 36323 9183 36329
rect 11882 36320 11888 36372
rect 11940 36360 11946 36372
rect 12161 36363 12219 36369
rect 12161 36360 12173 36363
rect 11940 36332 12173 36360
rect 11940 36320 11946 36332
rect 12161 36329 12173 36332
rect 12207 36360 12219 36363
rect 12434 36360 12440 36372
rect 12207 36332 12440 36360
rect 12207 36329 12219 36332
rect 12161 36323 12219 36329
rect 12434 36320 12440 36332
rect 12492 36320 12498 36372
rect 12526 36320 12532 36372
rect 12584 36360 12590 36372
rect 12713 36363 12771 36369
rect 12713 36360 12725 36363
rect 12584 36332 12725 36360
rect 12584 36320 12590 36332
rect 12713 36329 12725 36332
rect 12759 36329 12771 36363
rect 12713 36323 12771 36329
rect 14277 36363 14335 36369
rect 14277 36329 14289 36363
rect 14323 36360 14335 36363
rect 15378 36360 15384 36372
rect 14323 36332 15384 36360
rect 14323 36329 14335 36332
rect 14277 36323 14335 36329
rect 15378 36320 15384 36332
rect 15436 36320 15442 36372
rect 15838 36320 15844 36372
rect 15896 36360 15902 36372
rect 23658 36360 23664 36372
rect 15896 36332 23664 36360
rect 15896 36320 15902 36332
rect 23658 36320 23664 36332
rect 23716 36320 23722 36372
rect 11514 36252 11520 36304
rect 11572 36292 11578 36304
rect 15746 36292 15752 36304
rect 11572 36264 15752 36292
rect 11572 36252 11578 36264
rect 15746 36252 15752 36264
rect 15804 36252 15810 36304
rect 16117 36295 16175 36301
rect 16117 36261 16129 36295
rect 16163 36292 16175 36295
rect 16163 36264 18552 36292
rect 16163 36261 16175 36264
rect 16117 36255 16175 36261
rect 7466 36184 7472 36236
rect 7524 36224 7530 36236
rect 8205 36227 8263 36233
rect 8205 36224 8217 36227
rect 7524 36196 8217 36224
rect 7524 36184 7530 36196
rect 8205 36193 8217 36196
rect 8251 36193 8263 36227
rect 9677 36227 9735 36233
rect 9677 36224 9689 36227
rect 8205 36187 8263 36193
rect 8312 36196 9689 36224
rect 1762 36116 1768 36168
rect 1820 36156 1826 36168
rect 2041 36159 2099 36165
rect 2041 36156 2053 36159
rect 1820 36128 2053 36156
rect 1820 36116 1826 36128
rect 2041 36125 2053 36128
rect 2087 36125 2099 36159
rect 2041 36119 2099 36125
rect 7650 36116 7656 36168
rect 7708 36156 7714 36168
rect 8312 36156 8340 36196
rect 9677 36193 9689 36196
rect 9723 36193 9735 36227
rect 9677 36187 9735 36193
rect 12710 36184 12716 36236
rect 12768 36224 12774 36236
rect 13265 36227 13323 36233
rect 13265 36224 13277 36227
rect 12768 36196 13277 36224
rect 12768 36184 12774 36196
rect 13265 36193 13277 36196
rect 13311 36193 13323 36227
rect 13265 36187 13323 36193
rect 13814 36184 13820 36236
rect 13872 36224 13878 36236
rect 14737 36227 14795 36233
rect 14737 36224 14749 36227
rect 13872 36196 14749 36224
rect 13872 36184 13878 36196
rect 14737 36193 14749 36196
rect 14783 36193 14795 36227
rect 14737 36187 14795 36193
rect 14826 36184 14832 36236
rect 14884 36184 14890 36236
rect 16761 36227 16819 36233
rect 16761 36193 16773 36227
rect 16807 36224 16819 36227
rect 17494 36224 17500 36236
rect 16807 36196 17500 36224
rect 16807 36193 16819 36196
rect 16761 36187 16819 36193
rect 17494 36184 17500 36196
rect 17552 36184 17558 36236
rect 18524 36224 18552 36264
rect 19426 36252 19432 36304
rect 19484 36252 19490 36304
rect 20990 36292 20996 36304
rect 19536 36264 20996 36292
rect 19536 36224 19564 36264
rect 20990 36252 20996 36264
rect 21048 36252 21054 36304
rect 21818 36252 21824 36304
rect 21876 36292 21882 36304
rect 25133 36295 25191 36301
rect 25133 36292 25145 36295
rect 21876 36264 25145 36292
rect 21876 36252 21882 36264
rect 25133 36261 25145 36264
rect 25179 36261 25191 36295
rect 25133 36255 25191 36261
rect 18524 36196 19564 36224
rect 19981 36227 20039 36233
rect 19981 36193 19993 36227
rect 20027 36193 20039 36227
rect 19981 36187 20039 36193
rect 7708 36128 8340 36156
rect 9585 36159 9643 36165
rect 7708 36116 7714 36128
rect 9585 36125 9597 36159
rect 9631 36156 9643 36159
rect 10134 36156 10140 36168
rect 9631 36128 10140 36156
rect 9631 36125 9643 36128
rect 9585 36119 9643 36125
rect 10134 36116 10140 36128
rect 10192 36116 10198 36168
rect 12434 36116 12440 36168
rect 12492 36156 12498 36168
rect 13173 36159 13231 36165
rect 13173 36156 13185 36159
rect 12492 36128 13185 36156
rect 12492 36116 12498 36128
rect 13173 36125 13185 36128
rect 13219 36125 13231 36159
rect 16577 36159 16635 36165
rect 16577 36156 16589 36159
rect 13173 36119 13231 36125
rect 15764 36128 16589 36156
rect 9493 36091 9551 36097
rect 9493 36057 9505 36091
rect 9539 36088 9551 36091
rect 12710 36088 12716 36100
rect 9539 36060 12716 36088
rect 9539 36057 9551 36060
rect 9493 36051 9551 36057
rect 12710 36048 12716 36060
rect 12768 36048 12774 36100
rect 15764 36032 15792 36128
rect 16577 36125 16589 36128
rect 16623 36125 16635 36159
rect 19996 36156 20024 36187
rect 21266 36184 21272 36236
rect 21324 36184 21330 36236
rect 21361 36227 21419 36233
rect 21361 36193 21373 36227
rect 21407 36193 21419 36227
rect 21361 36187 21419 36193
rect 16577 36119 16635 36125
rect 17420 36128 20024 36156
rect 16485 36091 16543 36097
rect 16485 36057 16497 36091
rect 16531 36088 16543 36091
rect 17313 36091 17371 36097
rect 17313 36088 17325 36091
rect 16531 36060 17325 36088
rect 16531 36057 16543 36060
rect 16485 36051 16543 36057
rect 17313 36057 17325 36060
rect 17359 36057 17371 36091
rect 17313 36051 17371 36057
rect 1581 36023 1639 36029
rect 1581 35989 1593 36023
rect 1627 36020 1639 36023
rect 3418 36020 3424 36032
rect 1627 35992 3424 36020
rect 1627 35989 1639 35992
rect 1581 35983 1639 35989
rect 3418 35980 3424 35992
rect 3476 35980 3482 36032
rect 7742 35980 7748 36032
rect 7800 36020 7806 36032
rect 8021 36023 8079 36029
rect 8021 36020 8033 36023
rect 7800 35992 8033 36020
rect 7800 35980 7806 35992
rect 8021 35989 8033 35992
rect 8067 35989 8079 36023
rect 8021 35983 8079 35989
rect 8113 36023 8171 36029
rect 8113 35989 8125 36023
rect 8159 36020 8171 36023
rect 10318 36020 10324 36032
rect 8159 35992 10324 36020
rect 8159 35989 8171 35992
rect 8113 35983 8171 35989
rect 10318 35980 10324 35992
rect 10376 35980 10382 36032
rect 12434 35980 12440 36032
rect 12492 35980 12498 36032
rect 12618 35980 12624 36032
rect 12676 36020 12682 36032
rect 13081 36023 13139 36029
rect 13081 36020 13093 36023
rect 12676 35992 13093 36020
rect 12676 35980 12682 35992
rect 13081 35989 13093 35992
rect 13127 35989 13139 36023
rect 13081 35983 13139 35989
rect 14642 35980 14648 36032
rect 14700 35980 14706 36032
rect 15746 35980 15752 36032
rect 15804 35980 15810 36032
rect 15838 35980 15844 36032
rect 15896 36020 15902 36032
rect 17420 36020 17448 36128
rect 21174 36116 21180 36168
rect 21232 36156 21238 36168
rect 21376 36156 21404 36187
rect 23750 36184 23756 36236
rect 23808 36184 23814 36236
rect 23937 36227 23995 36233
rect 23937 36193 23949 36227
rect 23983 36224 23995 36227
rect 24486 36224 24492 36236
rect 23983 36196 24492 36224
rect 23983 36193 23995 36196
rect 23937 36187 23995 36193
rect 24486 36184 24492 36196
rect 24544 36184 24550 36236
rect 21232 36128 21404 36156
rect 24857 36159 24915 36165
rect 21232 36116 21238 36128
rect 24857 36125 24869 36159
rect 24903 36156 24915 36159
rect 25314 36156 25320 36168
rect 24903 36128 25320 36156
rect 24903 36125 24915 36128
rect 24857 36119 24915 36125
rect 25314 36116 25320 36128
rect 25372 36116 25378 36168
rect 19889 36091 19947 36097
rect 19889 36057 19901 36091
rect 19935 36088 19947 36091
rect 22094 36088 22100 36100
rect 19935 36060 22100 36088
rect 19935 36057 19947 36060
rect 19889 36051 19947 36057
rect 22094 36048 22100 36060
rect 22152 36088 22158 36100
rect 25130 36088 25136 36100
rect 22152 36060 25136 36088
rect 22152 36048 22158 36060
rect 25130 36048 25136 36060
rect 25188 36048 25194 36100
rect 15896 35992 17448 36020
rect 19797 36023 19855 36029
rect 15896 35980 15902 35992
rect 19797 35989 19809 36023
rect 19843 36020 19855 36023
rect 20346 36020 20352 36032
rect 19843 35992 20352 36020
rect 19843 35989 19855 35992
rect 19797 35983 19855 35989
rect 20346 35980 20352 35992
rect 20404 35980 20410 36032
rect 20438 35980 20444 36032
rect 20496 36020 20502 36032
rect 20809 36023 20867 36029
rect 20809 36020 20821 36023
rect 20496 35992 20821 36020
rect 20496 35980 20502 35992
rect 20809 35989 20821 35992
rect 20855 35989 20867 36023
rect 20809 35983 20867 35989
rect 21082 35980 21088 36032
rect 21140 36020 21146 36032
rect 21177 36023 21235 36029
rect 21177 36020 21189 36023
rect 21140 35992 21189 36020
rect 21140 35980 21146 35992
rect 21177 35989 21189 35992
rect 21223 35989 21235 36023
rect 21177 35983 21235 35989
rect 23290 35980 23296 36032
rect 23348 35980 23354 36032
rect 23658 35980 23664 36032
rect 23716 35980 23722 36032
rect 23750 35980 23756 36032
rect 23808 36020 23814 36032
rect 24394 36020 24400 36032
rect 23808 35992 24400 36020
rect 23808 35980 23814 35992
rect 24394 35980 24400 35992
rect 24452 35980 24458 36032
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 5534 35816 5540 35828
rect 4264 35788 5540 35816
rect 4264 35689 4292 35788
rect 5534 35776 5540 35788
rect 5592 35776 5598 35828
rect 5994 35776 6000 35828
rect 6052 35776 6058 35828
rect 6457 35819 6515 35825
rect 6457 35785 6469 35819
rect 6503 35816 6515 35819
rect 6914 35816 6920 35828
rect 6503 35788 6920 35816
rect 6503 35785 6515 35788
rect 6457 35779 6515 35785
rect 6472 35748 6500 35779
rect 6914 35776 6920 35788
rect 6972 35776 6978 35828
rect 13538 35816 13544 35828
rect 9876 35788 13544 35816
rect 5750 35720 6500 35748
rect 8662 35708 8668 35760
rect 8720 35748 8726 35760
rect 8720 35720 8878 35748
rect 8720 35708 8726 35720
rect 4249 35683 4307 35689
rect 4249 35649 4261 35683
rect 4295 35649 4307 35683
rect 4249 35643 4307 35649
rect 4525 35615 4583 35621
rect 4525 35581 4537 35615
rect 4571 35612 4583 35615
rect 5810 35612 5816 35624
rect 4571 35584 5816 35612
rect 4571 35581 4583 35584
rect 4525 35575 4583 35581
rect 5810 35572 5816 35584
rect 5868 35572 5874 35624
rect 8113 35615 8171 35621
rect 8113 35581 8125 35615
rect 8159 35581 8171 35615
rect 8113 35575 8171 35581
rect 8389 35615 8447 35621
rect 8389 35581 8401 35615
rect 8435 35612 8447 35615
rect 9582 35612 9588 35624
rect 8435 35584 9588 35612
rect 8435 35581 8447 35584
rect 8389 35575 8447 35581
rect 8128 35476 8156 35575
rect 9582 35572 9588 35584
rect 9640 35572 9646 35624
rect 8846 35476 8852 35488
rect 8128 35448 8852 35476
rect 8846 35436 8852 35448
rect 8904 35436 8910 35488
rect 9766 35436 9772 35488
rect 9824 35476 9830 35488
rect 9876 35485 9904 35788
rect 13538 35776 13544 35788
rect 13596 35776 13602 35828
rect 13817 35819 13875 35825
rect 13817 35785 13829 35819
rect 13863 35816 13875 35819
rect 13998 35816 14004 35828
rect 13863 35788 14004 35816
rect 13863 35785 13875 35788
rect 13817 35779 13875 35785
rect 13832 35748 13860 35779
rect 13998 35776 14004 35788
rect 14056 35816 14062 35828
rect 14366 35816 14372 35828
rect 14056 35788 14372 35816
rect 14056 35776 14062 35788
rect 14366 35776 14372 35788
rect 14424 35776 14430 35828
rect 14461 35819 14519 35825
rect 14461 35785 14473 35819
rect 14507 35816 14519 35819
rect 14642 35816 14648 35828
rect 14507 35788 14648 35816
rect 14507 35785 14519 35788
rect 14461 35779 14519 35785
rect 14642 35776 14648 35788
rect 14700 35776 14706 35828
rect 17770 35776 17776 35828
rect 17828 35816 17834 35828
rect 20165 35819 20223 35825
rect 20165 35816 20177 35819
rect 17828 35788 20177 35816
rect 17828 35776 17834 35788
rect 20165 35785 20177 35788
rect 20211 35816 20223 35819
rect 24394 35816 24400 35828
rect 20211 35788 24400 35816
rect 20211 35785 20223 35788
rect 20165 35779 20223 35785
rect 24394 35776 24400 35788
rect 24452 35776 24458 35828
rect 13202 35720 13860 35748
rect 14090 35708 14096 35760
rect 14148 35748 14154 35760
rect 17126 35748 17132 35760
rect 14148 35720 17132 35748
rect 14148 35708 14154 35720
rect 17126 35708 17132 35720
rect 17184 35708 17190 35760
rect 17862 35708 17868 35760
rect 17920 35708 17926 35760
rect 18414 35708 18420 35760
rect 18472 35708 18478 35760
rect 20257 35751 20315 35757
rect 20257 35717 20269 35751
rect 20303 35748 20315 35751
rect 20530 35748 20536 35760
rect 20303 35720 20536 35748
rect 20303 35717 20315 35720
rect 20257 35711 20315 35717
rect 20530 35708 20536 35720
rect 20588 35708 20594 35760
rect 23934 35708 23940 35760
rect 23992 35708 23998 35760
rect 19242 35640 19248 35692
rect 19300 35680 19306 35692
rect 21082 35680 21088 35692
rect 19300 35652 21088 35680
rect 19300 35640 19306 35652
rect 21082 35640 21088 35652
rect 21140 35640 21146 35692
rect 22186 35640 22192 35692
rect 22244 35680 22250 35692
rect 22830 35680 22836 35692
rect 22244 35652 22836 35680
rect 22244 35640 22250 35652
rect 22830 35640 22836 35652
rect 22888 35680 22894 35692
rect 23109 35683 23167 35689
rect 23109 35680 23121 35683
rect 22888 35652 23121 35680
rect 22888 35640 22894 35652
rect 23109 35649 23121 35652
rect 23155 35649 23167 35683
rect 23109 35643 23167 35649
rect 10962 35572 10968 35624
rect 11020 35612 11026 35624
rect 11701 35615 11759 35621
rect 11701 35612 11713 35615
rect 11020 35584 11713 35612
rect 11020 35572 11026 35584
rect 11701 35581 11713 35584
rect 11747 35581 11759 35615
rect 11701 35575 11759 35581
rect 11977 35615 12035 35621
rect 11977 35581 11989 35615
rect 12023 35612 12035 35615
rect 13814 35612 13820 35624
rect 12023 35584 13820 35612
rect 12023 35581 12035 35584
rect 11977 35575 12035 35581
rect 13814 35572 13820 35584
rect 13872 35572 13878 35624
rect 17589 35615 17647 35621
rect 17589 35581 17601 35615
rect 17635 35581 17647 35615
rect 17589 35575 17647 35581
rect 13449 35547 13507 35553
rect 13449 35513 13461 35547
rect 13495 35544 13507 35547
rect 13630 35544 13636 35556
rect 13495 35516 13636 35544
rect 13495 35513 13507 35516
rect 13449 35507 13507 35513
rect 13630 35504 13636 35516
rect 13688 35504 13694 35556
rect 9861 35479 9919 35485
rect 9861 35476 9873 35479
rect 9824 35448 9873 35476
rect 9824 35436 9830 35448
rect 9861 35445 9873 35448
rect 9907 35445 9919 35479
rect 9861 35439 9919 35445
rect 10226 35436 10232 35488
rect 10284 35436 10290 35488
rect 15930 35436 15936 35488
rect 15988 35476 15994 35488
rect 17604 35476 17632 35575
rect 18598 35572 18604 35624
rect 18656 35612 18662 35624
rect 20349 35615 20407 35621
rect 20349 35612 20361 35615
rect 18656 35584 20361 35612
rect 18656 35572 18662 35584
rect 20349 35581 20361 35584
rect 20395 35581 20407 35615
rect 20349 35575 20407 35581
rect 22465 35615 22523 35621
rect 22465 35581 22477 35615
rect 22511 35612 22523 35615
rect 22738 35612 22744 35624
rect 22511 35584 22744 35612
rect 22511 35581 22523 35584
rect 22465 35575 22523 35581
rect 22738 35572 22744 35584
rect 22796 35572 22802 35624
rect 23382 35572 23388 35624
rect 23440 35572 23446 35624
rect 23934 35572 23940 35624
rect 23992 35612 23998 35624
rect 25225 35615 25283 35621
rect 25225 35612 25237 35615
rect 23992 35584 25237 35612
rect 23992 35572 23998 35584
rect 25225 35581 25237 35584
rect 25271 35612 25283 35615
rect 25406 35612 25412 35624
rect 25271 35584 25412 35612
rect 25271 35581 25283 35584
rect 25225 35575 25283 35581
rect 25406 35572 25412 35584
rect 25464 35572 25470 35624
rect 19337 35547 19395 35553
rect 19337 35513 19349 35547
rect 19383 35544 19395 35547
rect 21542 35544 21548 35556
rect 19383 35516 21548 35544
rect 19383 35513 19395 35516
rect 19337 35507 19395 35513
rect 21542 35504 21548 35516
rect 21600 35504 21606 35556
rect 17954 35476 17960 35488
rect 15988 35448 17960 35476
rect 15988 35436 15994 35448
rect 17954 35436 17960 35448
rect 18012 35436 18018 35488
rect 19794 35436 19800 35488
rect 19852 35436 19858 35488
rect 20901 35479 20959 35485
rect 20901 35445 20913 35479
rect 20947 35476 20959 35479
rect 20990 35476 20996 35488
rect 20947 35448 20996 35476
rect 20947 35445 20959 35448
rect 20901 35439 20959 35445
rect 20990 35436 20996 35448
rect 21048 35436 21054 35488
rect 22370 35436 22376 35488
rect 22428 35476 22434 35488
rect 22830 35476 22836 35488
rect 22428 35448 22836 35476
rect 22428 35436 22434 35448
rect 22830 35436 22836 35448
rect 22888 35436 22894 35488
rect 23474 35436 23480 35488
rect 23532 35476 23538 35488
rect 24857 35479 24915 35485
rect 24857 35476 24869 35479
rect 23532 35448 24869 35476
rect 23532 35436 23538 35448
rect 24857 35445 24869 35448
rect 24903 35445 24915 35479
rect 24857 35439 24915 35445
rect 25314 35436 25320 35488
rect 25372 35476 25378 35488
rect 25409 35479 25467 35485
rect 25409 35476 25421 35479
rect 25372 35448 25421 35476
rect 25372 35436 25378 35448
rect 25409 35445 25421 35448
rect 25455 35445 25467 35479
rect 25409 35439 25467 35445
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 7650 35232 7656 35284
rect 7708 35272 7714 35284
rect 7837 35275 7895 35281
rect 7837 35272 7849 35275
rect 7708 35244 7849 35272
rect 7708 35232 7714 35244
rect 7837 35241 7849 35244
rect 7883 35241 7895 35275
rect 7837 35235 7895 35241
rect 8205 35275 8263 35281
rect 8205 35241 8217 35275
rect 8251 35272 8263 35275
rect 8662 35272 8668 35284
rect 8251 35244 8668 35272
rect 8251 35241 8263 35244
rect 8205 35235 8263 35241
rect 8662 35232 8668 35244
rect 8720 35232 8726 35284
rect 8754 35232 8760 35284
rect 8812 35272 8818 35284
rect 9309 35275 9367 35281
rect 9309 35272 9321 35275
rect 8812 35244 9321 35272
rect 8812 35232 8818 35244
rect 9309 35241 9321 35244
rect 9355 35241 9367 35275
rect 9309 35235 9367 35241
rect 10594 35232 10600 35284
rect 10652 35272 10658 35284
rect 12989 35275 13047 35281
rect 12989 35272 13001 35275
rect 10652 35244 13001 35272
rect 10652 35232 10658 35244
rect 12989 35241 13001 35244
rect 13035 35241 13047 35275
rect 12989 35235 13047 35241
rect 15654 35232 15660 35284
rect 15712 35272 15718 35284
rect 17129 35275 17187 35281
rect 17129 35272 17141 35275
rect 15712 35244 17141 35272
rect 15712 35232 15718 35244
rect 17129 35241 17141 35244
rect 17175 35241 17187 35275
rect 17129 35235 17187 35241
rect 17497 35275 17555 35281
rect 17497 35241 17509 35275
rect 17543 35272 17555 35275
rect 17862 35272 17868 35284
rect 17543 35244 17868 35272
rect 17543 35241 17555 35244
rect 17497 35235 17555 35241
rect 8570 35164 8576 35216
rect 8628 35204 8634 35216
rect 8628 35176 9904 35204
rect 8628 35164 8634 35176
rect 5534 35096 5540 35148
rect 5592 35136 5598 35148
rect 6086 35136 6092 35148
rect 5592 35108 6092 35136
rect 5592 35096 5598 35108
rect 6086 35096 6092 35108
rect 6144 35096 6150 35148
rect 6365 35139 6423 35145
rect 6365 35105 6377 35139
rect 6411 35136 6423 35139
rect 9766 35136 9772 35148
rect 6411 35108 9772 35136
rect 6411 35105 6423 35108
rect 6365 35099 6423 35105
rect 9766 35096 9772 35108
rect 9824 35096 9830 35148
rect 9876 35145 9904 35176
rect 12342 35164 12348 35216
rect 12400 35204 12406 35216
rect 13446 35204 13452 35216
rect 12400 35176 13452 35204
rect 12400 35164 12406 35176
rect 13446 35164 13452 35176
rect 13504 35164 13510 35216
rect 9861 35139 9919 35145
rect 9861 35105 9873 35139
rect 9907 35105 9919 35139
rect 9861 35099 9919 35105
rect 11054 35096 11060 35148
rect 11112 35136 11118 35148
rect 13541 35139 13599 35145
rect 13541 35136 13553 35139
rect 11112 35108 13553 35136
rect 11112 35096 11118 35108
rect 13541 35105 13553 35108
rect 13587 35105 13599 35139
rect 13541 35099 13599 35105
rect 15381 35139 15439 35145
rect 15381 35105 15393 35139
rect 15427 35136 15439 35139
rect 15746 35136 15752 35148
rect 15427 35108 15752 35136
rect 15427 35105 15439 35108
rect 15381 35099 15439 35105
rect 15746 35096 15752 35108
rect 15804 35096 15810 35148
rect 13449 35071 13507 35077
rect 13449 35037 13461 35071
rect 13495 35068 13507 35071
rect 14550 35068 14556 35080
rect 13495 35040 14556 35068
rect 13495 35037 13507 35040
rect 13449 35031 13507 35037
rect 14550 35028 14556 35040
rect 14608 35028 14614 35080
rect 17512 35068 17540 35235
rect 17862 35232 17868 35244
rect 17920 35272 17926 35284
rect 18322 35272 18328 35284
rect 17920 35244 18328 35272
rect 17920 35232 17926 35244
rect 18322 35232 18328 35244
rect 18380 35232 18386 35284
rect 18414 35232 18420 35284
rect 18472 35272 18478 35284
rect 19692 35275 19750 35281
rect 19692 35272 19704 35275
rect 18472 35244 19704 35272
rect 18472 35232 18478 35244
rect 19692 35241 19704 35244
rect 19738 35272 19750 35275
rect 20898 35272 20904 35284
rect 19738 35244 20904 35272
rect 19738 35241 19750 35244
rect 19692 35235 19750 35241
rect 20898 35232 20904 35244
rect 20956 35232 20962 35284
rect 21082 35232 21088 35284
rect 21140 35272 21146 35284
rect 22370 35272 22376 35284
rect 21140 35244 22376 35272
rect 21140 35232 21146 35244
rect 22370 35232 22376 35244
rect 22428 35232 22434 35284
rect 17954 35096 17960 35148
rect 18012 35136 18018 35148
rect 18322 35136 18328 35148
rect 18012 35108 18328 35136
rect 18012 35096 18018 35108
rect 18322 35096 18328 35108
rect 18380 35136 18386 35148
rect 19429 35139 19487 35145
rect 19429 35136 19441 35139
rect 18380 35108 19441 35136
rect 18380 35096 18386 35108
rect 19429 35105 19441 35108
rect 19475 35136 19487 35139
rect 20162 35136 20168 35148
rect 19475 35108 20168 35136
rect 19475 35105 19487 35108
rect 19429 35099 19487 35105
rect 20162 35096 20168 35108
rect 20220 35096 20226 35148
rect 23014 35096 23020 35148
rect 23072 35136 23078 35148
rect 23934 35136 23940 35148
rect 23072 35108 23940 35136
rect 23072 35096 23078 35108
rect 23934 35096 23940 35108
rect 23992 35136 23998 35148
rect 24210 35136 24216 35148
rect 23992 35108 24216 35136
rect 23992 35096 23998 35108
rect 24210 35096 24216 35108
rect 24268 35136 24274 35148
rect 24397 35139 24455 35145
rect 24397 35136 24409 35139
rect 24268 35108 24409 35136
rect 24268 35096 24274 35108
rect 24397 35105 24409 35108
rect 24443 35105 24455 35139
rect 24397 35099 24455 35105
rect 16790 35040 17540 35068
rect 22186 35028 22192 35080
rect 22244 35068 22250 35080
rect 22281 35071 22339 35077
rect 22281 35068 22293 35071
rect 22244 35040 22293 35068
rect 22244 35028 22250 35040
rect 22281 35037 22293 35040
rect 22327 35037 22339 35071
rect 22281 35031 22339 35037
rect 25314 35028 25320 35080
rect 25372 35028 25378 35080
rect 6914 34960 6920 35012
rect 6972 34960 6978 35012
rect 8662 34960 8668 35012
rect 8720 35000 8726 35012
rect 9677 35003 9735 35009
rect 9677 35000 9689 35003
rect 8720 34972 9689 35000
rect 8720 34960 8726 34972
rect 9677 34969 9689 34972
rect 9723 34969 9735 35003
rect 9677 34963 9735 34969
rect 15657 35003 15715 35009
rect 15657 34969 15669 35003
rect 15703 34969 15715 35003
rect 19610 35000 19616 35012
rect 15657 34963 15715 34969
rect 17052 34972 19616 35000
rect 9769 34935 9827 34941
rect 9769 34901 9781 34935
rect 9815 34932 9827 34935
rect 10134 34932 10140 34944
rect 9815 34904 10140 34932
rect 9815 34901 9827 34904
rect 9769 34895 9827 34901
rect 10134 34892 10140 34904
rect 10192 34892 10198 34944
rect 13357 34935 13415 34941
rect 13357 34901 13369 34935
rect 13403 34932 13415 34935
rect 15562 34932 15568 34944
rect 13403 34904 15568 34932
rect 13403 34901 13415 34904
rect 13357 34895 13415 34901
rect 15562 34892 15568 34904
rect 15620 34892 15626 34944
rect 15672 34932 15700 34963
rect 17052 34932 17080 34972
rect 19610 34960 19616 34972
rect 19668 34960 19674 35012
rect 20990 35000 20996 35012
rect 20930 34972 20996 35000
rect 20990 34960 20996 34972
rect 21048 35000 21054 35012
rect 21048 34972 21588 35000
rect 21048 34960 21054 34972
rect 15672 34904 17080 34932
rect 21174 34892 21180 34944
rect 21232 34892 21238 34944
rect 21560 34941 21588 34972
rect 22554 34960 22560 35012
rect 22612 34960 22618 35012
rect 23014 35000 23020 35012
rect 22940 34972 23020 35000
rect 21545 34935 21603 34941
rect 21545 34901 21557 34935
rect 21591 34932 21603 34935
rect 22940 34932 22968 34972
rect 23014 34960 23020 34972
rect 23072 34960 23078 35012
rect 21591 34904 22968 34932
rect 21591 34901 21603 34904
rect 21545 34895 21603 34901
rect 23382 34892 23388 34944
rect 23440 34932 23446 34944
rect 24029 34935 24087 34941
rect 24029 34932 24041 34935
rect 23440 34904 24041 34932
rect 23440 34892 23446 34904
rect 24029 34901 24041 34904
rect 24075 34901 24087 34935
rect 24029 34895 24087 34901
rect 24946 34892 24952 34944
rect 25004 34932 25010 34944
rect 25133 34935 25191 34941
rect 25133 34932 25145 34935
rect 25004 34904 25145 34932
rect 25004 34892 25010 34904
rect 25133 34901 25145 34904
rect 25179 34901 25191 34935
rect 25133 34895 25191 34901
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 8754 34688 8760 34740
rect 8812 34728 8818 34740
rect 8812 34700 9536 34728
rect 8812 34688 8818 34700
rect 5994 34620 6000 34672
rect 6052 34660 6058 34672
rect 6825 34663 6883 34669
rect 6825 34660 6837 34663
rect 6052 34632 6837 34660
rect 6052 34620 6058 34632
rect 6825 34629 6837 34632
rect 6871 34629 6883 34663
rect 6825 34623 6883 34629
rect 6914 34620 6920 34672
rect 6972 34660 6978 34672
rect 7282 34660 7288 34672
rect 6972 34632 7288 34660
rect 6972 34620 6978 34632
rect 7282 34620 7288 34632
rect 7340 34620 7346 34672
rect 9508 34660 9536 34700
rect 9766 34688 9772 34740
rect 9824 34728 9830 34740
rect 10597 34731 10655 34737
rect 10597 34728 10609 34731
rect 9824 34700 10609 34728
rect 9824 34688 9830 34700
rect 10597 34697 10609 34700
rect 10643 34697 10655 34731
rect 12802 34728 12808 34740
rect 10597 34691 10655 34697
rect 11072 34700 12808 34728
rect 9508 34632 9614 34660
rect 6086 34552 6092 34604
rect 6144 34592 6150 34604
rect 6549 34595 6607 34601
rect 6549 34592 6561 34595
rect 6144 34564 6561 34592
rect 6144 34552 6150 34564
rect 6549 34561 6561 34564
rect 6595 34561 6607 34595
rect 8846 34592 8852 34604
rect 8904 34601 8910 34604
rect 8814 34564 8852 34592
rect 6549 34555 6607 34561
rect 8846 34552 8852 34564
rect 8904 34555 8914 34601
rect 11072 34592 11100 34700
rect 12802 34688 12808 34700
rect 12860 34728 12866 34740
rect 13722 34728 13728 34740
rect 12860 34700 13728 34728
rect 12860 34688 12866 34700
rect 13722 34688 13728 34700
rect 13780 34688 13786 34740
rect 13817 34731 13875 34737
rect 13817 34697 13829 34731
rect 13863 34728 13875 34731
rect 13998 34728 14004 34740
rect 13863 34700 14004 34728
rect 13863 34697 13875 34700
rect 13817 34691 13875 34697
rect 13832 34660 13860 34691
rect 13998 34688 14004 34700
rect 14056 34688 14062 34740
rect 14182 34688 14188 34740
rect 14240 34728 14246 34740
rect 15565 34731 15623 34737
rect 15565 34728 15577 34731
rect 14240 34700 15577 34728
rect 14240 34688 14246 34700
rect 15565 34697 15577 34700
rect 15611 34697 15623 34731
rect 15565 34691 15623 34697
rect 15933 34731 15991 34737
rect 15933 34697 15945 34731
rect 15979 34728 15991 34731
rect 19794 34728 19800 34740
rect 15979 34700 19800 34728
rect 15979 34697 15991 34700
rect 15933 34691 15991 34697
rect 19794 34688 19800 34700
rect 19852 34688 19858 34740
rect 20714 34688 20720 34740
rect 20772 34728 20778 34740
rect 21085 34731 21143 34737
rect 21085 34728 21097 34731
rect 20772 34700 21097 34728
rect 20772 34688 20778 34700
rect 21085 34697 21097 34700
rect 21131 34697 21143 34731
rect 21085 34691 21143 34697
rect 21177 34731 21235 34737
rect 21177 34697 21189 34731
rect 21223 34728 21235 34731
rect 21634 34728 21640 34740
rect 21223 34700 21640 34728
rect 21223 34697 21235 34700
rect 21177 34691 21235 34697
rect 21634 34688 21640 34700
rect 21692 34688 21698 34740
rect 22094 34688 22100 34740
rect 22152 34728 22158 34740
rect 22373 34731 22431 34737
rect 22373 34728 22385 34731
rect 22152 34700 22385 34728
rect 22152 34688 22158 34700
rect 22373 34697 22385 34700
rect 22419 34697 22431 34731
rect 22373 34691 22431 34697
rect 22462 34688 22468 34740
rect 22520 34688 22526 34740
rect 22738 34688 22744 34740
rect 22796 34728 22802 34740
rect 23569 34731 23627 34737
rect 23569 34728 23581 34731
rect 22796 34700 23581 34728
rect 22796 34688 22802 34700
rect 23569 34697 23581 34700
rect 23615 34697 23627 34731
rect 23569 34691 23627 34697
rect 24397 34731 24455 34737
rect 24397 34697 24409 34731
rect 24443 34728 24455 34731
rect 24670 34728 24676 34740
rect 24443 34700 24676 34728
rect 24443 34697 24455 34700
rect 24397 34691 24455 34697
rect 24670 34688 24676 34700
rect 24728 34688 24734 34740
rect 25133 34731 25191 34737
rect 25133 34697 25145 34731
rect 25179 34697 25191 34731
rect 25133 34691 25191 34697
rect 13202 34646 13860 34660
rect 10336 34564 11100 34592
rect 13188 34632 13860 34646
rect 16025 34663 16083 34669
rect 8904 34552 8910 34555
rect 6914 34484 6920 34536
rect 6972 34524 6978 34536
rect 8297 34527 8355 34533
rect 8297 34524 8309 34527
rect 6972 34496 8309 34524
rect 6972 34484 6978 34496
rect 8297 34493 8309 34496
rect 8343 34524 8355 34527
rect 10336 34524 10364 34564
rect 8343 34496 10364 34524
rect 8343 34493 8355 34496
rect 8297 34487 8355 34493
rect 10410 34484 10416 34536
rect 10468 34524 10474 34536
rect 10962 34524 10968 34536
rect 10468 34496 10968 34524
rect 10468 34484 10474 34496
rect 10962 34484 10968 34496
rect 11020 34524 11026 34536
rect 11701 34527 11759 34533
rect 11701 34524 11713 34527
rect 11020 34496 11713 34524
rect 11020 34484 11026 34496
rect 11701 34493 11713 34496
rect 11747 34493 11759 34527
rect 13188 34524 13216 34632
rect 16025 34629 16037 34663
rect 16071 34660 16083 34663
rect 16206 34660 16212 34672
rect 16071 34632 16212 34660
rect 16071 34629 16083 34632
rect 16025 34623 16083 34629
rect 16206 34620 16212 34632
rect 16264 34620 16270 34672
rect 20254 34620 20260 34672
rect 20312 34660 20318 34672
rect 25148 34660 25176 34691
rect 20312 34632 25176 34660
rect 20312 34620 20318 34632
rect 15562 34552 15568 34604
rect 15620 34592 15626 34604
rect 18506 34592 18512 34604
rect 15620 34564 18512 34592
rect 15620 34552 15626 34564
rect 18506 34552 18512 34564
rect 18564 34552 18570 34604
rect 20622 34552 20628 34604
rect 20680 34592 20686 34604
rect 21634 34592 21640 34604
rect 20680 34564 21640 34592
rect 20680 34552 20686 34564
rect 21634 34552 21640 34564
rect 21692 34552 21698 34604
rect 24026 34552 24032 34604
rect 24084 34592 24090 34604
rect 24581 34595 24639 34601
rect 24581 34592 24593 34595
rect 24084 34564 24593 34592
rect 24084 34552 24090 34564
rect 24581 34561 24593 34564
rect 24627 34561 24639 34595
rect 24581 34555 24639 34561
rect 25314 34552 25320 34604
rect 25372 34552 25378 34604
rect 11701 34487 11759 34493
rect 11808 34496 13216 34524
rect 13449 34527 13507 34533
rect 5258 34416 5264 34468
rect 5316 34456 5322 34468
rect 5626 34456 5632 34468
rect 5316 34428 5632 34456
rect 5316 34416 5322 34428
rect 5626 34416 5632 34428
rect 5684 34416 5690 34468
rect 10226 34416 10232 34468
rect 10284 34456 10290 34468
rect 10873 34459 10931 34465
rect 10873 34456 10885 34459
rect 10284 34428 10885 34456
rect 10284 34416 10290 34428
rect 10873 34425 10885 34428
rect 10919 34456 10931 34459
rect 11808 34456 11836 34496
rect 13449 34493 13461 34527
rect 13495 34524 13507 34527
rect 13814 34524 13820 34536
rect 13495 34496 13820 34524
rect 13495 34493 13507 34496
rect 13449 34487 13507 34493
rect 13814 34484 13820 34496
rect 13872 34524 13878 34536
rect 14826 34524 14832 34536
rect 13872 34496 14832 34524
rect 13872 34484 13878 34496
rect 14826 34484 14832 34496
rect 14884 34484 14890 34536
rect 16117 34527 16175 34533
rect 16117 34493 16129 34527
rect 16163 34493 16175 34527
rect 16117 34487 16175 34493
rect 21269 34527 21327 34533
rect 21269 34493 21281 34527
rect 21315 34493 21327 34527
rect 21269 34487 21327 34493
rect 22557 34527 22615 34533
rect 22557 34493 22569 34527
rect 22603 34493 22615 34527
rect 23566 34524 23572 34536
rect 22557 34487 22615 34493
rect 23216 34496 23572 34524
rect 10919 34428 11836 34456
rect 10919 34425 10931 34428
rect 10873 34419 10931 34425
rect 15838 34416 15844 34468
rect 15896 34456 15902 34468
rect 16132 34456 16160 34487
rect 15896 34428 16160 34456
rect 15896 34416 15902 34428
rect 19794 34416 19800 34468
rect 19852 34456 19858 34468
rect 21284 34456 21312 34487
rect 19852 34428 21312 34456
rect 19852 34416 19858 34428
rect 22094 34416 22100 34468
rect 22152 34456 22158 34468
rect 22572 34456 22600 34487
rect 23216 34465 23244 34496
rect 23566 34484 23572 34496
rect 23624 34484 23630 34536
rect 23658 34484 23664 34536
rect 23716 34484 23722 34536
rect 23753 34527 23811 34533
rect 23753 34493 23765 34527
rect 23799 34493 23811 34527
rect 23753 34487 23811 34493
rect 22152 34428 22600 34456
rect 23201 34459 23259 34465
rect 22152 34416 22158 34428
rect 23201 34425 23213 34459
rect 23247 34425 23259 34459
rect 23768 34456 23796 34487
rect 23842 34456 23848 34468
rect 23768 34428 23848 34456
rect 23201 34419 23259 34425
rect 23842 34416 23848 34428
rect 23900 34416 23906 34468
rect 9112 34391 9170 34397
rect 9112 34357 9124 34391
rect 9158 34388 9170 34391
rect 9858 34388 9864 34400
rect 9158 34360 9864 34388
rect 9158 34357 9170 34360
rect 9112 34351 9170 34357
rect 9858 34348 9864 34360
rect 9916 34388 9922 34400
rect 10962 34388 10968 34400
rect 9916 34360 10968 34388
rect 9916 34348 9922 34360
rect 10962 34348 10968 34360
rect 11020 34348 11026 34400
rect 11974 34397 11980 34400
rect 11964 34391 11980 34397
rect 11964 34357 11976 34391
rect 11964 34351 11980 34357
rect 11974 34348 11980 34351
rect 12032 34348 12038 34400
rect 20714 34348 20720 34400
rect 20772 34348 20778 34400
rect 22002 34348 22008 34400
rect 22060 34348 22066 34400
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 7282 34144 7288 34196
rect 7340 34184 7346 34196
rect 7561 34187 7619 34193
rect 7561 34184 7573 34187
rect 7340 34156 7573 34184
rect 7340 34144 7346 34156
rect 7561 34153 7573 34156
rect 7607 34184 7619 34187
rect 8481 34187 8539 34193
rect 8481 34184 8493 34187
rect 7607 34156 8493 34184
rect 7607 34153 7619 34156
rect 7561 34147 7619 34153
rect 8481 34153 8493 34156
rect 8527 34153 8539 34187
rect 8481 34147 8539 34153
rect 9122 34144 9128 34196
rect 9180 34144 9186 34196
rect 10686 34144 10692 34196
rect 10744 34184 10750 34196
rect 12161 34187 12219 34193
rect 12161 34184 12173 34187
rect 10744 34156 12173 34184
rect 10744 34144 10750 34156
rect 12161 34153 12173 34156
rect 12207 34184 12219 34187
rect 12207 34156 12434 34184
rect 12207 34153 12219 34156
rect 12161 34147 12219 34153
rect 12406 34116 12434 34156
rect 13814 34144 13820 34196
rect 13872 34184 13878 34196
rect 17681 34187 17739 34193
rect 13872 34156 17632 34184
rect 13872 34144 13878 34156
rect 17604 34116 17632 34156
rect 17681 34153 17693 34187
rect 17727 34184 17739 34187
rect 18414 34184 18420 34196
rect 17727 34156 18420 34184
rect 17727 34153 17739 34156
rect 17681 34147 17739 34153
rect 18414 34144 18420 34156
rect 18472 34144 18478 34196
rect 19426 34144 19432 34196
rect 19484 34184 19490 34196
rect 20441 34187 20499 34193
rect 20441 34184 20453 34187
rect 19484 34156 20453 34184
rect 19484 34144 19490 34156
rect 20441 34153 20453 34156
rect 20487 34153 20499 34187
rect 20441 34147 20499 34153
rect 25314 34144 25320 34196
rect 25372 34144 25378 34196
rect 25406 34144 25412 34196
rect 25464 34144 25470 34196
rect 20254 34116 20260 34128
rect 12406 34088 13584 34116
rect 17604 34088 20260 34116
rect 5534 34008 5540 34060
rect 5592 34008 5598 34060
rect 5810 34008 5816 34060
rect 5868 34048 5874 34060
rect 7285 34051 7343 34057
rect 7285 34048 7297 34051
rect 5868 34020 7297 34048
rect 5868 34008 5874 34020
rect 7285 34017 7297 34020
rect 7331 34048 7343 34051
rect 9214 34048 9220 34060
rect 7331 34020 9220 34048
rect 7331 34017 7343 34020
rect 7285 34011 7343 34017
rect 9214 34008 9220 34020
rect 9272 34048 9278 34060
rect 9677 34051 9735 34057
rect 9677 34048 9689 34051
rect 9272 34020 9689 34048
rect 9272 34008 9278 34020
rect 9677 34017 9689 34020
rect 9723 34017 9735 34051
rect 12805 34051 12863 34057
rect 12805 34048 12817 34051
rect 9677 34011 9735 34017
rect 10689 34051 10747 34057
rect 10689 34017 10701 34051
rect 10735 34048 10747 34051
rect 10735 34020 12434 34048
rect 10735 34017 10747 34020
rect 10689 34011 10747 34017
rect 10410 33980 10416 33992
rect 9692 33952 10416 33980
rect 9692 33924 9720 33952
rect 10410 33940 10416 33952
rect 10468 33940 10474 33992
rect 12066 33980 12072 33992
rect 11822 33952 12072 33980
rect 12066 33940 12072 33952
rect 12124 33940 12130 33992
rect 12406 33980 12434 34020
rect 13354 34008 13360 34060
rect 13412 34048 13418 34060
rect 13556 34057 13584 34088
rect 20254 34076 20260 34088
rect 20312 34076 20318 34128
rect 20530 34076 20536 34128
rect 20588 34116 20594 34128
rect 21085 34119 21143 34125
rect 21085 34116 21097 34119
rect 20588 34088 21097 34116
rect 20588 34076 20594 34088
rect 21085 34085 21097 34088
rect 21131 34085 21143 34119
rect 21085 34079 21143 34085
rect 13449 34051 13507 34057
rect 13449 34048 13461 34051
rect 13412 34020 13461 34048
rect 13412 34008 13418 34020
rect 13449 34017 13461 34020
rect 13495 34017 13507 34051
rect 13449 34011 13507 34017
rect 13541 34051 13599 34057
rect 13541 34017 13553 34051
rect 13587 34017 13599 34051
rect 13541 34011 13599 34017
rect 15930 34008 15936 34060
rect 15988 34008 15994 34060
rect 17770 34008 17776 34060
rect 17828 34048 17834 34060
rect 19981 34051 20039 34057
rect 19981 34048 19993 34051
rect 17828 34020 19993 34048
rect 17828 34008 17834 34020
rect 19981 34017 19993 34020
rect 20027 34017 20039 34051
rect 19981 34011 20039 34017
rect 21174 34008 21180 34060
rect 21232 34048 21238 34060
rect 21637 34051 21695 34057
rect 21637 34048 21649 34051
rect 21232 34020 21649 34048
rect 21232 34008 21238 34020
rect 21637 34017 21649 34020
rect 21683 34017 21695 34051
rect 21637 34011 21695 34017
rect 22278 34008 22284 34060
rect 22336 34048 22342 34060
rect 22741 34051 22799 34057
rect 22741 34048 22753 34051
rect 22336 34020 22753 34048
rect 22336 34008 22342 34020
rect 22741 34017 22753 34020
rect 22787 34017 22799 34051
rect 22741 34011 22799 34017
rect 22925 34051 22983 34057
rect 22925 34017 22937 34051
rect 22971 34048 22983 34051
rect 23382 34048 23388 34060
rect 22971 34020 23388 34048
rect 22971 34017 22983 34020
rect 22925 34011 22983 34017
rect 23382 34008 23388 34020
rect 23440 34008 23446 34060
rect 13630 33980 13636 33992
rect 12406 33952 13636 33980
rect 13630 33940 13636 33952
rect 13688 33940 13694 33992
rect 14090 33980 14096 33992
rect 13924 33952 14096 33980
rect 5813 33915 5871 33921
rect 5813 33881 5825 33915
rect 5859 33881 5871 33915
rect 7282 33912 7288 33924
rect 7038 33884 7288 33912
rect 5813 33875 5871 33881
rect 5828 33844 5856 33875
rect 7282 33872 7288 33884
rect 7340 33872 7346 33924
rect 7650 33872 7656 33924
rect 7708 33912 7714 33924
rect 9493 33915 9551 33921
rect 9493 33912 9505 33915
rect 7708 33884 9505 33912
rect 7708 33872 7714 33884
rect 9493 33881 9505 33884
rect 9539 33881 9551 33915
rect 9493 33875 9551 33881
rect 9674 33872 9680 33924
rect 9732 33872 9738 33924
rect 12526 33912 12532 33924
rect 11992 33884 12532 33912
rect 7374 33844 7380 33856
rect 5828 33816 7380 33844
rect 7374 33804 7380 33816
rect 7432 33844 7438 33856
rect 8478 33844 8484 33856
rect 7432 33816 8484 33844
rect 7432 33804 7438 33816
rect 8478 33804 8484 33816
rect 8536 33804 8542 33856
rect 9585 33847 9643 33853
rect 9585 33813 9597 33847
rect 9631 33844 9643 33847
rect 11992 33844 12020 33884
rect 12526 33872 12532 33884
rect 12584 33872 12590 33924
rect 13924 33912 13952 33952
rect 14090 33940 14096 33952
rect 14148 33940 14154 33992
rect 17862 33980 17868 33992
rect 17342 33952 17868 33980
rect 17862 33940 17868 33952
rect 17920 33980 17926 33992
rect 17957 33983 18015 33989
rect 17957 33980 17969 33983
rect 17920 33952 17969 33980
rect 17920 33940 17926 33952
rect 17957 33949 17969 33952
rect 18003 33980 18015 33983
rect 19426 33980 19432 33992
rect 18003 33952 19432 33980
rect 18003 33949 18015 33952
rect 17957 33943 18015 33949
rect 19426 33940 19432 33952
rect 19484 33940 19490 33992
rect 19702 33940 19708 33992
rect 19760 33980 19766 33992
rect 19889 33983 19947 33989
rect 19889 33980 19901 33983
rect 19760 33952 19901 33980
rect 19760 33940 19766 33952
rect 19889 33949 19901 33952
rect 19935 33949 19947 33983
rect 19889 33943 19947 33949
rect 21545 33983 21603 33989
rect 21545 33949 21557 33983
rect 21591 33980 21603 33983
rect 21726 33980 21732 33992
rect 21591 33952 21732 33980
rect 21591 33949 21603 33952
rect 21545 33943 21603 33949
rect 21726 33940 21732 33952
rect 21784 33980 21790 33992
rect 21784 33952 22784 33980
rect 21784 33940 21790 33952
rect 13372 33884 13952 33912
rect 9631 33816 12020 33844
rect 9631 33813 9643 33816
rect 9585 33807 9643 33813
rect 12066 33804 12072 33856
rect 12124 33844 12130 33856
rect 12437 33847 12495 33853
rect 12437 33844 12449 33847
rect 12124 33816 12449 33844
rect 12124 33804 12130 33816
rect 12437 33813 12449 33816
rect 12483 33813 12495 33847
rect 12437 33807 12495 33813
rect 12802 33804 12808 33856
rect 12860 33844 12866 33856
rect 12989 33847 13047 33853
rect 12989 33844 13001 33847
rect 12860 33816 13001 33844
rect 12860 33804 12866 33816
rect 12989 33813 13001 33816
rect 13035 33813 13047 33847
rect 12989 33807 13047 33813
rect 13170 33804 13176 33856
rect 13228 33844 13234 33856
rect 13372 33853 13400 33884
rect 14734 33872 14740 33924
rect 14792 33912 14798 33924
rect 16209 33915 16267 33921
rect 16209 33912 16221 33915
rect 14792 33884 16221 33912
rect 14792 33872 14798 33884
rect 16209 33881 16221 33884
rect 16255 33881 16267 33915
rect 19797 33915 19855 33921
rect 16209 33875 16267 33881
rect 17512 33884 19748 33912
rect 13357 33847 13415 33853
rect 13357 33844 13369 33847
rect 13228 33816 13369 33844
rect 13228 33804 13234 33816
rect 13357 33813 13369 33816
rect 13403 33813 13415 33847
rect 13357 33807 13415 33813
rect 13630 33804 13636 33856
rect 13688 33844 13694 33856
rect 13906 33844 13912 33856
rect 13688 33816 13912 33844
rect 13688 33804 13694 33816
rect 13906 33804 13912 33816
rect 13964 33804 13970 33856
rect 13998 33804 14004 33856
rect 14056 33844 14062 33856
rect 17512 33844 17540 33884
rect 14056 33816 17540 33844
rect 14056 33804 14062 33816
rect 19242 33804 19248 33856
rect 19300 33844 19306 33856
rect 19429 33847 19487 33853
rect 19429 33844 19441 33847
rect 19300 33816 19441 33844
rect 19300 33804 19306 33816
rect 19429 33813 19441 33816
rect 19475 33813 19487 33847
rect 19720 33844 19748 33884
rect 19797 33881 19809 33915
rect 19843 33912 19855 33915
rect 20070 33912 20076 33924
rect 19843 33884 20076 33912
rect 19843 33881 19855 33884
rect 19797 33875 19855 33881
rect 20070 33872 20076 33884
rect 20128 33872 20134 33924
rect 20898 33872 20904 33924
rect 20956 33912 20962 33924
rect 22649 33915 22707 33921
rect 22649 33912 22661 33915
rect 20956 33884 22661 33912
rect 20956 33872 20962 33884
rect 22649 33881 22661 33884
rect 22695 33881 22707 33915
rect 22756 33912 22784 33952
rect 24578 33940 24584 33992
rect 24636 33980 24642 33992
rect 24765 33983 24823 33989
rect 24765 33980 24777 33983
rect 24636 33952 24777 33980
rect 24636 33940 24642 33952
rect 24765 33949 24777 33952
rect 24811 33949 24823 33983
rect 24765 33943 24823 33949
rect 25130 33912 25136 33924
rect 22756 33884 25136 33912
rect 22649 33875 22707 33881
rect 25130 33872 25136 33884
rect 25188 33872 25194 33924
rect 20622 33844 20628 33856
rect 19720 33816 20628 33844
rect 19429 33807 19487 33813
rect 20622 33804 20628 33816
rect 20680 33804 20686 33856
rect 21450 33804 21456 33856
rect 21508 33804 21514 33856
rect 22281 33847 22339 33853
rect 22281 33813 22293 33847
rect 22327 33844 22339 33847
rect 22462 33844 22468 33856
rect 22327 33816 22468 33844
rect 22327 33813 22339 33816
rect 22281 33807 22339 33813
rect 22462 33804 22468 33816
rect 22520 33804 22526 33856
rect 24578 33804 24584 33856
rect 24636 33804 24642 33856
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 7193 33643 7251 33649
rect 7193 33609 7205 33643
rect 7239 33640 7251 33643
rect 7282 33640 7288 33652
rect 7239 33612 7288 33640
rect 7239 33609 7251 33612
rect 7193 33603 7251 33609
rect 7282 33600 7288 33612
rect 7340 33600 7346 33652
rect 10318 33600 10324 33652
rect 10376 33640 10382 33652
rect 10413 33643 10471 33649
rect 10413 33640 10425 33643
rect 10376 33612 10425 33640
rect 10376 33600 10382 33612
rect 10413 33609 10425 33612
rect 10459 33609 10471 33643
rect 10413 33603 10471 33609
rect 10778 33600 10784 33652
rect 10836 33640 10842 33652
rect 10873 33643 10931 33649
rect 10873 33640 10885 33643
rect 10836 33612 10885 33640
rect 10836 33600 10842 33612
rect 10873 33609 10885 33612
rect 10919 33609 10931 33643
rect 10873 33603 10931 33609
rect 12710 33600 12716 33652
rect 12768 33640 12774 33652
rect 12897 33643 12955 33649
rect 12897 33640 12909 33643
rect 12768 33612 12909 33640
rect 12768 33600 12774 33612
rect 12897 33609 12909 33612
rect 12943 33609 12955 33643
rect 12897 33603 12955 33609
rect 13357 33643 13415 33649
rect 13357 33609 13369 33643
rect 13403 33640 13415 33643
rect 13814 33640 13820 33652
rect 13403 33612 13820 33640
rect 13403 33609 13415 33612
rect 13357 33603 13415 33609
rect 13814 33600 13820 33612
rect 13872 33600 13878 33652
rect 14550 33640 14556 33652
rect 14108 33612 14556 33640
rect 11790 33532 11796 33584
rect 11848 33572 11854 33584
rect 13998 33572 14004 33584
rect 11848 33544 14004 33572
rect 11848 33532 11854 33544
rect 13998 33532 14004 33544
rect 14056 33532 14062 33584
rect 1302 33464 1308 33516
rect 1360 33504 1366 33516
rect 1765 33507 1823 33513
rect 1765 33504 1777 33507
rect 1360 33476 1777 33504
rect 1360 33464 1366 33476
rect 1765 33473 1777 33476
rect 1811 33504 1823 33507
rect 2041 33507 2099 33513
rect 2041 33504 2053 33507
rect 1811 33476 2053 33504
rect 1811 33473 1823 33476
rect 1765 33467 1823 33473
rect 2041 33473 2053 33476
rect 2087 33473 2099 33507
rect 2041 33467 2099 33473
rect 10781 33507 10839 33513
rect 10781 33473 10793 33507
rect 10827 33504 10839 33507
rect 11606 33504 11612 33516
rect 10827 33476 11612 33504
rect 10827 33473 10839 33476
rect 10781 33467 10839 33473
rect 11606 33464 11612 33476
rect 11664 33464 11670 33516
rect 12434 33464 12440 33516
rect 12492 33504 12498 33516
rect 12618 33504 12624 33516
rect 12492 33476 12624 33504
rect 12492 33464 12498 33476
rect 12618 33464 12624 33476
rect 12676 33464 12682 33516
rect 12710 33464 12716 33516
rect 12768 33504 12774 33516
rect 13170 33504 13176 33516
rect 12768 33476 13176 33504
rect 12768 33464 12774 33476
rect 13170 33464 13176 33476
rect 13228 33464 13234 33516
rect 14108 33513 14136 33612
rect 14550 33600 14556 33612
rect 14608 33640 14614 33652
rect 15930 33640 15936 33652
rect 14608 33612 15936 33640
rect 14608 33600 14614 33612
rect 15930 33600 15936 33612
rect 15988 33600 15994 33652
rect 16209 33643 16267 33649
rect 16209 33609 16221 33643
rect 16255 33640 16267 33643
rect 17862 33640 17868 33652
rect 16255 33612 17868 33640
rect 16255 33609 16267 33612
rect 16209 33603 16267 33609
rect 16224 33572 16252 33603
rect 17862 33600 17868 33612
rect 17920 33640 17926 33652
rect 17920 33612 18460 33640
rect 17920 33600 17926 33612
rect 18322 33572 18328 33584
rect 15594 33544 16252 33572
rect 18064 33544 18328 33572
rect 15948 33516 15976 33544
rect 13265 33507 13323 33513
rect 13265 33473 13277 33507
rect 13311 33473 13323 33507
rect 13265 33467 13323 33473
rect 14093 33507 14151 33513
rect 14093 33473 14105 33507
rect 14139 33473 14151 33507
rect 14093 33467 14151 33473
rect 5350 33396 5356 33448
rect 5408 33396 5414 33448
rect 9766 33396 9772 33448
rect 9824 33396 9830 33448
rect 10965 33439 11023 33445
rect 10965 33405 10977 33439
rect 11011 33405 11023 33439
rect 10965 33399 11023 33405
rect 8294 33328 8300 33380
rect 8352 33368 8358 33380
rect 10980 33368 11008 33399
rect 11422 33396 11428 33448
rect 11480 33436 11486 33448
rect 12529 33439 12587 33445
rect 12529 33436 12541 33439
rect 11480 33408 12541 33436
rect 11480 33396 11486 33408
rect 12529 33405 12541 33408
rect 12575 33436 12587 33439
rect 13280 33436 13308 33467
rect 15930 33464 15936 33516
rect 15988 33464 15994 33516
rect 18064 33513 18092 33544
rect 18322 33532 18328 33544
rect 18380 33532 18386 33584
rect 18432 33572 18460 33612
rect 19610 33600 19616 33652
rect 19668 33640 19674 33652
rect 19797 33643 19855 33649
rect 19797 33640 19809 33643
rect 19668 33612 19809 33640
rect 19668 33600 19674 33612
rect 19797 33609 19809 33612
rect 19843 33609 19855 33643
rect 19797 33603 19855 33609
rect 20257 33643 20315 33649
rect 20257 33609 20269 33643
rect 20303 33609 20315 33643
rect 20257 33603 20315 33609
rect 20272 33572 20300 33603
rect 20622 33600 20628 33652
rect 20680 33600 20686 33652
rect 21450 33600 21456 33652
rect 21508 33640 21514 33652
rect 22649 33643 22707 33649
rect 22649 33640 22661 33643
rect 21508 33612 22661 33640
rect 21508 33600 21514 33612
rect 22649 33609 22661 33612
rect 22695 33609 22707 33643
rect 22649 33603 22707 33609
rect 23658 33572 23664 33584
rect 18432 33544 18814 33572
rect 20272 33544 23664 33572
rect 23658 33532 23664 33544
rect 23716 33532 23722 33584
rect 25406 33572 25412 33584
rect 24978 33558 25412 33572
rect 24964 33544 25412 33558
rect 18049 33507 18107 33513
rect 18049 33473 18061 33507
rect 18095 33473 18107 33507
rect 18049 33467 18107 33473
rect 20717 33507 20775 33513
rect 20717 33473 20729 33507
rect 20763 33504 20775 33507
rect 21266 33504 21272 33516
rect 20763 33476 21272 33504
rect 20763 33473 20775 33476
rect 20717 33467 20775 33473
rect 21266 33464 21272 33476
rect 21324 33464 21330 33516
rect 22186 33464 22192 33516
rect 22244 33504 22250 33516
rect 23477 33507 23535 33513
rect 23477 33504 23489 33507
rect 22244 33476 23489 33504
rect 22244 33464 22250 33476
rect 23477 33473 23489 33476
rect 23523 33473 23535 33507
rect 23477 33467 23535 33473
rect 12575 33408 13308 33436
rect 12575 33405 12587 33408
rect 12529 33399 12587 33405
rect 12636 33380 12664 33408
rect 13538 33396 13544 33448
rect 13596 33396 13602 33448
rect 14369 33439 14427 33445
rect 14369 33405 14381 33439
rect 14415 33436 14427 33439
rect 16298 33436 16304 33448
rect 14415 33408 16304 33436
rect 14415 33405 14427 33408
rect 14369 33399 14427 33405
rect 16298 33396 16304 33408
rect 16356 33396 16362 33448
rect 18325 33439 18383 33445
rect 18325 33405 18337 33439
rect 18371 33436 18383 33439
rect 20901 33439 20959 33445
rect 18371 33408 20668 33436
rect 18371 33405 18383 33408
rect 18325 33399 18383 33405
rect 8352 33340 11008 33368
rect 8352 33328 8358 33340
rect 12618 33328 12624 33380
rect 12676 33328 12682 33380
rect 19426 33328 19432 33380
rect 19484 33368 19490 33380
rect 19886 33368 19892 33380
rect 19484 33340 19892 33368
rect 19484 33328 19490 33340
rect 19886 33328 19892 33340
rect 19944 33328 19950 33380
rect 1581 33303 1639 33309
rect 1581 33269 1593 33303
rect 1627 33300 1639 33303
rect 3510 33300 3516 33312
rect 1627 33272 3516 33300
rect 1627 33269 1639 33272
rect 1581 33263 1639 33269
rect 3510 33260 3516 33272
rect 3568 33260 3574 33312
rect 7190 33260 7196 33312
rect 7248 33300 7254 33312
rect 10594 33300 10600 33312
rect 7248 33272 10600 33300
rect 7248 33260 7254 33272
rect 10594 33260 10600 33272
rect 10652 33260 10658 33312
rect 13446 33260 13452 33312
rect 13504 33300 13510 33312
rect 15838 33300 15844 33312
rect 13504 33272 15844 33300
rect 13504 33260 13510 33272
rect 15838 33260 15844 33272
rect 15896 33260 15902 33312
rect 20640 33300 20668 33408
rect 20901 33405 20913 33439
rect 20947 33405 20959 33439
rect 20901 33399 20959 33405
rect 20916 33368 20944 33399
rect 20990 33396 20996 33448
rect 21048 33436 21054 33448
rect 22005 33439 22063 33445
rect 22005 33436 22017 33439
rect 21048 33408 22017 33436
rect 21048 33396 21054 33408
rect 22005 33405 22017 33408
rect 22051 33405 22063 33439
rect 22005 33399 22063 33405
rect 23750 33396 23756 33448
rect 23808 33396 23814 33448
rect 24210 33396 24216 33448
rect 24268 33436 24274 33448
rect 24964 33436 24992 33544
rect 25406 33532 25412 33544
rect 25464 33532 25470 33584
rect 24268 33408 24992 33436
rect 24268 33396 24274 33408
rect 23474 33368 23480 33380
rect 20916 33340 23480 33368
rect 23474 33328 23480 33340
rect 23532 33328 23538 33380
rect 21174 33300 21180 33312
rect 20640 33272 21180 33300
rect 21174 33260 21180 33272
rect 21232 33260 21238 33312
rect 21266 33260 21272 33312
rect 21324 33260 21330 33312
rect 21358 33260 21364 33312
rect 21416 33300 21422 33312
rect 25225 33303 25283 33309
rect 25225 33300 25237 33303
rect 21416 33272 25237 33300
rect 21416 33260 21422 33272
rect 25225 33269 25237 33272
rect 25271 33269 25283 33303
rect 25225 33263 25283 33269
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 7469 33099 7527 33105
rect 7469 33065 7481 33099
rect 7515 33096 7527 33099
rect 7742 33096 7748 33108
rect 7515 33068 7748 33096
rect 7515 33065 7527 33068
rect 7469 33059 7527 33065
rect 7742 33056 7748 33068
rect 7800 33056 7806 33108
rect 9306 33056 9312 33108
rect 9364 33096 9370 33108
rect 9401 33099 9459 33105
rect 9401 33096 9413 33099
rect 9364 33068 9413 33096
rect 9364 33056 9370 33068
rect 9401 33065 9413 33068
rect 9447 33065 9459 33099
rect 9401 33059 9459 33065
rect 10594 33056 10600 33108
rect 10652 33056 10658 33108
rect 10870 33056 10876 33108
rect 10928 33096 10934 33108
rect 11149 33099 11207 33105
rect 11149 33096 11161 33099
rect 10928 33068 11161 33096
rect 10928 33056 10934 33068
rect 11149 33065 11161 33068
rect 11195 33065 11207 33099
rect 15102 33096 15108 33108
rect 11149 33059 11207 33065
rect 12406 33068 15108 33096
rect 9674 32988 9680 33040
rect 9732 33028 9738 33040
rect 12406 33028 12434 33068
rect 15102 33056 15108 33068
rect 15160 33056 15166 33108
rect 17402 33096 17408 33108
rect 16592 33068 17408 33096
rect 9732 33000 12434 33028
rect 9732 32988 9738 33000
rect 13630 32988 13636 33040
rect 13688 33028 13694 33040
rect 15749 33031 15807 33037
rect 15749 33028 15761 33031
rect 13688 33000 15761 33028
rect 13688 32988 13694 33000
rect 5261 32963 5319 32969
rect 5261 32929 5273 32963
rect 5307 32960 5319 32963
rect 5534 32960 5540 32972
rect 5307 32932 5540 32960
rect 5307 32929 5319 32932
rect 5261 32923 5319 32929
rect 5534 32920 5540 32932
rect 5592 32920 5598 32972
rect 7009 32963 7067 32969
rect 7009 32929 7021 32963
rect 7055 32960 7067 32963
rect 7466 32960 7472 32972
rect 7055 32932 7472 32960
rect 7055 32929 7067 32932
rect 7009 32923 7067 32929
rect 7466 32920 7472 32932
rect 7524 32920 7530 32972
rect 8113 32963 8171 32969
rect 8113 32929 8125 32963
rect 8159 32960 8171 32963
rect 8294 32960 8300 32972
rect 8159 32932 8300 32960
rect 8159 32929 8171 32932
rect 8113 32923 8171 32929
rect 7282 32892 7288 32904
rect 6670 32864 7288 32892
rect 7282 32852 7288 32864
rect 7340 32852 7346 32904
rect 8128 32892 8156 32923
rect 8294 32920 8300 32932
rect 8352 32920 8358 32972
rect 9858 32920 9864 32972
rect 9916 32960 9922 32972
rect 9953 32963 10011 32969
rect 9953 32960 9965 32963
rect 9916 32932 9965 32960
rect 9916 32920 9922 32932
rect 9953 32929 9965 32932
rect 9999 32960 10011 32963
rect 11146 32960 11152 32972
rect 9999 32932 11152 32960
rect 9999 32929 10011 32932
rect 9953 32923 10011 32929
rect 11146 32920 11152 32932
rect 11204 32920 11210 32972
rect 11514 32920 11520 32972
rect 11572 32960 11578 32972
rect 11701 32963 11759 32969
rect 11701 32960 11713 32963
rect 11572 32932 11713 32960
rect 11572 32920 11578 32932
rect 11701 32929 11713 32932
rect 11747 32929 11759 32963
rect 11701 32923 11759 32929
rect 14458 32920 14464 32972
rect 14516 32960 14522 32972
rect 14737 32963 14795 32969
rect 14737 32960 14749 32963
rect 14516 32932 14749 32960
rect 14516 32920 14522 32932
rect 14737 32929 14749 32932
rect 14783 32929 14795 32963
rect 14737 32923 14795 32929
rect 14826 32920 14832 32972
rect 14884 32920 14890 32972
rect 7668 32864 8156 32892
rect 5537 32827 5595 32833
rect 5537 32793 5549 32827
rect 5583 32793 5595 32827
rect 5537 32787 5595 32793
rect 5552 32756 5580 32787
rect 7668 32756 7696 32864
rect 9766 32852 9772 32904
rect 9824 32852 9830 32904
rect 15396 32892 15424 33000
rect 15749 32997 15761 33000
rect 15795 32997 15807 33031
rect 15749 32991 15807 32997
rect 15470 32920 15476 32972
rect 15528 32960 15534 32972
rect 16592 32969 16620 33068
rect 17402 33056 17408 33068
rect 17460 33056 17466 33108
rect 19797 33099 19855 33105
rect 19797 33065 19809 33099
rect 19843 33096 19855 33099
rect 20898 33096 20904 33108
rect 19843 33068 20904 33096
rect 19843 33065 19855 33068
rect 19797 33059 19855 33065
rect 20898 33056 20904 33068
rect 20956 33056 20962 33108
rect 21174 33056 21180 33108
rect 21232 33096 21238 33108
rect 21818 33096 21824 33108
rect 21232 33068 21824 33096
rect 21232 33056 21238 33068
rect 21818 33056 21824 33068
rect 21876 33056 21882 33108
rect 22189 33099 22247 33105
rect 22189 33065 22201 33099
rect 22235 33096 22247 33099
rect 23934 33096 23940 33108
rect 22235 33068 23940 33096
rect 22235 33065 22247 33068
rect 22189 33059 22247 33065
rect 23934 33056 23940 33068
rect 23992 33056 23998 33108
rect 17221 33031 17279 33037
rect 17221 32997 17233 33031
rect 17267 33028 17279 33031
rect 17862 33028 17868 33040
rect 17267 33000 17868 33028
rect 17267 32997 17279 33000
rect 17221 32991 17279 32997
rect 17862 32988 17868 33000
rect 17920 32988 17926 33040
rect 22554 33028 22560 33040
rect 21376 33000 22560 33028
rect 16577 32963 16635 32969
rect 16577 32960 16589 32963
rect 15528 32932 16589 32960
rect 15528 32920 15534 32932
rect 16577 32929 16589 32932
rect 16623 32929 16635 32963
rect 16577 32923 16635 32929
rect 16761 32963 16819 32969
rect 16761 32929 16773 32963
rect 16807 32960 16819 32963
rect 16942 32960 16948 32972
rect 16807 32932 16948 32960
rect 16807 32929 16819 32932
rect 16761 32923 16819 32929
rect 16942 32920 16948 32932
rect 17000 32920 17006 32972
rect 20441 32963 20499 32969
rect 20441 32929 20453 32963
rect 20487 32960 20499 32963
rect 21376 32960 21404 33000
rect 22554 32988 22560 33000
rect 22612 32988 22618 33040
rect 20487 32932 21404 32960
rect 20487 32929 20499 32932
rect 20441 32923 20499 32929
rect 21450 32920 21456 32972
rect 21508 32920 21514 32972
rect 21542 32920 21548 32972
rect 21600 32920 21606 32972
rect 16485 32895 16543 32901
rect 16485 32892 16497 32895
rect 15396 32864 16497 32892
rect 16485 32861 16497 32864
rect 16531 32861 16543 32895
rect 16485 32855 16543 32861
rect 20165 32895 20223 32901
rect 20165 32861 20177 32895
rect 20211 32892 20223 32895
rect 20990 32892 20996 32904
rect 20211 32864 20996 32892
rect 20211 32861 20223 32864
rect 20165 32855 20223 32861
rect 20990 32852 20996 32864
rect 21048 32852 21054 32904
rect 22370 32852 22376 32904
rect 22428 32852 22434 32904
rect 22738 32852 22744 32904
rect 22796 32852 22802 32904
rect 24857 32895 24915 32901
rect 24857 32861 24869 32895
rect 24903 32892 24915 32895
rect 25314 32892 25320 32904
rect 24903 32864 25320 32892
rect 24903 32861 24915 32864
rect 24857 32855 24915 32861
rect 25314 32852 25320 32864
rect 25372 32852 25378 32904
rect 7742 32784 7748 32836
rect 7800 32824 7806 32836
rect 7929 32827 7987 32833
rect 7929 32824 7941 32827
rect 7800 32796 7941 32824
rect 7800 32784 7806 32796
rect 7929 32793 7941 32796
rect 7975 32793 7987 32827
rect 7929 32787 7987 32793
rect 10873 32827 10931 32833
rect 10873 32793 10885 32827
rect 10919 32824 10931 32827
rect 11609 32827 11667 32833
rect 11609 32824 11621 32827
rect 10919 32796 11621 32824
rect 10919 32793 10931 32796
rect 10873 32787 10931 32793
rect 11609 32793 11621 32796
rect 11655 32824 11667 32827
rect 11698 32824 11704 32836
rect 11655 32796 11704 32824
rect 11655 32793 11667 32796
rect 11609 32787 11667 32793
rect 11698 32784 11704 32796
rect 11756 32824 11762 32836
rect 19429 32827 19487 32833
rect 19429 32824 19441 32827
rect 11756 32796 12434 32824
rect 11756 32784 11762 32796
rect 5552 32728 7696 32756
rect 7834 32716 7840 32768
rect 7892 32716 7898 32768
rect 9490 32716 9496 32768
rect 9548 32756 9554 32768
rect 9861 32759 9919 32765
rect 9861 32756 9873 32759
rect 9548 32728 9873 32756
rect 9548 32716 9554 32728
rect 9861 32725 9873 32728
rect 9907 32725 9919 32759
rect 9861 32719 9919 32725
rect 10594 32716 10600 32768
rect 10652 32756 10658 32768
rect 11517 32759 11575 32765
rect 11517 32756 11529 32759
rect 10652 32728 11529 32756
rect 10652 32716 10658 32728
rect 11517 32725 11529 32728
rect 11563 32756 11575 32759
rect 11882 32756 11888 32768
rect 11563 32728 11888 32756
rect 11563 32725 11575 32728
rect 11517 32719 11575 32725
rect 11882 32716 11888 32728
rect 11940 32716 11946 32768
rect 12406 32756 12434 32796
rect 14016 32796 19441 32824
rect 14016 32768 14044 32796
rect 19429 32793 19441 32796
rect 19475 32824 19487 32827
rect 20257 32827 20315 32833
rect 20257 32824 20269 32827
rect 19475 32796 20269 32824
rect 19475 32793 19487 32796
rect 19429 32787 19487 32793
rect 20257 32793 20269 32796
rect 20303 32793 20315 32827
rect 20257 32787 20315 32793
rect 20364 32796 25176 32824
rect 13998 32756 14004 32768
rect 12406 32728 14004 32756
rect 13998 32716 14004 32728
rect 14056 32716 14062 32768
rect 14277 32759 14335 32765
rect 14277 32725 14289 32759
rect 14323 32756 14335 32759
rect 14458 32756 14464 32768
rect 14323 32728 14464 32756
rect 14323 32725 14335 32728
rect 14277 32719 14335 32725
rect 14458 32716 14464 32728
rect 14516 32716 14522 32768
rect 14642 32716 14648 32768
rect 14700 32716 14706 32768
rect 16114 32716 16120 32768
rect 16172 32716 16178 32768
rect 16206 32716 16212 32768
rect 16264 32756 16270 32768
rect 20364 32756 20392 32796
rect 16264 32728 20392 32756
rect 16264 32716 16270 32728
rect 20898 32716 20904 32768
rect 20956 32756 20962 32768
rect 20993 32759 21051 32765
rect 20993 32756 21005 32759
rect 20956 32728 21005 32756
rect 20956 32716 20962 32728
rect 20993 32725 21005 32728
rect 21039 32725 21051 32759
rect 20993 32719 21051 32725
rect 21082 32716 21088 32768
rect 21140 32756 21146 32768
rect 21266 32756 21272 32768
rect 21140 32728 21272 32756
rect 21140 32716 21146 32728
rect 21266 32716 21272 32728
rect 21324 32756 21330 32768
rect 21361 32759 21419 32765
rect 21361 32756 21373 32759
rect 21324 32728 21373 32756
rect 21324 32716 21330 32728
rect 21361 32725 21373 32728
rect 21407 32756 21419 32759
rect 22833 32759 22891 32765
rect 22833 32756 22845 32759
rect 21407 32728 22845 32756
rect 21407 32725 21419 32728
rect 21361 32719 21419 32725
rect 22833 32725 22845 32728
rect 22879 32756 22891 32759
rect 24118 32756 24124 32768
rect 22879 32728 24124 32756
rect 22879 32725 22891 32728
rect 22833 32719 22891 32725
rect 24118 32716 24124 32728
rect 24176 32716 24182 32768
rect 25148 32765 25176 32796
rect 25133 32759 25191 32765
rect 25133 32725 25145 32759
rect 25179 32725 25191 32759
rect 25133 32719 25191 32725
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 4614 32512 4620 32564
rect 4672 32512 4678 32564
rect 4982 32512 4988 32564
rect 5040 32512 5046 32564
rect 5350 32512 5356 32564
rect 5408 32512 5414 32564
rect 6917 32555 6975 32561
rect 6917 32521 6929 32555
rect 6963 32552 6975 32555
rect 7834 32552 7840 32564
rect 6963 32524 7840 32552
rect 6963 32521 6975 32524
rect 6917 32515 6975 32521
rect 7834 32512 7840 32524
rect 7892 32512 7898 32564
rect 8478 32552 8484 32564
rect 8220 32524 8484 32552
rect 4632 32484 4660 32512
rect 4890 32484 4896 32496
rect 4632 32456 4896 32484
rect 4890 32444 4896 32456
rect 4948 32484 4954 32496
rect 5445 32487 5503 32493
rect 5445 32484 5457 32487
rect 4948 32456 5457 32484
rect 4948 32444 4954 32456
rect 5445 32453 5457 32456
rect 5491 32453 5503 32487
rect 5445 32447 5503 32453
rect 5534 32444 5540 32496
rect 5592 32444 5598 32496
rect 7282 32444 7288 32496
rect 7340 32484 7346 32496
rect 8220 32484 8248 32524
rect 8478 32512 8484 32524
rect 8536 32512 8542 32564
rect 9309 32555 9367 32561
rect 9309 32521 9321 32555
rect 9355 32552 9367 32555
rect 9674 32552 9680 32564
rect 9355 32524 9680 32552
rect 9355 32521 9367 32524
rect 9309 32515 9367 32521
rect 9674 32512 9680 32524
rect 9732 32512 9738 32564
rect 11977 32555 12035 32561
rect 11977 32521 11989 32555
rect 12023 32552 12035 32555
rect 14642 32552 14648 32564
rect 12023 32524 14648 32552
rect 12023 32521 12035 32524
rect 11977 32515 12035 32521
rect 14642 32512 14648 32524
rect 14700 32512 14706 32564
rect 15212 32524 16160 32552
rect 7340 32456 8326 32484
rect 7340 32444 7346 32456
rect 12250 32444 12256 32496
rect 12308 32484 12314 32496
rect 15212 32484 15240 32524
rect 12308 32456 15240 32484
rect 16132 32484 16160 32524
rect 16206 32512 16212 32564
rect 16264 32552 16270 32564
rect 17313 32555 17371 32561
rect 17313 32552 17325 32555
rect 16264 32524 17325 32552
rect 16264 32512 16270 32524
rect 17313 32521 17325 32524
rect 17359 32521 17371 32555
rect 17313 32515 17371 32521
rect 17678 32512 17684 32564
rect 17736 32552 17742 32564
rect 21177 32555 21235 32561
rect 17736 32524 20300 32552
rect 17736 32512 17742 32524
rect 18417 32487 18475 32493
rect 18417 32484 18429 32487
rect 16132 32456 18429 32484
rect 12308 32444 12314 32456
rect 18417 32453 18429 32456
rect 18463 32453 18475 32487
rect 18417 32447 18475 32453
rect 18509 32487 18567 32493
rect 18509 32453 18521 32487
rect 18555 32484 18567 32487
rect 18690 32484 18696 32496
rect 18555 32456 18696 32484
rect 18555 32453 18567 32456
rect 18509 32447 18567 32453
rect 5552 32416 5580 32444
rect 6178 32416 6184 32428
rect 5552 32388 6184 32416
rect 6178 32376 6184 32388
rect 6236 32416 6242 32428
rect 7561 32419 7619 32425
rect 7561 32416 7573 32419
rect 6236 32388 7573 32416
rect 6236 32376 6242 32388
rect 7561 32385 7573 32388
rect 7607 32385 7619 32419
rect 7561 32379 7619 32385
rect 12345 32419 12403 32425
rect 12345 32385 12357 32419
rect 12391 32416 12403 32419
rect 13173 32419 13231 32425
rect 13173 32416 13185 32419
rect 12391 32388 13185 32416
rect 12391 32385 12403 32388
rect 12345 32379 12403 32385
rect 13173 32385 13185 32388
rect 13219 32385 13231 32419
rect 13173 32379 13231 32385
rect 14550 32376 14556 32428
rect 14608 32376 14614 32428
rect 15930 32376 15936 32428
rect 15988 32376 15994 32428
rect 17218 32376 17224 32428
rect 17276 32376 17282 32428
rect 5442 32308 5448 32360
rect 5500 32348 5506 32360
rect 5537 32351 5595 32357
rect 5537 32348 5549 32351
rect 5500 32320 5549 32348
rect 5500 32308 5506 32320
rect 5537 32317 5549 32320
rect 5583 32317 5595 32351
rect 5537 32311 5595 32317
rect 7466 32308 7472 32360
rect 7524 32348 7530 32360
rect 7837 32351 7895 32357
rect 7837 32348 7849 32351
rect 7524 32320 7849 32348
rect 7524 32308 7530 32320
rect 7837 32317 7849 32320
rect 7883 32317 7895 32351
rect 7837 32311 7895 32317
rect 9858 32308 9864 32360
rect 9916 32308 9922 32360
rect 11054 32308 11060 32360
rect 11112 32348 11118 32360
rect 11701 32351 11759 32357
rect 11701 32348 11713 32351
rect 11112 32320 11713 32348
rect 11112 32308 11118 32320
rect 11701 32317 11713 32320
rect 11747 32348 11759 32351
rect 12158 32348 12164 32360
rect 11747 32320 12164 32348
rect 11747 32317 11759 32320
rect 11701 32311 11759 32317
rect 12158 32308 12164 32320
rect 12216 32348 12222 32360
rect 12437 32351 12495 32357
rect 12437 32348 12449 32351
rect 12216 32320 12449 32348
rect 12216 32308 12222 32320
rect 12437 32317 12449 32320
rect 12483 32317 12495 32351
rect 12437 32311 12495 32317
rect 12529 32351 12587 32357
rect 12529 32317 12541 32351
rect 12575 32317 12587 32351
rect 12529 32311 12587 32317
rect 14829 32351 14887 32357
rect 14829 32317 14841 32351
rect 14875 32348 14887 32351
rect 16206 32348 16212 32360
rect 14875 32320 16212 32348
rect 14875 32317 14887 32320
rect 14829 32311 14887 32317
rect 11974 32240 11980 32292
rect 12032 32280 12038 32292
rect 12544 32280 12572 32311
rect 16206 32308 16212 32320
rect 16264 32308 16270 32360
rect 17497 32351 17555 32357
rect 17497 32317 17509 32351
rect 17543 32348 17555 32351
rect 17862 32348 17868 32360
rect 17543 32320 17868 32348
rect 17543 32317 17555 32320
rect 17497 32311 17555 32317
rect 17862 32308 17868 32320
rect 17920 32308 17926 32360
rect 12032 32252 12572 32280
rect 12032 32240 12038 32252
rect 16298 32240 16304 32292
rect 16356 32280 16362 32292
rect 18432 32280 18460 32447
rect 18690 32444 18696 32456
rect 18748 32444 18754 32496
rect 20272 32425 20300 32524
rect 21177 32521 21189 32555
rect 21223 32552 21235 32555
rect 21266 32552 21272 32564
rect 21223 32524 21272 32552
rect 21223 32521 21235 32524
rect 21177 32515 21235 32521
rect 21266 32512 21272 32524
rect 21324 32552 21330 32564
rect 21910 32552 21916 32564
rect 21324 32524 21916 32552
rect 21324 32512 21330 32524
rect 21910 32512 21916 32524
rect 21968 32512 21974 32564
rect 22189 32555 22247 32561
rect 22189 32521 22201 32555
rect 22235 32552 22247 32555
rect 22833 32555 22891 32561
rect 22235 32524 22784 32552
rect 22235 32521 22247 32524
rect 22189 32515 22247 32521
rect 22756 32484 22784 32524
rect 22833 32521 22845 32555
rect 22879 32552 22891 32555
rect 24486 32552 24492 32564
rect 22879 32524 24492 32552
rect 22879 32521 22891 32524
rect 22833 32515 22891 32521
rect 24486 32512 24492 32524
rect 24544 32512 24550 32564
rect 24762 32512 24768 32564
rect 24820 32552 24826 32564
rect 24857 32555 24915 32561
rect 24857 32552 24869 32555
rect 24820 32524 24869 32552
rect 24820 32512 24826 32524
rect 24857 32521 24869 32524
rect 24903 32521 24915 32555
rect 24857 32515 24915 32521
rect 24026 32484 24032 32496
rect 20364 32456 22508 32484
rect 22756 32456 24032 32484
rect 20257 32419 20315 32425
rect 20257 32385 20269 32419
rect 20303 32385 20315 32419
rect 20257 32379 20315 32385
rect 18690 32308 18696 32360
rect 18748 32308 18754 32360
rect 19518 32308 19524 32360
rect 19576 32348 19582 32360
rect 20364 32348 20392 32456
rect 21082 32376 21088 32428
rect 21140 32376 21146 32428
rect 21634 32376 21640 32428
rect 21692 32416 21698 32428
rect 22373 32419 22431 32425
rect 22373 32416 22385 32419
rect 21692 32388 22385 32416
rect 21692 32376 21698 32388
rect 22373 32385 22385 32388
rect 22419 32385 22431 32419
rect 22480 32416 22508 32456
rect 24026 32444 24032 32456
rect 24084 32444 24090 32496
rect 23017 32419 23075 32425
rect 23017 32416 23029 32419
rect 22480 32388 23029 32416
rect 22373 32379 22431 32385
rect 23017 32385 23029 32388
rect 23063 32385 23075 32419
rect 24872 32416 24900 32515
rect 25317 32419 25375 32425
rect 25317 32416 25329 32419
rect 24872 32388 25329 32416
rect 23017 32379 23075 32385
rect 25317 32385 25329 32388
rect 25363 32385 25375 32419
rect 25317 32379 25375 32385
rect 19576 32320 20392 32348
rect 21361 32351 21419 32357
rect 19576 32308 19582 32320
rect 21361 32317 21373 32351
rect 21407 32348 21419 32351
rect 21542 32348 21548 32360
rect 21407 32320 21548 32348
rect 21407 32317 21419 32320
rect 21361 32311 21419 32317
rect 21542 32308 21548 32320
rect 21600 32308 21606 32360
rect 23198 32308 23204 32360
rect 23256 32348 23262 32360
rect 23293 32351 23351 32357
rect 23293 32348 23305 32351
rect 23256 32320 23305 32348
rect 23256 32308 23262 32320
rect 23293 32317 23305 32320
rect 23339 32317 23351 32351
rect 23293 32311 23351 32317
rect 25133 32283 25191 32289
rect 25133 32280 25145 32283
rect 16356 32252 18184 32280
rect 18432 32252 25145 32280
rect 16356 32240 16362 32252
rect 10413 32215 10471 32221
rect 10413 32181 10425 32215
rect 10459 32212 10471 32215
rect 10962 32212 10968 32224
rect 10459 32184 10968 32212
rect 10459 32181 10471 32184
rect 10413 32175 10471 32181
rect 10962 32172 10968 32184
rect 11020 32172 11026 32224
rect 14550 32172 14556 32224
rect 14608 32212 14614 32224
rect 15194 32212 15200 32224
rect 14608 32184 15200 32212
rect 14608 32172 14614 32184
rect 15194 32172 15200 32184
rect 15252 32172 15258 32224
rect 16850 32172 16856 32224
rect 16908 32172 16914 32224
rect 17678 32172 17684 32224
rect 17736 32212 17742 32224
rect 18049 32215 18107 32221
rect 18049 32212 18061 32215
rect 17736 32184 18061 32212
rect 17736 32172 17742 32184
rect 18049 32181 18061 32184
rect 18095 32181 18107 32215
rect 18156 32212 18184 32252
rect 25133 32249 25145 32252
rect 25179 32249 25191 32283
rect 25133 32243 25191 32249
rect 18598 32212 18604 32224
rect 18156 32184 18604 32212
rect 18049 32175 18107 32181
rect 18598 32172 18604 32184
rect 18656 32172 18662 32224
rect 20070 32172 20076 32224
rect 20128 32172 20134 32224
rect 20717 32215 20775 32221
rect 20717 32181 20729 32215
rect 20763 32212 20775 32215
rect 21358 32212 21364 32224
rect 20763 32184 21364 32212
rect 20763 32181 20775 32184
rect 20717 32175 20775 32181
rect 21358 32172 21364 32184
rect 21416 32172 21422 32224
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 7929 32011 7987 32017
rect 7929 31977 7941 32011
rect 7975 32008 7987 32011
rect 8294 32008 8300 32020
rect 7975 31980 8300 32008
rect 7975 31977 7987 31980
rect 7929 31971 7987 31977
rect 8294 31968 8300 31980
rect 8352 31968 8358 32020
rect 9674 32017 9680 32020
rect 9664 32011 9680 32017
rect 9664 31977 9676 32011
rect 9664 31971 9680 31977
rect 9674 31968 9680 31971
rect 9732 31968 9738 32020
rect 10134 31968 10140 32020
rect 10192 32008 10198 32020
rect 10192 31980 11100 32008
rect 10192 31968 10198 31980
rect 8386 31900 8392 31952
rect 8444 31940 8450 31952
rect 11072 31940 11100 31980
rect 11146 31968 11152 32020
rect 11204 31968 11210 32020
rect 11606 31968 11612 32020
rect 11664 32008 11670 32020
rect 16393 32011 16451 32017
rect 16393 32008 16405 32011
rect 11664 31980 16405 32008
rect 11664 31968 11670 31980
rect 16393 31977 16405 31980
rect 16439 31977 16451 32011
rect 21174 32008 21180 32020
rect 16393 31971 16451 31977
rect 17052 31980 21180 32008
rect 14277 31943 14335 31949
rect 14277 31940 14289 31943
rect 8444 31912 9444 31940
rect 11072 31912 14289 31940
rect 8444 31900 8450 31912
rect 6178 31832 6184 31884
rect 6236 31832 6242 31884
rect 6457 31875 6515 31881
rect 6457 31841 6469 31875
rect 6503 31872 6515 31875
rect 6914 31872 6920 31884
rect 6503 31844 6920 31872
rect 6503 31841 6515 31844
rect 6457 31835 6515 31841
rect 6914 31832 6920 31844
rect 6972 31832 6978 31884
rect 8297 31875 8355 31881
rect 8297 31872 8309 31875
rect 7576 31844 8309 31872
rect 7576 31790 7604 31844
rect 8297 31841 8309 31844
rect 8343 31872 8355 31875
rect 8478 31872 8484 31884
rect 8343 31844 8484 31872
rect 8343 31841 8355 31844
rect 8297 31835 8355 31841
rect 8478 31832 8484 31844
rect 8536 31872 8542 31884
rect 9416 31872 9444 31912
rect 14277 31909 14289 31912
rect 14323 31909 14335 31943
rect 14277 31903 14335 31909
rect 14384 31912 16988 31940
rect 8536 31844 9352 31872
rect 9416 31844 13676 31872
rect 8536 31832 8542 31844
rect 5718 31628 5724 31680
rect 5776 31668 5782 31680
rect 8478 31668 8484 31680
rect 5776 31640 8484 31668
rect 5776 31628 5782 31640
rect 8478 31628 8484 31640
rect 8536 31628 8542 31680
rect 9324 31668 9352 31844
rect 9398 31764 9404 31816
rect 9456 31764 9462 31816
rect 11054 31764 11060 31816
rect 11112 31804 11118 31816
rect 11330 31804 11336 31816
rect 11112 31776 11336 31804
rect 11112 31764 11118 31776
rect 11330 31764 11336 31776
rect 11388 31764 11394 31816
rect 11517 31807 11575 31813
rect 11517 31773 11529 31807
rect 11563 31804 11575 31807
rect 11606 31804 11612 31816
rect 11563 31776 11612 31804
rect 11563 31773 11575 31776
rect 11517 31767 11575 31773
rect 10962 31736 10968 31748
rect 10902 31708 10968 31736
rect 10962 31696 10968 31708
rect 11020 31736 11026 31748
rect 11532 31736 11560 31767
rect 11606 31764 11612 31776
rect 11664 31804 11670 31816
rect 12066 31804 12072 31816
rect 11664 31776 12072 31804
rect 11664 31764 11670 31776
rect 12066 31764 12072 31776
rect 12124 31764 12130 31816
rect 13648 31804 13676 31844
rect 13722 31832 13728 31884
rect 13780 31872 13786 31884
rect 14384 31872 14412 31912
rect 14921 31875 14979 31881
rect 14921 31872 14933 31875
rect 13780 31844 14412 31872
rect 14476 31844 14933 31872
rect 13780 31832 13786 31844
rect 14476 31804 14504 31844
rect 14921 31841 14933 31844
rect 14967 31872 14979 31875
rect 16574 31872 16580 31884
rect 14967 31844 16580 31872
rect 14967 31841 14979 31844
rect 14921 31835 14979 31841
rect 16574 31832 16580 31844
rect 16632 31832 16638 31884
rect 16960 31881 16988 31912
rect 16945 31875 17003 31881
rect 16945 31841 16957 31875
rect 16991 31841 17003 31875
rect 16945 31835 17003 31841
rect 13648 31776 14504 31804
rect 14737 31807 14795 31813
rect 14737 31773 14749 31807
rect 14783 31804 14795 31807
rect 16853 31807 16911 31813
rect 14783 31776 16804 31804
rect 14783 31773 14795 31776
rect 14737 31767 14795 31773
rect 11020 31708 11560 31736
rect 16776 31736 16804 31776
rect 16853 31773 16865 31807
rect 16899 31804 16911 31807
rect 17052 31804 17080 31980
rect 21174 31968 21180 31980
rect 21232 31968 21238 32020
rect 24121 32011 24179 32017
rect 24121 31977 24133 32011
rect 24167 32008 24179 32011
rect 24210 32008 24216 32020
rect 24167 31980 24216 32008
rect 24167 31977 24179 31980
rect 24121 31971 24179 31977
rect 24210 31968 24216 31980
rect 24268 31968 24274 32020
rect 25130 31968 25136 32020
rect 25188 31968 25194 32020
rect 21913 31943 21971 31949
rect 19168 31912 21220 31940
rect 18414 31872 18420 31884
rect 17236 31844 18420 31872
rect 17236 31804 17264 31844
rect 18414 31832 18420 31844
rect 18472 31832 18478 31884
rect 19168 31872 19196 31912
rect 19076 31844 19196 31872
rect 18049 31807 18107 31813
rect 18049 31804 18061 31807
rect 16899 31776 17080 31804
rect 17144 31776 17264 31804
rect 18007 31776 18061 31804
rect 16899 31773 16911 31776
rect 16853 31767 16911 31773
rect 17144 31736 17172 31776
rect 18049 31773 18061 31776
rect 18095 31804 18107 31807
rect 18874 31804 18880 31816
rect 18095 31776 18880 31804
rect 18095 31773 18107 31776
rect 18049 31767 18107 31773
rect 16776 31708 17172 31736
rect 11020 31696 11026 31708
rect 17586 31696 17592 31748
rect 17644 31736 17650 31748
rect 18064 31736 18092 31767
rect 18874 31764 18880 31776
rect 18932 31764 18938 31816
rect 18966 31764 18972 31816
rect 19024 31764 19030 31816
rect 18984 31736 19012 31764
rect 17644 31708 18092 31736
rect 18800 31708 19012 31736
rect 17644 31696 17650 31708
rect 9766 31668 9772 31680
rect 9324 31640 9772 31668
rect 9766 31628 9772 31640
rect 9824 31668 9830 31680
rect 10980 31668 11008 31696
rect 18800 31680 18828 31708
rect 9824 31640 11008 31668
rect 9824 31628 9830 31640
rect 13906 31628 13912 31680
rect 13964 31668 13970 31680
rect 14645 31671 14703 31677
rect 14645 31668 14657 31671
rect 13964 31640 14657 31668
rect 13964 31628 13970 31640
rect 14645 31637 14657 31640
rect 14691 31668 14703 31671
rect 14826 31668 14832 31680
rect 14691 31640 14832 31668
rect 14691 31637 14703 31640
rect 14645 31631 14703 31637
rect 14826 31628 14832 31640
rect 14884 31628 14890 31680
rect 16758 31628 16764 31680
rect 16816 31628 16822 31680
rect 16942 31628 16948 31680
rect 17000 31668 17006 31680
rect 18782 31668 18788 31680
rect 17000 31640 18788 31668
rect 17000 31628 17006 31640
rect 18782 31628 18788 31640
rect 18840 31628 18846 31680
rect 18966 31628 18972 31680
rect 19024 31668 19030 31680
rect 19076 31668 19104 31844
rect 19610 31832 19616 31884
rect 19668 31872 19674 31884
rect 21192 31881 21220 31912
rect 21913 31909 21925 31943
rect 21959 31940 21971 31943
rect 23382 31940 23388 31952
rect 21959 31912 23388 31940
rect 21959 31909 21971 31912
rect 21913 31903 21971 31909
rect 23382 31900 23388 31912
rect 23440 31900 23446 31952
rect 19981 31875 20039 31881
rect 19981 31872 19993 31875
rect 19668 31844 19993 31872
rect 19668 31832 19674 31844
rect 19981 31841 19993 31844
rect 20027 31841 20039 31875
rect 19981 31835 20039 31841
rect 21177 31875 21235 31881
rect 21177 31841 21189 31875
rect 21223 31841 21235 31875
rect 21177 31835 21235 31841
rect 21358 31832 21364 31884
rect 21416 31872 21422 31884
rect 22373 31875 22431 31881
rect 22373 31872 22385 31875
rect 21416 31844 22385 31872
rect 21416 31832 21422 31844
rect 22373 31841 22385 31844
rect 22419 31841 22431 31875
rect 22373 31835 22431 31841
rect 22557 31875 22615 31881
rect 22557 31841 22569 31875
rect 22603 31872 22615 31875
rect 23474 31872 23480 31884
rect 22603 31844 23480 31872
rect 22603 31841 22615 31844
rect 22557 31835 22615 31841
rect 23474 31832 23480 31844
rect 23532 31832 23538 31884
rect 19889 31807 19947 31813
rect 19889 31773 19901 31807
rect 19935 31804 19947 31807
rect 20438 31804 20444 31816
rect 19935 31776 20444 31804
rect 19935 31773 19947 31776
rect 19889 31767 19947 31773
rect 20438 31764 20444 31776
rect 20496 31764 20502 31816
rect 21085 31807 21143 31813
rect 21085 31773 21097 31807
rect 21131 31804 21143 31807
rect 21818 31804 21824 31816
rect 21131 31776 21824 31804
rect 21131 31773 21143 31776
rect 21085 31767 21143 31773
rect 21818 31764 21824 31776
rect 21876 31764 21882 31816
rect 24857 31807 24915 31813
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 25314 31804 25320 31816
rect 24903 31776 25320 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 19797 31739 19855 31745
rect 19797 31705 19809 31739
rect 19843 31736 19855 31739
rect 20530 31736 20536 31748
rect 19843 31708 20536 31736
rect 19843 31705 19855 31708
rect 19797 31699 19855 31705
rect 20530 31696 20536 31708
rect 20588 31696 20594 31748
rect 20993 31739 21051 31745
rect 20993 31705 21005 31739
rect 21039 31736 21051 31739
rect 21174 31736 21180 31748
rect 21039 31708 21180 31736
rect 21039 31705 21051 31708
rect 20993 31699 21051 31705
rect 21174 31696 21180 31708
rect 21232 31696 21238 31748
rect 19024 31640 19104 31668
rect 19024 31628 19030 31640
rect 19150 31628 19156 31680
rect 19208 31668 19214 31680
rect 19429 31671 19487 31677
rect 19429 31668 19441 31671
rect 19208 31640 19441 31668
rect 19208 31628 19214 31640
rect 19429 31637 19441 31640
rect 19475 31637 19487 31671
rect 19429 31631 19487 31637
rect 20622 31628 20628 31680
rect 20680 31628 20686 31680
rect 20898 31628 20904 31680
rect 20956 31668 20962 31680
rect 22281 31671 22339 31677
rect 22281 31668 22293 31671
rect 20956 31640 22293 31668
rect 20956 31628 20962 31640
rect 22281 31637 22293 31640
rect 22327 31637 22339 31671
rect 22281 31631 22339 31637
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 7469 31467 7527 31473
rect 7469 31433 7481 31467
rect 7515 31464 7527 31467
rect 7650 31464 7656 31476
rect 7515 31436 7656 31464
rect 7515 31433 7527 31436
rect 7469 31427 7527 31433
rect 7650 31424 7656 31436
rect 7708 31424 7714 31476
rect 8662 31424 8668 31476
rect 8720 31424 8726 31476
rect 9033 31467 9091 31473
rect 9033 31433 9045 31467
rect 9079 31464 9091 31467
rect 9858 31464 9864 31476
rect 9079 31436 9864 31464
rect 9079 31433 9091 31436
rect 9033 31427 9091 31433
rect 9858 31424 9864 31436
rect 9916 31424 9922 31476
rect 13354 31424 13360 31476
rect 13412 31464 13418 31476
rect 13538 31464 13544 31476
rect 13412 31436 13544 31464
rect 13412 31424 13418 31436
rect 13538 31424 13544 31436
rect 13596 31424 13602 31476
rect 15013 31467 15071 31473
rect 15013 31433 15025 31467
rect 15059 31464 15071 31467
rect 15930 31464 15936 31476
rect 15059 31436 15936 31464
rect 15059 31433 15071 31436
rect 15013 31427 15071 31433
rect 8386 31356 8392 31408
rect 8444 31396 8450 31408
rect 15028 31396 15056 31427
rect 15930 31424 15936 31436
rect 15988 31424 15994 31476
rect 17586 31424 17592 31476
rect 17644 31424 17650 31476
rect 18325 31467 18383 31473
rect 18325 31433 18337 31467
rect 18371 31464 18383 31467
rect 18506 31464 18512 31476
rect 18371 31436 18512 31464
rect 18371 31433 18383 31436
rect 18325 31427 18383 31433
rect 18506 31424 18512 31436
rect 18564 31424 18570 31476
rect 19521 31467 19579 31473
rect 19521 31433 19533 31467
rect 19567 31464 19579 31467
rect 21450 31464 21456 31476
rect 19567 31436 21456 31464
rect 19567 31433 19579 31436
rect 19521 31427 19579 31433
rect 21450 31424 21456 31436
rect 21508 31424 21514 31476
rect 21545 31467 21603 31473
rect 21545 31433 21557 31467
rect 21591 31464 21603 31467
rect 21818 31464 21824 31476
rect 21591 31436 21824 31464
rect 21591 31433 21603 31436
rect 21545 31427 21603 31433
rect 21818 31424 21824 31436
rect 21876 31424 21882 31476
rect 23290 31424 23296 31476
rect 23348 31464 23354 31476
rect 23348 31436 24348 31464
rect 23348 31424 23354 31436
rect 8444 31368 9260 31396
rect 14398 31368 15056 31396
rect 8444 31356 8450 31368
rect 1765 31331 1823 31337
rect 1765 31297 1777 31331
rect 1811 31328 1823 31331
rect 1946 31328 1952 31340
rect 1811 31300 1952 31328
rect 1811 31297 1823 31300
rect 1765 31291 1823 31297
rect 1946 31288 1952 31300
rect 2004 31288 2010 31340
rect 7834 31288 7840 31340
rect 7892 31288 7898 31340
rect 7929 31331 7987 31337
rect 7929 31297 7941 31331
rect 7975 31328 7987 31331
rect 8938 31328 8944 31340
rect 7975 31300 8944 31328
rect 7975 31297 7987 31300
rect 7929 31291 7987 31297
rect 1302 31220 1308 31272
rect 1360 31260 1366 31272
rect 2041 31263 2099 31269
rect 2041 31260 2053 31263
rect 1360 31232 2053 31260
rect 1360 31220 1366 31232
rect 2041 31229 2053 31232
rect 2087 31229 2099 31263
rect 2041 31223 2099 31229
rect 5626 31220 5632 31272
rect 5684 31260 5690 31272
rect 7193 31263 7251 31269
rect 7193 31260 7205 31263
rect 5684 31232 7205 31260
rect 5684 31220 5690 31232
rect 7193 31229 7205 31232
rect 7239 31260 7251 31263
rect 7944 31260 7972 31291
rect 8938 31288 8944 31300
rect 8996 31288 9002 31340
rect 7239 31232 7972 31260
rect 7239 31229 7251 31232
rect 7193 31223 7251 31229
rect 8110 31220 8116 31272
rect 8168 31220 8174 31272
rect 8478 31220 8484 31272
rect 8536 31260 8542 31272
rect 9232 31269 9260 31368
rect 15102 31356 15108 31408
rect 15160 31396 15166 31408
rect 15160 31368 18920 31396
rect 15160 31356 15166 31368
rect 17497 31331 17555 31337
rect 17497 31297 17509 31331
rect 17543 31297 17555 31331
rect 17497 31291 17555 31297
rect 9125 31263 9183 31269
rect 9125 31260 9137 31263
rect 8536 31232 9137 31260
rect 8536 31220 8542 31232
rect 9125 31229 9137 31232
rect 9171 31229 9183 31263
rect 9125 31223 9183 31229
rect 9217 31263 9275 31269
rect 9217 31229 9229 31263
rect 9263 31229 9275 31263
rect 9217 31223 9275 31229
rect 9398 31220 9404 31272
rect 9456 31260 9462 31272
rect 12897 31263 12955 31269
rect 12897 31260 12909 31263
rect 9456 31232 12909 31260
rect 9456 31220 9462 31232
rect 12897 31229 12909 31232
rect 12943 31260 12955 31263
rect 13173 31263 13231 31269
rect 12943 31232 13032 31260
rect 12943 31229 12955 31232
rect 12897 31223 12955 31229
rect 7374 31152 7380 31204
rect 7432 31192 7438 31204
rect 8128 31192 8156 31220
rect 7432 31164 8156 31192
rect 7432 31152 7438 31164
rect 13004 31124 13032 31232
rect 13173 31229 13185 31263
rect 13219 31260 13231 31263
rect 13262 31260 13268 31272
rect 13219 31232 13268 31260
rect 13219 31229 13231 31232
rect 13173 31223 13231 31229
rect 13262 31220 13268 31232
rect 13320 31220 13326 31272
rect 14366 31220 14372 31272
rect 14424 31260 14430 31272
rect 16761 31263 16819 31269
rect 16761 31260 16773 31263
rect 14424 31232 16773 31260
rect 14424 31220 14430 31232
rect 16761 31229 16773 31232
rect 16807 31260 16819 31263
rect 17512 31260 17540 31291
rect 18322 31288 18328 31340
rect 18380 31328 18386 31340
rect 18693 31331 18751 31337
rect 18693 31328 18705 31331
rect 18380 31300 18705 31328
rect 18380 31288 18386 31300
rect 18693 31297 18705 31300
rect 18739 31297 18751 31331
rect 18693 31291 18751 31297
rect 16807 31232 17540 31260
rect 16807 31229 16819 31232
rect 16761 31223 16819 31229
rect 17770 31220 17776 31272
rect 17828 31220 17834 31272
rect 18892 31269 18920 31368
rect 19886 31356 19892 31408
rect 19944 31356 19950 31408
rect 21634 31356 21640 31408
rect 21692 31396 21698 31408
rect 22465 31399 22523 31405
rect 22465 31396 22477 31399
rect 21692 31368 22477 31396
rect 21692 31356 21698 31368
rect 22465 31365 22477 31368
rect 22511 31365 22523 31399
rect 24210 31396 24216 31408
rect 23690 31368 24216 31396
rect 22465 31359 22523 31365
rect 24210 31356 24216 31368
rect 24268 31356 24274 31408
rect 20717 31331 20775 31337
rect 20717 31328 20729 31331
rect 19996 31300 20729 31328
rect 19996 31272 20024 31300
rect 20717 31297 20729 31300
rect 20763 31297 20775 31331
rect 24320 31328 24348 31436
rect 24394 31424 24400 31476
rect 24452 31464 24458 31476
rect 25133 31467 25191 31473
rect 25133 31464 25145 31467
rect 24452 31436 25145 31464
rect 24452 31424 24458 31436
rect 25133 31433 25145 31436
rect 25179 31433 25191 31467
rect 25133 31427 25191 31433
rect 24581 31331 24639 31337
rect 24581 31328 24593 31331
rect 24320 31300 24593 31328
rect 20717 31291 20775 31297
rect 24581 31297 24593 31300
rect 24627 31297 24639 31331
rect 24581 31291 24639 31297
rect 25314 31288 25320 31340
rect 25372 31288 25378 31340
rect 18785 31263 18843 31269
rect 18785 31229 18797 31263
rect 18831 31229 18843 31263
rect 18785 31223 18843 31229
rect 18877 31263 18935 31269
rect 18877 31229 18889 31263
rect 18923 31229 18935 31263
rect 18877 31223 18935 31229
rect 16482 31152 16488 31204
rect 16540 31192 16546 31204
rect 18800 31192 18828 31223
rect 19058 31220 19064 31272
rect 19116 31260 19122 31272
rect 19978 31260 19984 31272
rect 19116 31232 19984 31260
rect 19116 31220 19122 31232
rect 19978 31220 19984 31232
rect 20036 31220 20042 31272
rect 20165 31263 20223 31269
rect 20165 31229 20177 31263
rect 20211 31260 20223 31263
rect 20530 31260 20536 31272
rect 20211 31232 20536 31260
rect 20211 31229 20223 31232
rect 20165 31223 20223 31229
rect 20530 31220 20536 31232
rect 20588 31260 20594 31272
rect 22094 31260 22100 31272
rect 20588 31232 22100 31260
rect 20588 31220 20594 31232
rect 22094 31220 22100 31232
rect 22152 31220 22158 31272
rect 22186 31220 22192 31272
rect 22244 31220 22250 31272
rect 24946 31260 24952 31272
rect 22296 31232 24952 31260
rect 22296 31192 22324 31232
rect 24946 31220 24952 31232
rect 25004 31220 25010 31272
rect 16540 31164 18644 31192
rect 18800 31164 22324 31192
rect 16540 31152 16546 31164
rect 14458 31124 14464 31136
rect 13004 31096 14464 31124
rect 14458 31084 14464 31096
rect 14516 31084 14522 31136
rect 14642 31084 14648 31136
rect 14700 31084 14706 31136
rect 17126 31084 17132 31136
rect 17184 31084 17190 31136
rect 18616 31124 18644 31164
rect 22296 31136 22324 31164
rect 19886 31124 19892 31136
rect 18616 31096 19892 31124
rect 19886 31084 19892 31096
rect 19944 31124 19950 31136
rect 20533 31127 20591 31133
rect 20533 31124 20545 31127
rect 19944 31096 20545 31124
rect 19944 31084 19950 31096
rect 20533 31093 20545 31096
rect 20579 31093 20591 31127
rect 20533 31087 20591 31093
rect 22278 31084 22284 31136
rect 22336 31084 22342 31136
rect 23566 31084 23572 31136
rect 23624 31124 23630 31136
rect 23937 31127 23995 31133
rect 23937 31124 23949 31127
rect 23624 31096 23949 31124
rect 23624 31084 23630 31096
rect 23937 31093 23949 31096
rect 23983 31093 23995 31127
rect 23937 31087 23995 31093
rect 24394 31084 24400 31136
rect 24452 31084 24458 31136
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 8110 30880 8116 30932
rect 8168 30920 8174 30932
rect 8168 30892 12434 30920
rect 8168 30880 8174 30892
rect 11606 30852 11612 30864
rect 10980 30824 11612 30852
rect 1578 30744 1584 30796
rect 1636 30784 1642 30796
rect 3973 30787 4031 30793
rect 3973 30784 3985 30787
rect 1636 30756 3985 30784
rect 1636 30744 1642 30756
rect 3973 30753 3985 30756
rect 4019 30753 4031 30787
rect 3973 30747 4031 30753
rect 7834 30744 7840 30796
rect 7892 30784 7898 30796
rect 7929 30787 7987 30793
rect 7929 30784 7941 30787
rect 7892 30756 7941 30784
rect 7892 30744 7898 30756
rect 7929 30753 7941 30756
rect 7975 30753 7987 30787
rect 7929 30747 7987 30753
rect 9398 30744 9404 30796
rect 9456 30784 9462 30796
rect 9585 30787 9643 30793
rect 9585 30784 9597 30787
rect 9456 30756 9597 30784
rect 9456 30744 9462 30756
rect 9585 30753 9597 30756
rect 9631 30753 9643 30787
rect 9585 30747 9643 30753
rect 9861 30787 9919 30793
rect 9861 30753 9873 30787
rect 9907 30784 9919 30787
rect 10594 30784 10600 30796
rect 9907 30756 10600 30784
rect 9907 30753 9919 30756
rect 9861 30747 9919 30753
rect 10594 30744 10600 30756
rect 10652 30744 10658 30796
rect 10980 30702 11008 30824
rect 11606 30812 11612 30824
rect 11664 30812 11670 30864
rect 12406 30784 12434 30892
rect 12526 30880 12532 30932
rect 12584 30920 12590 30932
rect 12805 30923 12863 30929
rect 12805 30920 12817 30923
rect 12584 30892 12817 30920
rect 12584 30880 12590 30892
rect 12805 30889 12817 30892
rect 12851 30889 12863 30923
rect 12805 30883 12863 30889
rect 15930 30880 15936 30932
rect 15988 30920 15994 30932
rect 18233 30923 18291 30929
rect 18233 30920 18245 30923
rect 15988 30892 18245 30920
rect 15988 30880 15994 30892
rect 13357 30787 13415 30793
rect 13357 30784 13369 30787
rect 12406 30756 13369 30784
rect 13357 30753 13369 30756
rect 13403 30753 13415 30787
rect 13357 30747 13415 30753
rect 15194 30744 15200 30796
rect 15252 30784 15258 30796
rect 16209 30787 16267 30793
rect 16209 30784 16221 30787
rect 15252 30756 16221 30784
rect 15252 30744 15258 30756
rect 16209 30753 16221 30756
rect 16255 30753 16267 30787
rect 16209 30747 16267 30753
rect 16485 30787 16543 30793
rect 16485 30753 16497 30787
rect 16531 30784 16543 30787
rect 16942 30784 16948 30796
rect 16531 30756 16948 30784
rect 16531 30753 16543 30756
rect 16485 30747 16543 30753
rect 16942 30744 16948 30756
rect 17000 30744 17006 30796
rect 11238 30676 11244 30728
rect 11296 30716 11302 30728
rect 12529 30719 12587 30725
rect 12529 30716 12541 30719
rect 11296 30688 12541 30716
rect 11296 30676 11302 30688
rect 12529 30685 12541 30688
rect 12575 30716 12587 30719
rect 13173 30719 13231 30725
rect 13173 30716 13185 30719
rect 12575 30688 13185 30716
rect 12575 30685 12587 30688
rect 12529 30679 12587 30685
rect 13173 30685 13185 30688
rect 13219 30716 13231 30719
rect 13538 30716 13544 30728
rect 13219 30688 13544 30716
rect 13219 30685 13231 30688
rect 13173 30679 13231 30685
rect 13538 30676 13544 30688
rect 13596 30676 13602 30728
rect 17604 30702 17632 30892
rect 18233 30889 18245 30892
rect 18279 30889 18291 30923
rect 18233 30883 18291 30889
rect 18598 30880 18604 30932
rect 18656 30920 18662 30932
rect 19242 30920 19248 30932
rect 18656 30892 19248 30920
rect 18656 30880 18662 30892
rect 19242 30880 19248 30892
rect 19300 30880 19306 30932
rect 20438 30920 20444 30932
rect 19904 30892 20444 30920
rect 19904 30793 19932 30892
rect 20438 30880 20444 30892
rect 20496 30880 20502 30932
rect 23109 30923 23167 30929
rect 23109 30889 23121 30923
rect 23155 30920 23167 30923
rect 23474 30920 23480 30932
rect 23155 30892 23480 30920
rect 23155 30889 23167 30892
rect 23109 30883 23167 30889
rect 23474 30880 23480 30892
rect 23532 30920 23538 30932
rect 23842 30920 23848 30932
rect 23532 30892 23848 30920
rect 23532 30880 23538 30892
rect 23842 30880 23848 30892
rect 23900 30880 23906 30932
rect 24857 30923 24915 30929
rect 24857 30889 24869 30923
rect 24903 30920 24915 30923
rect 25314 30920 25320 30932
rect 24903 30892 25320 30920
rect 24903 30889 24915 30892
rect 24857 30883 24915 30889
rect 25314 30880 25320 30892
rect 25372 30880 25378 30932
rect 19889 30787 19947 30793
rect 19889 30753 19901 30787
rect 19935 30753 19947 30787
rect 19889 30747 19947 30753
rect 19978 30744 19984 30796
rect 20036 30744 20042 30796
rect 20162 30744 20168 30796
rect 20220 30784 20226 30796
rect 22557 30787 22615 30793
rect 22557 30784 22569 30787
rect 20220 30756 22569 30784
rect 20220 30744 20226 30756
rect 22557 30753 22569 30756
rect 22603 30753 22615 30787
rect 22557 30747 22615 30753
rect 19797 30719 19855 30725
rect 19797 30685 19809 30719
rect 19843 30716 19855 30719
rect 20254 30716 20260 30728
rect 19843 30688 20260 30716
rect 19843 30685 19855 30688
rect 19797 30679 19855 30685
rect 20254 30676 20260 30688
rect 20312 30676 20318 30728
rect 22278 30676 22284 30728
rect 22336 30716 22342 30728
rect 22373 30719 22431 30725
rect 22373 30716 22385 30719
rect 22336 30688 22385 30716
rect 22336 30676 22342 30688
rect 22373 30685 22385 30688
rect 22419 30685 22431 30719
rect 22373 30679 22431 30685
rect 22462 30676 22468 30728
rect 22520 30716 22526 30728
rect 23845 30719 23903 30725
rect 23845 30716 23857 30719
rect 22520 30688 23857 30716
rect 22520 30676 22526 30688
rect 23845 30685 23857 30688
rect 23891 30685 23903 30719
rect 23845 30679 23903 30685
rect 25317 30719 25375 30725
rect 25317 30685 25329 30719
rect 25363 30716 25375 30719
rect 25498 30716 25504 30728
rect 25363 30688 25504 30716
rect 25363 30685 25375 30688
rect 25317 30679 25375 30685
rect 25498 30676 25504 30688
rect 25556 30676 25562 30728
rect 3786 30608 3792 30660
rect 3844 30648 3850 30660
rect 4157 30651 4215 30657
rect 4157 30648 4169 30651
rect 3844 30620 4169 30648
rect 3844 30608 3850 30620
rect 4157 30617 4169 30620
rect 4203 30617 4215 30651
rect 4157 30611 4215 30617
rect 5813 30651 5871 30657
rect 5813 30617 5825 30651
rect 5859 30648 5871 30651
rect 6270 30648 6276 30660
rect 5859 30620 6276 30648
rect 5859 30617 5871 30620
rect 5813 30611 5871 30617
rect 6270 30608 6276 30620
rect 6328 30608 6334 30660
rect 13265 30651 13323 30657
rect 13265 30617 13277 30651
rect 13311 30648 13323 30651
rect 16574 30648 16580 30660
rect 13311 30620 16580 30648
rect 13311 30617 13323 30620
rect 13265 30611 13323 30617
rect 16574 30608 16580 30620
rect 16632 30608 16638 30660
rect 18506 30608 18512 30660
rect 18564 30648 18570 30660
rect 18690 30648 18696 30660
rect 18564 30620 18696 30648
rect 18564 30608 18570 30620
rect 18690 30608 18696 30620
rect 18748 30608 18754 30660
rect 8478 30540 8484 30592
rect 8536 30540 8542 30592
rect 11330 30540 11336 30592
rect 11388 30540 11394 30592
rect 17862 30540 17868 30592
rect 17920 30580 17926 30592
rect 17957 30583 18015 30589
rect 17957 30580 17969 30583
rect 17920 30552 17969 30580
rect 17920 30540 17926 30552
rect 17957 30549 17969 30552
rect 18003 30549 18015 30583
rect 17957 30543 18015 30549
rect 19426 30540 19432 30592
rect 19484 30540 19490 30592
rect 22005 30583 22063 30589
rect 22005 30549 22017 30583
rect 22051 30580 22063 30583
rect 22278 30580 22284 30592
rect 22051 30552 22284 30580
rect 22051 30549 22063 30552
rect 22005 30543 22063 30549
rect 22278 30540 22284 30552
rect 22336 30540 22342 30592
rect 22465 30583 22523 30589
rect 22465 30549 22477 30583
rect 22511 30580 22523 30583
rect 23474 30580 23480 30592
rect 22511 30552 23480 30580
rect 22511 30549 22523 30552
rect 22465 30543 22523 30549
rect 23474 30540 23480 30552
rect 23532 30540 23538 30592
rect 23661 30583 23719 30589
rect 23661 30549 23673 30583
rect 23707 30580 23719 30583
rect 25038 30580 25044 30592
rect 23707 30552 25044 30580
rect 23707 30549 23719 30552
rect 23661 30543 23719 30549
rect 25038 30540 25044 30552
rect 25096 30540 25102 30592
rect 25130 30540 25136 30592
rect 25188 30540 25194 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 11790 30336 11796 30388
rect 11848 30376 11854 30388
rect 12529 30379 12587 30385
rect 12529 30376 12541 30379
rect 11848 30348 12541 30376
rect 11848 30336 11854 30348
rect 12529 30345 12541 30348
rect 12575 30376 12587 30379
rect 16942 30376 16948 30388
rect 12575 30348 16948 30376
rect 12575 30345 12587 30348
rect 12529 30339 12587 30345
rect 16942 30336 16948 30348
rect 17000 30336 17006 30388
rect 18322 30336 18328 30388
rect 18380 30376 18386 30388
rect 18690 30376 18696 30388
rect 18380 30348 18696 30376
rect 18380 30336 18386 30348
rect 18690 30336 18696 30348
rect 18748 30336 18754 30388
rect 20438 30336 20444 30388
rect 20496 30376 20502 30388
rect 25130 30376 25136 30388
rect 20496 30348 25136 30376
rect 20496 30336 20502 30348
rect 25130 30336 25136 30348
rect 25188 30336 25194 30388
rect 8386 30268 8392 30320
rect 8444 30308 8450 30320
rect 11238 30308 11244 30320
rect 8444 30280 11244 30308
rect 8444 30268 8450 30280
rect 11238 30268 11244 30280
rect 11296 30268 11302 30320
rect 16390 30268 16396 30320
rect 16448 30308 16454 30320
rect 16448 30280 19656 30308
rect 16448 30268 16454 30280
rect 10781 30243 10839 30249
rect 10781 30209 10793 30243
rect 10827 30240 10839 30243
rect 11701 30243 11759 30249
rect 11701 30240 11713 30243
rect 10827 30212 11713 30240
rect 10827 30209 10839 30212
rect 10781 30203 10839 30209
rect 11701 30209 11713 30212
rect 11747 30209 11759 30243
rect 14366 30240 14372 30252
rect 11701 30203 11759 30209
rect 12406 30212 14372 30240
rect 10042 30132 10048 30184
rect 10100 30172 10106 30184
rect 10137 30175 10195 30181
rect 10137 30172 10149 30175
rect 10100 30144 10149 30172
rect 10100 30132 10106 30144
rect 10137 30141 10149 30144
rect 10183 30172 10195 30175
rect 10594 30172 10600 30184
rect 10183 30144 10600 30172
rect 10183 30141 10195 30144
rect 10137 30135 10195 30141
rect 10594 30132 10600 30144
rect 10652 30172 10658 30184
rect 10873 30175 10931 30181
rect 10873 30172 10885 30175
rect 10652 30144 10885 30172
rect 10652 30132 10658 30144
rect 10873 30141 10885 30144
rect 10919 30141 10931 30175
rect 10873 30135 10931 30141
rect 10965 30175 11023 30181
rect 10965 30141 10977 30175
rect 11011 30141 11023 30175
rect 10965 30135 11023 30141
rect 10686 30064 10692 30116
rect 10744 30104 10750 30116
rect 10980 30104 11008 30135
rect 10744 30076 11008 30104
rect 10744 30064 10750 30076
rect 10410 29996 10416 30048
rect 10468 29996 10474 30048
rect 11882 29996 11888 30048
rect 11940 30036 11946 30048
rect 12253 30039 12311 30045
rect 12253 30036 12265 30039
rect 11940 30008 12265 30036
rect 11940 29996 11946 30008
rect 12253 30005 12265 30008
rect 12299 30036 12311 30039
rect 12406 30036 12434 30212
rect 14366 30200 14372 30212
rect 14424 30200 14430 30252
rect 14458 30200 14464 30252
rect 14516 30200 14522 30252
rect 15838 30200 15844 30252
rect 15896 30200 15902 30252
rect 17402 30240 17408 30252
rect 16132 30212 17408 30240
rect 14737 30175 14795 30181
rect 14737 30141 14749 30175
rect 14783 30172 14795 30175
rect 16132 30172 16160 30212
rect 17402 30200 17408 30212
rect 17460 30240 17466 30252
rect 17862 30240 17868 30252
rect 17460 30212 17868 30240
rect 17460 30200 17466 30212
rect 17862 30200 17868 30212
rect 17920 30200 17926 30252
rect 17957 30243 18015 30249
rect 17957 30209 17969 30243
rect 18003 30240 18015 30243
rect 18601 30243 18659 30249
rect 18601 30240 18613 30243
rect 18003 30212 18613 30240
rect 18003 30209 18015 30212
rect 17957 30203 18015 30209
rect 18601 30209 18613 30212
rect 18647 30209 18659 30243
rect 18601 30203 18659 30209
rect 18877 30243 18935 30249
rect 18877 30209 18889 30243
rect 18923 30240 18935 30243
rect 19058 30240 19064 30252
rect 18923 30212 19064 30240
rect 18923 30209 18935 30212
rect 18877 30203 18935 30209
rect 14783 30144 16160 30172
rect 14783 30141 14795 30144
rect 14737 30135 14795 30141
rect 16206 30132 16212 30184
rect 16264 30132 16270 30184
rect 16945 30175 17003 30181
rect 16945 30141 16957 30175
rect 16991 30172 17003 30175
rect 17218 30172 17224 30184
rect 16991 30144 17224 30172
rect 16991 30141 17003 30144
rect 16945 30135 17003 30141
rect 17218 30132 17224 30144
rect 17276 30132 17282 30184
rect 17972 30104 18000 30203
rect 19058 30200 19064 30212
rect 19116 30200 19122 30252
rect 19628 30249 19656 30280
rect 23566 30268 23572 30320
rect 23624 30308 23630 30320
rect 23661 30311 23719 30317
rect 23661 30308 23673 30311
rect 23624 30280 23673 30308
rect 23624 30268 23630 30280
rect 23661 30277 23673 30280
rect 23707 30277 23719 30311
rect 23661 30271 23719 30277
rect 24210 30268 24216 30320
rect 24268 30268 24274 30320
rect 19613 30243 19671 30249
rect 19613 30209 19625 30243
rect 19659 30209 19671 30243
rect 19613 30203 19671 30209
rect 22186 30200 22192 30252
rect 22244 30240 22250 30252
rect 23385 30243 23443 30249
rect 23385 30240 23397 30243
rect 22244 30212 23397 30240
rect 22244 30200 22250 30212
rect 23385 30209 23397 30212
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 18049 30175 18107 30181
rect 18049 30141 18061 30175
rect 18095 30141 18107 30175
rect 18049 30135 18107 30141
rect 18233 30175 18291 30181
rect 18233 30141 18245 30175
rect 18279 30172 18291 30175
rect 19794 30172 19800 30184
rect 18279 30144 19800 30172
rect 18279 30141 18291 30144
rect 18233 30135 18291 30141
rect 17512 30076 18000 30104
rect 12299 30008 12434 30036
rect 12299 30005 12311 30008
rect 12253 29999 12311 30005
rect 14366 29996 14372 30048
rect 14424 30036 14430 30048
rect 17512 30036 17540 30076
rect 14424 30008 17540 30036
rect 14424 29996 14430 30008
rect 17586 29996 17592 30048
rect 17644 29996 17650 30048
rect 18064 30036 18092 30135
rect 19794 30132 19800 30144
rect 19852 30132 19858 30184
rect 23750 30132 23756 30184
rect 23808 30172 23814 30184
rect 25133 30175 25191 30181
rect 25133 30172 25145 30175
rect 23808 30144 25145 30172
rect 23808 30132 23814 30144
rect 25133 30141 25145 30144
rect 25179 30141 25191 30175
rect 25133 30135 25191 30141
rect 18322 30064 18328 30116
rect 18380 30104 18386 30116
rect 21082 30104 21088 30116
rect 18380 30076 21088 30104
rect 18380 30064 18386 30076
rect 21082 30064 21088 30076
rect 21140 30064 21146 30116
rect 19058 30036 19064 30048
rect 18064 30008 19064 30036
rect 19058 29996 19064 30008
rect 19116 30036 19122 30048
rect 19242 30036 19248 30048
rect 19116 30008 19248 30036
rect 19116 29996 19122 30008
rect 19242 29996 19248 30008
rect 19300 29996 19306 30048
rect 19429 30039 19487 30045
rect 19429 30005 19441 30039
rect 19475 30036 19487 30039
rect 21818 30036 21824 30048
rect 19475 30008 21824 30036
rect 19475 30005 19487 30008
rect 19429 29999 19487 30005
rect 21818 29996 21824 30008
rect 21876 29996 21882 30048
rect 24210 29996 24216 30048
rect 24268 30036 24274 30048
rect 25409 30039 25467 30045
rect 25409 30036 25421 30039
rect 24268 30008 25421 30036
rect 24268 29996 24274 30008
rect 25409 30005 25421 30008
rect 25455 30005 25467 30039
rect 25409 29999 25467 30005
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 4246 29792 4252 29844
rect 4304 29832 4310 29844
rect 7285 29835 7343 29841
rect 7285 29832 7297 29835
rect 4304 29804 7297 29832
rect 4304 29792 4310 29804
rect 7285 29801 7297 29804
rect 7331 29832 7343 29835
rect 7650 29832 7656 29844
rect 7331 29804 7656 29832
rect 7331 29801 7343 29804
rect 7285 29795 7343 29801
rect 7650 29792 7656 29804
rect 7708 29792 7714 29844
rect 7742 29792 7748 29844
rect 7800 29832 7806 29844
rect 7837 29835 7895 29841
rect 7837 29832 7849 29835
rect 7800 29804 7849 29832
rect 7800 29792 7806 29804
rect 7837 29801 7849 29804
rect 7883 29801 7895 29835
rect 7837 29795 7895 29801
rect 9490 29792 9496 29844
rect 9548 29792 9554 29844
rect 10410 29792 10416 29844
rect 10468 29832 10474 29844
rect 12986 29832 12992 29844
rect 10468 29804 12992 29832
rect 10468 29792 10474 29804
rect 12986 29792 12992 29804
rect 13044 29792 13050 29844
rect 16022 29792 16028 29844
rect 16080 29832 16086 29844
rect 16482 29832 16488 29844
rect 16080 29804 16488 29832
rect 16080 29792 16086 29804
rect 16482 29792 16488 29804
rect 16540 29792 16546 29844
rect 16574 29792 16580 29844
rect 16632 29832 16638 29844
rect 21726 29832 21732 29844
rect 16632 29804 21732 29832
rect 16632 29792 16638 29804
rect 21726 29792 21732 29804
rect 21784 29792 21790 29844
rect 6362 29724 6368 29776
rect 6420 29764 6426 29776
rect 8941 29767 8999 29773
rect 8941 29764 8953 29767
rect 6420 29736 8953 29764
rect 6420 29724 6426 29736
rect 8941 29733 8953 29736
rect 8987 29764 8999 29767
rect 9306 29764 9312 29776
rect 8987 29736 9312 29764
rect 8987 29733 8999 29736
rect 8941 29727 8999 29733
rect 9306 29724 9312 29736
rect 9364 29764 9370 29776
rect 9582 29764 9588 29776
rect 9364 29736 9588 29764
rect 9364 29724 9370 29736
rect 9582 29724 9588 29736
rect 9640 29724 9646 29776
rect 11330 29724 11336 29776
rect 11388 29764 11394 29776
rect 12621 29767 12679 29773
rect 11388 29736 12434 29764
rect 11388 29724 11394 29736
rect 4062 29656 4068 29708
rect 4120 29696 4126 29708
rect 4249 29699 4307 29705
rect 4249 29696 4261 29699
rect 4120 29668 4261 29696
rect 4120 29656 4126 29668
rect 4249 29665 4261 29668
rect 4295 29665 4307 29699
rect 4249 29659 4307 29665
rect 6914 29656 6920 29708
rect 6972 29696 6978 29708
rect 8389 29699 8447 29705
rect 8389 29696 8401 29699
rect 6972 29668 8401 29696
rect 6972 29656 6978 29668
rect 8389 29665 8401 29668
rect 8435 29665 8447 29699
rect 8389 29659 8447 29665
rect 9674 29656 9680 29708
rect 9732 29696 9738 29708
rect 10045 29699 10103 29705
rect 10045 29696 10057 29699
rect 9732 29668 10057 29696
rect 9732 29656 9738 29668
rect 10045 29665 10057 29668
rect 10091 29665 10103 29699
rect 11977 29699 12035 29705
rect 11977 29696 11989 29699
rect 10045 29659 10103 29665
rect 10152 29668 11989 29696
rect 7834 29588 7840 29640
rect 7892 29628 7898 29640
rect 10152 29628 10180 29668
rect 11977 29665 11989 29668
rect 12023 29665 12035 29699
rect 12406 29696 12434 29736
rect 12621 29733 12633 29767
rect 12667 29764 12679 29767
rect 17310 29764 17316 29776
rect 12667 29736 17316 29764
rect 12667 29733 12679 29736
rect 12621 29727 12679 29733
rect 17310 29724 17316 29736
rect 17368 29724 17374 29776
rect 17586 29724 17592 29776
rect 17644 29764 17650 29776
rect 25133 29767 25191 29773
rect 25133 29764 25145 29767
rect 17644 29736 20116 29764
rect 17644 29724 17650 29736
rect 13173 29699 13231 29705
rect 13173 29696 13185 29699
rect 12406 29668 13185 29696
rect 11977 29659 12035 29665
rect 13173 29665 13185 29668
rect 13219 29665 13231 29699
rect 13173 29659 13231 29665
rect 14918 29656 14924 29708
rect 14976 29696 14982 29708
rect 17497 29699 17555 29705
rect 17497 29696 17509 29699
rect 14976 29668 17509 29696
rect 14976 29656 14982 29668
rect 17497 29665 17509 29668
rect 17543 29665 17555 29699
rect 17497 29659 17555 29665
rect 18782 29656 18788 29708
rect 18840 29656 18846 29708
rect 20088 29705 20116 29736
rect 21284 29736 25145 29764
rect 20073 29699 20131 29705
rect 20073 29665 20085 29699
rect 20119 29665 20131 29699
rect 20073 29659 20131 29665
rect 20257 29699 20315 29705
rect 20257 29665 20269 29699
rect 20303 29696 20315 29699
rect 21174 29696 21180 29708
rect 20303 29668 21180 29696
rect 20303 29665 20315 29668
rect 20257 29659 20315 29665
rect 21174 29656 21180 29668
rect 21232 29656 21238 29708
rect 7892 29600 10180 29628
rect 7892 29588 7898 29600
rect 11790 29588 11796 29640
rect 11848 29588 11854 29640
rect 12802 29588 12808 29640
rect 12860 29628 12866 29640
rect 13081 29631 13139 29637
rect 13081 29628 13093 29631
rect 12860 29600 13093 29628
rect 12860 29588 12866 29600
rect 13081 29597 13093 29600
rect 13127 29597 13139 29631
rect 13081 29591 13139 29597
rect 13722 29588 13728 29640
rect 13780 29628 13786 29640
rect 17034 29628 17040 29640
rect 13780 29600 17040 29628
rect 13780 29588 13786 29600
rect 17034 29588 17040 29600
rect 17092 29588 17098 29640
rect 19981 29631 20039 29637
rect 19981 29597 19993 29631
rect 20027 29628 20039 29631
rect 20714 29628 20720 29640
rect 20027 29600 20720 29628
rect 20027 29597 20039 29600
rect 19981 29591 20039 29597
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 3878 29520 3884 29572
rect 3936 29560 3942 29572
rect 4433 29563 4491 29569
rect 4433 29560 4445 29563
rect 3936 29532 4445 29560
rect 3936 29520 3942 29532
rect 4433 29529 4445 29532
rect 4479 29529 4491 29563
rect 4433 29523 4491 29529
rect 6086 29520 6092 29572
rect 6144 29520 6150 29572
rect 7098 29520 7104 29572
rect 7156 29560 7162 29572
rect 8297 29563 8355 29569
rect 8297 29560 8309 29563
rect 7156 29532 8309 29560
rect 7156 29520 7162 29532
rect 7374 29452 7380 29504
rect 7432 29492 7438 29504
rect 7484 29501 7512 29532
rect 8297 29529 8309 29532
rect 8343 29529 8355 29563
rect 8297 29523 8355 29529
rect 9582 29520 9588 29572
rect 9640 29560 9646 29572
rect 9861 29563 9919 29569
rect 9861 29560 9873 29563
rect 9640 29532 9873 29560
rect 9640 29520 9646 29532
rect 9861 29529 9873 29532
rect 9907 29529 9919 29563
rect 9861 29523 9919 29529
rect 9950 29520 9956 29572
rect 10008 29520 10014 29572
rect 12986 29520 12992 29572
rect 13044 29520 13050 29572
rect 14734 29520 14740 29572
rect 14792 29520 14798 29572
rect 16390 29520 16396 29572
rect 16448 29560 16454 29572
rect 17313 29563 17371 29569
rect 16448 29532 17264 29560
rect 16448 29520 16454 29532
rect 7469 29495 7527 29501
rect 7469 29492 7481 29495
rect 7432 29464 7481 29492
rect 7432 29452 7438 29464
rect 7469 29461 7481 29464
rect 7515 29461 7527 29495
rect 7469 29455 7527 29461
rect 7650 29452 7656 29504
rect 7708 29492 7714 29504
rect 8205 29495 8263 29501
rect 8205 29492 8217 29495
rect 7708 29464 8217 29492
rect 7708 29452 7714 29464
rect 8205 29461 8217 29464
rect 8251 29461 8263 29495
rect 8205 29455 8263 29461
rect 9217 29495 9275 29501
rect 9217 29461 9229 29495
rect 9263 29492 9275 29495
rect 9968 29492 9996 29520
rect 10686 29492 10692 29504
rect 9263 29464 10692 29492
rect 9263 29461 9275 29464
rect 9217 29455 9275 29461
rect 10686 29452 10692 29464
rect 10744 29452 10750 29504
rect 10778 29452 10784 29504
rect 10836 29492 10842 29504
rect 11425 29495 11483 29501
rect 11425 29492 11437 29495
rect 10836 29464 11437 29492
rect 10836 29452 10842 29464
rect 11425 29461 11437 29464
rect 11471 29461 11483 29495
rect 11425 29455 11483 29461
rect 11882 29452 11888 29504
rect 11940 29452 11946 29504
rect 15102 29452 15108 29504
rect 15160 29492 15166 29504
rect 16945 29495 17003 29501
rect 16945 29492 16957 29495
rect 15160 29464 16957 29492
rect 15160 29452 15166 29464
rect 16945 29461 16957 29464
rect 16991 29461 17003 29495
rect 17236 29492 17264 29532
rect 17313 29529 17325 29563
rect 17359 29560 17371 29563
rect 17586 29560 17592 29572
rect 17359 29532 17592 29560
rect 17359 29529 17371 29532
rect 17313 29523 17371 29529
rect 17586 29520 17592 29532
rect 17644 29520 17650 29572
rect 18601 29563 18659 29569
rect 18601 29529 18613 29563
rect 18647 29560 18659 29563
rect 19334 29560 19340 29572
rect 18647 29532 19340 29560
rect 18647 29529 18659 29532
rect 18601 29523 18659 29529
rect 19334 29520 19340 29532
rect 19392 29560 19398 29572
rect 21284 29560 21312 29736
rect 25133 29733 25145 29736
rect 25179 29733 25191 29767
rect 25133 29727 25191 29733
rect 22189 29699 22247 29705
rect 22189 29665 22201 29699
rect 22235 29696 22247 29699
rect 22554 29696 22560 29708
rect 22235 29668 22560 29696
rect 22235 29665 22247 29668
rect 22189 29659 22247 29665
rect 22554 29656 22560 29668
rect 22612 29656 22618 29708
rect 23382 29656 23388 29708
rect 23440 29656 23446 29708
rect 23569 29699 23627 29705
rect 23569 29665 23581 29699
rect 23615 29696 23627 29699
rect 23750 29696 23756 29708
rect 23615 29668 23756 29696
rect 23615 29665 23627 29668
rect 23569 29659 23627 29665
rect 23750 29656 23756 29668
rect 23808 29656 23814 29708
rect 21913 29631 21971 29637
rect 21913 29597 21925 29631
rect 21959 29628 21971 29631
rect 22002 29628 22008 29640
rect 21959 29600 22008 29628
rect 21959 29597 21971 29600
rect 21913 29591 21971 29597
rect 22002 29588 22008 29600
rect 22060 29588 22066 29640
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 19392 29532 21312 29560
rect 19392 29520 19398 29532
rect 21450 29520 21456 29572
rect 21508 29560 21514 29572
rect 21508 29532 21680 29560
rect 21508 29520 21514 29532
rect 17405 29495 17463 29501
rect 17405 29492 17417 29495
rect 17236 29464 17417 29492
rect 16945 29455 17003 29461
rect 17405 29461 17417 29464
rect 17451 29461 17463 29495
rect 17405 29455 17463 29461
rect 17494 29452 17500 29504
rect 17552 29492 17558 29504
rect 18141 29495 18199 29501
rect 18141 29492 18153 29495
rect 17552 29464 18153 29492
rect 17552 29452 17558 29464
rect 18141 29461 18153 29464
rect 18187 29461 18199 29495
rect 18141 29455 18199 29461
rect 18509 29495 18567 29501
rect 18509 29461 18521 29495
rect 18555 29492 18567 29495
rect 19058 29492 19064 29504
rect 18555 29464 19064 29492
rect 18555 29461 18567 29464
rect 18509 29455 18567 29461
rect 19058 29452 19064 29464
rect 19116 29452 19122 29504
rect 19613 29495 19671 29501
rect 19613 29461 19625 29495
rect 19659 29492 19671 29495
rect 20346 29492 20352 29504
rect 19659 29464 20352 29492
rect 19659 29461 19671 29464
rect 19613 29455 19671 29461
rect 20346 29452 20352 29464
rect 20404 29452 20410 29504
rect 20898 29452 20904 29504
rect 20956 29452 20962 29504
rect 21542 29452 21548 29504
rect 21600 29452 21606 29504
rect 21652 29492 21680 29532
rect 21726 29520 21732 29572
rect 21784 29560 21790 29572
rect 23842 29560 23848 29572
rect 21784 29532 23848 29560
rect 21784 29520 21790 29532
rect 23842 29520 23848 29532
rect 23900 29520 23906 29572
rect 22005 29495 22063 29501
rect 22005 29492 22017 29495
rect 21652 29464 22017 29492
rect 22005 29461 22017 29464
rect 22051 29461 22063 29495
rect 22005 29455 22063 29461
rect 22830 29452 22836 29504
rect 22888 29492 22894 29504
rect 22925 29495 22983 29501
rect 22925 29492 22937 29495
rect 22888 29464 22937 29492
rect 22888 29452 22894 29464
rect 22925 29461 22937 29464
rect 22971 29461 22983 29495
rect 22925 29455 22983 29461
rect 23290 29452 23296 29504
rect 23348 29452 23354 29504
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 7650 29248 7656 29300
rect 7708 29288 7714 29300
rect 7708 29260 9352 29288
rect 7708 29248 7714 29260
rect 9030 29180 9036 29232
rect 9088 29180 9094 29232
rect 9324 29220 9352 29260
rect 9766 29248 9772 29300
rect 9824 29248 9830 29300
rect 11238 29248 11244 29300
rect 11296 29288 11302 29300
rect 14921 29291 14979 29297
rect 14921 29288 14933 29291
rect 11296 29260 14933 29288
rect 11296 29248 11302 29260
rect 14921 29257 14933 29260
rect 14967 29257 14979 29291
rect 14921 29251 14979 29257
rect 15289 29291 15347 29297
rect 15289 29257 15301 29291
rect 15335 29288 15347 29291
rect 15654 29288 15660 29300
rect 15335 29260 15660 29288
rect 15335 29257 15347 29260
rect 15289 29251 15347 29257
rect 15654 29248 15660 29260
rect 15712 29288 15718 29300
rect 15933 29291 15991 29297
rect 15933 29288 15945 29291
rect 15712 29260 15945 29288
rect 15712 29248 15718 29260
rect 15933 29257 15945 29260
rect 15979 29257 15991 29291
rect 15933 29251 15991 29257
rect 17218 29248 17224 29300
rect 17276 29248 17282 29300
rect 17313 29291 17371 29297
rect 17313 29257 17325 29291
rect 17359 29288 17371 29291
rect 17494 29288 17500 29300
rect 17359 29260 17500 29288
rect 17359 29257 17371 29260
rect 17313 29251 17371 29257
rect 17494 29248 17500 29260
rect 17552 29248 17558 29300
rect 17586 29248 17592 29300
rect 17644 29288 17650 29300
rect 17957 29291 18015 29297
rect 17957 29288 17969 29291
rect 17644 29260 17969 29288
rect 17644 29248 17650 29260
rect 17957 29257 17969 29260
rect 18003 29288 18015 29291
rect 19518 29288 19524 29300
rect 18003 29260 19524 29288
rect 18003 29257 18015 29260
rect 17957 29251 18015 29257
rect 19518 29248 19524 29260
rect 19576 29248 19582 29300
rect 20073 29291 20131 29297
rect 20073 29257 20085 29291
rect 20119 29257 20131 29291
rect 20073 29251 20131 29257
rect 20533 29291 20591 29297
rect 20533 29257 20545 29291
rect 20579 29288 20591 29291
rect 20806 29288 20812 29300
rect 20579 29260 20812 29288
rect 20579 29257 20591 29260
rect 20533 29251 20591 29257
rect 9324 29192 14320 29220
rect 12897 29155 12955 29161
rect 9508 29124 12480 29152
rect 6546 29044 6552 29096
rect 6604 29084 6610 29096
rect 7745 29087 7803 29093
rect 7745 29084 7757 29087
rect 6604 29056 7757 29084
rect 6604 29044 6610 29056
rect 7745 29053 7757 29056
rect 7791 29053 7803 29087
rect 7745 29047 7803 29053
rect 9398 29044 9404 29096
rect 9456 29084 9462 29096
rect 9508 29093 9536 29124
rect 9493 29087 9551 29093
rect 9493 29084 9505 29087
rect 9456 29056 9505 29084
rect 9456 29044 9462 29056
rect 9493 29053 9505 29056
rect 9539 29053 9551 29087
rect 9766 29084 9772 29096
rect 9493 29047 9551 29053
rect 9600 29056 9772 29084
rect 9030 28976 9036 29028
rect 9088 29016 9094 29028
rect 9600 29016 9628 29056
rect 9766 29044 9772 29056
rect 9824 29044 9830 29096
rect 12452 29084 12480 29124
rect 12897 29121 12909 29155
rect 12943 29152 12955 29155
rect 13722 29152 13728 29164
rect 12943 29124 13728 29152
rect 12943 29121 12955 29124
rect 12897 29115 12955 29121
rect 13722 29112 13728 29124
rect 13780 29112 13786 29164
rect 14090 29112 14096 29164
rect 14148 29112 14154 29164
rect 14182 29112 14188 29164
rect 14240 29112 14246 29164
rect 14292 29152 14320 29192
rect 15562 29180 15568 29232
rect 15620 29220 15626 29232
rect 16209 29223 16267 29229
rect 16209 29220 16221 29223
rect 15620 29192 16221 29220
rect 15620 29180 15626 29192
rect 16209 29189 16221 29192
rect 16255 29220 16267 29223
rect 16298 29220 16304 29232
rect 16255 29192 16304 29220
rect 16255 29189 16267 29192
rect 16209 29183 16267 29189
rect 16298 29180 16304 29192
rect 16356 29220 16362 29232
rect 18322 29220 18328 29232
rect 16356 29192 18328 29220
rect 16356 29180 16362 29192
rect 18322 29180 18328 29192
rect 18380 29180 18386 29232
rect 20088 29220 20116 29251
rect 20806 29248 20812 29260
rect 20864 29248 20870 29300
rect 20898 29248 20904 29300
rect 20956 29288 20962 29300
rect 22373 29291 22431 29297
rect 22373 29288 22385 29291
rect 20956 29260 22385 29288
rect 20956 29248 20962 29260
rect 22373 29257 22385 29260
rect 22419 29257 22431 29291
rect 22373 29251 22431 29257
rect 23842 29248 23848 29300
rect 23900 29288 23906 29300
rect 23937 29291 23995 29297
rect 23937 29288 23949 29291
rect 23900 29260 23949 29288
rect 23900 29248 23906 29260
rect 23937 29257 23949 29260
rect 23983 29257 23995 29291
rect 23937 29251 23995 29257
rect 25314 29248 25320 29300
rect 25372 29248 25378 29300
rect 25498 29248 25504 29300
rect 25556 29248 25562 29300
rect 22462 29220 22468 29232
rect 20088 29192 22468 29220
rect 22462 29180 22468 29192
rect 22520 29180 22526 29232
rect 24578 29180 24584 29232
rect 24636 29220 24642 29232
rect 24673 29223 24731 29229
rect 24673 29220 24685 29223
rect 24636 29192 24685 29220
rect 24636 29180 24642 29192
rect 24673 29189 24685 29192
rect 24719 29189 24731 29223
rect 24673 29183 24731 29189
rect 14292 29124 15516 29152
rect 12989 29087 13047 29093
rect 12452 29056 12756 29084
rect 9088 28988 9628 29016
rect 9088 28976 9094 28988
rect 10870 28976 10876 29028
rect 10928 29016 10934 29028
rect 12529 29019 12587 29025
rect 12529 29016 12541 29019
rect 10928 28988 12541 29016
rect 10928 28976 10934 28988
rect 12529 28985 12541 28988
rect 12575 28985 12587 29019
rect 12728 29016 12756 29056
rect 12989 29053 13001 29087
rect 13035 29084 13047 29087
rect 13078 29084 13084 29096
rect 13035 29056 13084 29084
rect 13035 29053 13047 29056
rect 12989 29047 13047 29053
rect 13078 29044 13084 29056
rect 13136 29044 13142 29096
rect 13173 29087 13231 29093
rect 13173 29053 13185 29087
rect 13219 29053 13231 29087
rect 13173 29047 13231 29053
rect 13188 29016 13216 29047
rect 13262 29044 13268 29096
rect 13320 29084 13326 29096
rect 13906 29084 13912 29096
rect 13320 29056 13912 29084
rect 13320 29044 13326 29056
rect 13906 29044 13912 29056
rect 13964 29084 13970 29096
rect 14274 29084 14280 29096
rect 13964 29056 14280 29084
rect 13964 29044 13970 29056
rect 14274 29044 14280 29056
rect 14332 29044 14338 29096
rect 14369 29087 14427 29093
rect 14369 29053 14381 29087
rect 14415 29084 14427 29087
rect 14642 29084 14648 29096
rect 14415 29056 14648 29084
rect 14415 29053 14427 29056
rect 14369 29047 14427 29053
rect 14642 29044 14648 29056
rect 14700 29044 14706 29096
rect 15194 29044 15200 29096
rect 15252 29084 15258 29096
rect 15488 29093 15516 29124
rect 16390 29112 16396 29164
rect 16448 29152 16454 29164
rect 16485 29155 16543 29161
rect 16485 29152 16497 29155
rect 16448 29124 16497 29152
rect 16448 29112 16454 29124
rect 16485 29121 16497 29124
rect 16531 29152 16543 29155
rect 19705 29155 19763 29161
rect 19705 29152 19717 29155
rect 16531 29124 19717 29152
rect 16531 29121 16543 29124
rect 16485 29115 16543 29121
rect 19705 29121 19717 29124
rect 19751 29152 19763 29155
rect 20441 29155 20499 29161
rect 20441 29152 20453 29155
rect 19751 29124 20453 29152
rect 19751 29121 19763 29124
rect 19705 29115 19763 29121
rect 20441 29121 20453 29124
rect 20487 29121 20499 29155
rect 20441 29115 20499 29121
rect 21450 29112 21456 29164
rect 21508 29152 21514 29164
rect 21545 29155 21603 29161
rect 21545 29152 21557 29155
rect 21508 29124 21557 29152
rect 21508 29112 21514 29124
rect 21545 29121 21557 29124
rect 21591 29121 21603 29155
rect 21545 29115 21603 29121
rect 23661 29155 23719 29161
rect 23661 29121 23673 29155
rect 23707 29152 23719 29155
rect 24118 29152 24124 29164
rect 23707 29124 24124 29152
rect 23707 29121 23719 29124
rect 23661 29115 23719 29121
rect 15381 29087 15439 29093
rect 15381 29084 15393 29087
rect 15252 29056 15393 29084
rect 15252 29044 15258 29056
rect 15381 29053 15393 29056
rect 15427 29053 15439 29087
rect 15381 29047 15439 29053
rect 15473 29087 15531 29093
rect 15473 29053 15485 29087
rect 15519 29053 15531 29087
rect 15473 29047 15531 29053
rect 17402 29044 17408 29096
rect 17460 29044 17466 29096
rect 17586 29044 17592 29096
rect 17644 29084 17650 29096
rect 17770 29084 17776 29096
rect 17644 29056 17776 29084
rect 17644 29044 17650 29056
rect 17770 29044 17776 29056
rect 17828 29044 17834 29096
rect 17880 29056 19656 29084
rect 12728 28988 13216 29016
rect 12529 28979 12587 28985
rect 13446 28976 13452 29028
rect 13504 29016 13510 29028
rect 13725 29019 13783 29025
rect 13725 29016 13737 29019
rect 13504 28988 13737 29016
rect 13504 28976 13510 28988
rect 13725 28985 13737 28988
rect 13771 28985 13783 29019
rect 13725 28979 13783 28985
rect 16022 28976 16028 29028
rect 16080 29016 16086 29028
rect 16853 29019 16911 29025
rect 16853 29016 16865 29019
rect 16080 28988 16865 29016
rect 16080 28976 16086 28988
rect 16853 28985 16865 28988
rect 16899 28985 16911 29019
rect 16853 28979 16911 28985
rect 16942 28976 16948 29028
rect 17000 29016 17006 29028
rect 17880 29016 17908 29056
rect 19628 29028 19656 29056
rect 20162 29044 20168 29096
rect 20220 29084 20226 29096
rect 20625 29087 20683 29093
rect 20625 29084 20637 29087
rect 20220 29056 20637 29084
rect 20220 29044 20226 29056
rect 20625 29053 20637 29056
rect 20671 29053 20683 29087
rect 21560 29084 21588 29115
rect 24118 29112 24124 29124
rect 24176 29112 24182 29164
rect 22465 29087 22523 29093
rect 22465 29084 22477 29087
rect 21560 29056 22477 29084
rect 20625 29047 20683 29053
rect 22465 29053 22477 29056
rect 22511 29053 22523 29087
rect 22465 29047 22523 29053
rect 22649 29087 22707 29093
rect 22649 29053 22661 29087
rect 22695 29084 22707 29087
rect 23566 29084 23572 29096
rect 22695 29056 23572 29084
rect 22695 29053 22707 29056
rect 22649 29047 22707 29053
rect 23566 29044 23572 29056
rect 23624 29044 23630 29096
rect 17000 28988 17908 29016
rect 18049 29019 18107 29025
rect 17000 28976 17006 28988
rect 18049 28985 18061 29019
rect 18095 29016 18107 29019
rect 19058 29016 19064 29028
rect 18095 28988 19064 29016
rect 18095 28985 18107 28988
rect 18049 28979 18107 28985
rect 8008 28951 8066 28957
rect 8008 28917 8020 28951
rect 8054 28948 8066 28951
rect 8662 28948 8668 28960
rect 8054 28920 8668 28948
rect 8054 28917 8066 28920
rect 8008 28911 8066 28917
rect 8662 28908 8668 28920
rect 8720 28908 8726 28960
rect 16114 28908 16120 28960
rect 16172 28948 16178 28960
rect 18064 28948 18092 28979
rect 19058 28976 19064 28988
rect 19116 28976 19122 29028
rect 19610 28976 19616 29028
rect 19668 29016 19674 29028
rect 20806 29016 20812 29028
rect 19668 28988 20812 29016
rect 19668 28976 19674 28988
rect 20806 28976 20812 28988
rect 20864 28976 20870 29028
rect 20898 28976 20904 29028
rect 20956 29016 20962 29028
rect 21085 29019 21143 29025
rect 21085 29016 21097 29019
rect 20956 28988 21097 29016
rect 20956 28976 20962 28988
rect 21085 28985 21097 28988
rect 21131 28985 21143 29019
rect 21085 28979 21143 28985
rect 22005 29019 22063 29025
rect 22005 28985 22017 29019
rect 22051 29016 22063 29019
rect 23290 29016 23296 29028
rect 22051 28988 23296 29016
rect 22051 28985 22063 28988
rect 22005 28979 22063 28985
rect 23290 28976 23296 28988
rect 23348 28976 23354 29028
rect 23474 28976 23480 29028
rect 23532 29016 23538 29028
rect 24857 29019 24915 29025
rect 24857 29016 24869 29019
rect 23532 28988 24869 29016
rect 23532 28976 23538 28988
rect 24857 28985 24869 28988
rect 24903 28985 24915 29019
rect 24857 28979 24915 28985
rect 16172 28920 18092 28948
rect 16172 28908 16178 28920
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 12805 28747 12863 28753
rect 12805 28713 12817 28747
rect 12851 28744 12863 28747
rect 14090 28744 14096 28756
rect 12851 28716 14096 28744
rect 12851 28713 12863 28716
rect 12805 28707 12863 28713
rect 14090 28704 14096 28716
rect 14148 28704 14154 28756
rect 14734 28704 14740 28756
rect 14792 28744 14798 28756
rect 16761 28747 16819 28753
rect 16761 28744 16773 28747
rect 14792 28716 16773 28744
rect 14792 28704 14798 28716
rect 16761 28713 16773 28716
rect 16807 28744 16819 28747
rect 21266 28744 21272 28756
rect 16807 28716 21272 28744
rect 16807 28713 16819 28716
rect 16761 28707 16819 28713
rect 21266 28704 21272 28716
rect 21324 28704 21330 28756
rect 21450 28704 21456 28756
rect 21508 28744 21514 28756
rect 24302 28744 24308 28756
rect 21508 28716 24308 28744
rect 21508 28704 21514 28716
rect 24302 28704 24308 28716
rect 24360 28704 24366 28756
rect 21174 28636 21180 28688
rect 21232 28636 21238 28688
rect 1302 28568 1308 28620
rect 1360 28608 1366 28620
rect 2041 28611 2099 28617
rect 2041 28608 2053 28611
rect 1360 28580 2053 28608
rect 1360 28568 1366 28580
rect 2041 28577 2053 28580
rect 2087 28577 2099 28611
rect 2041 28571 2099 28577
rect 3418 28568 3424 28620
rect 3476 28608 3482 28620
rect 4249 28611 4307 28617
rect 4249 28608 4261 28611
rect 3476 28580 4261 28608
rect 3476 28568 3482 28580
rect 4249 28577 4261 28580
rect 4295 28577 4307 28611
rect 4249 28571 4307 28577
rect 5902 28568 5908 28620
rect 5960 28568 5966 28620
rect 6546 28568 6552 28620
rect 6604 28568 6610 28620
rect 6825 28611 6883 28617
rect 6825 28577 6837 28611
rect 6871 28608 6883 28611
rect 8297 28611 8355 28617
rect 6871 28580 8248 28608
rect 6871 28577 6883 28580
rect 6825 28571 6883 28577
rect 1762 28500 1768 28552
rect 1820 28500 1826 28552
rect 8220 28540 8248 28580
rect 8297 28577 8309 28611
rect 8343 28608 8355 28611
rect 9858 28608 9864 28620
rect 8343 28580 9864 28608
rect 8343 28577 8355 28580
rect 8297 28571 8355 28577
rect 9858 28568 9864 28580
rect 9916 28568 9922 28620
rect 10873 28611 10931 28617
rect 10873 28577 10885 28611
rect 10919 28608 10931 28611
rect 11330 28608 11336 28620
rect 10919 28580 11336 28608
rect 10919 28577 10931 28580
rect 10873 28571 10931 28577
rect 11330 28568 11336 28580
rect 11388 28568 11394 28620
rect 13354 28568 13360 28620
rect 13412 28568 13418 28620
rect 13630 28568 13636 28620
rect 13688 28608 13694 28620
rect 14829 28611 14887 28617
rect 14829 28608 14841 28611
rect 13688 28580 14841 28608
rect 13688 28568 13694 28580
rect 14829 28577 14841 28580
rect 14875 28577 14887 28611
rect 14829 28571 14887 28577
rect 16206 28568 16212 28620
rect 16264 28568 16270 28620
rect 17126 28568 17132 28620
rect 17184 28608 17190 28620
rect 17681 28611 17739 28617
rect 17681 28608 17693 28611
rect 17184 28580 17693 28608
rect 17184 28568 17190 28580
rect 17681 28577 17693 28580
rect 17727 28577 17739 28611
rect 17681 28571 17739 28577
rect 17770 28568 17776 28620
rect 17828 28568 17834 28620
rect 19429 28611 19487 28617
rect 19429 28577 19441 28611
rect 19475 28608 19487 28611
rect 22002 28608 22008 28620
rect 19475 28580 22008 28608
rect 19475 28577 19487 28580
rect 19429 28571 19487 28577
rect 22002 28568 22008 28580
rect 22060 28568 22066 28620
rect 22830 28568 22836 28620
rect 22888 28608 22894 28620
rect 22888 28580 24808 28608
rect 22888 28568 22894 28580
rect 9398 28540 9404 28552
rect 8220 28512 9404 28540
rect 9398 28500 9404 28512
rect 9456 28500 9462 28552
rect 9950 28500 9956 28552
rect 10008 28540 10014 28552
rect 10597 28543 10655 28549
rect 10597 28540 10609 28543
rect 10008 28512 10609 28540
rect 10008 28500 10014 28512
rect 10597 28509 10609 28512
rect 10643 28509 10655 28543
rect 10597 28503 10655 28509
rect 14645 28543 14703 28549
rect 14645 28509 14657 28543
rect 14691 28540 14703 28543
rect 15562 28540 15568 28552
rect 14691 28512 15568 28540
rect 14691 28509 14703 28512
rect 14645 28503 14703 28509
rect 15562 28500 15568 28512
rect 15620 28500 15626 28552
rect 16022 28500 16028 28552
rect 16080 28500 16086 28552
rect 16117 28543 16175 28549
rect 16117 28509 16129 28543
rect 16163 28540 16175 28543
rect 16850 28540 16856 28552
rect 16163 28512 16856 28540
rect 16163 28509 16175 28512
rect 16117 28503 16175 28509
rect 16850 28500 16856 28512
rect 16908 28500 16914 28552
rect 17589 28543 17647 28549
rect 17589 28509 17601 28543
rect 17635 28540 17647 28543
rect 18598 28540 18604 28552
rect 17635 28512 18604 28540
rect 17635 28509 17647 28512
rect 17589 28503 17647 28509
rect 18598 28500 18604 28512
rect 18656 28500 18662 28552
rect 24780 28549 24808 28580
rect 24029 28543 24087 28549
rect 24029 28509 24041 28543
rect 24075 28509 24087 28543
rect 24029 28503 24087 28509
rect 24765 28543 24823 28549
rect 24765 28509 24777 28543
rect 24811 28509 24823 28543
rect 24765 28503 24823 28509
rect 3970 28432 3976 28484
rect 4028 28472 4034 28484
rect 4433 28475 4491 28481
rect 4433 28472 4445 28475
rect 4028 28444 4445 28472
rect 4028 28432 4034 28444
rect 4433 28441 4445 28444
rect 4479 28441 4491 28475
rect 12526 28472 12532 28484
rect 8050 28444 8708 28472
rect 12098 28444 12532 28472
rect 4433 28435 4491 28441
rect 8680 28413 8708 28444
rect 12526 28432 12532 28444
rect 12584 28432 12590 28484
rect 13078 28432 13084 28484
rect 13136 28472 13142 28484
rect 13265 28475 13323 28481
rect 13265 28472 13277 28475
rect 13136 28444 13277 28472
rect 13136 28432 13142 28444
rect 13265 28441 13277 28444
rect 13311 28441 13323 28475
rect 13265 28435 13323 28441
rect 19705 28475 19763 28481
rect 19705 28441 19717 28475
rect 19751 28472 19763 28475
rect 19794 28472 19800 28484
rect 19751 28444 19800 28472
rect 19751 28441 19763 28444
rect 19705 28435 19763 28441
rect 19794 28432 19800 28444
rect 19852 28432 19858 28484
rect 21450 28472 21456 28484
rect 20930 28444 21456 28472
rect 21450 28432 21456 28444
rect 21508 28432 21514 28484
rect 24044 28472 24072 28503
rect 24210 28472 24216 28484
rect 24044 28444 24216 28472
rect 24210 28432 24216 28444
rect 24268 28472 24274 28484
rect 24854 28472 24860 28484
rect 24268 28444 24860 28472
rect 24268 28432 24274 28444
rect 24854 28432 24860 28444
rect 24912 28432 24918 28484
rect 8665 28407 8723 28413
rect 8665 28373 8677 28407
rect 8711 28404 8723 28407
rect 9030 28404 9036 28416
rect 8711 28376 9036 28404
rect 8711 28373 8723 28376
rect 8665 28367 8723 28373
rect 9030 28364 9036 28376
rect 9088 28404 9094 28416
rect 9582 28404 9588 28416
rect 9088 28376 9588 28404
rect 9088 28364 9094 28376
rect 9582 28364 9588 28376
rect 9640 28364 9646 28416
rect 12345 28407 12403 28413
rect 12345 28373 12357 28407
rect 12391 28404 12403 28407
rect 12802 28404 12808 28416
rect 12391 28376 12808 28404
rect 12391 28373 12403 28376
rect 12345 28367 12403 28373
rect 12802 28364 12808 28376
rect 12860 28364 12866 28416
rect 13170 28364 13176 28416
rect 13228 28364 13234 28416
rect 13909 28407 13967 28413
rect 13909 28373 13921 28407
rect 13955 28404 13967 28407
rect 13998 28404 14004 28416
rect 13955 28376 14004 28404
rect 13955 28373 13967 28376
rect 13909 28367 13967 28373
rect 13998 28364 14004 28376
rect 14056 28364 14062 28416
rect 14274 28364 14280 28416
rect 14332 28364 14338 28416
rect 14734 28364 14740 28416
rect 14792 28364 14798 28416
rect 15194 28364 15200 28416
rect 15252 28404 15258 28416
rect 15289 28407 15347 28413
rect 15289 28404 15301 28407
rect 15252 28376 15301 28404
rect 15252 28364 15258 28376
rect 15289 28373 15301 28376
rect 15335 28373 15347 28407
rect 15289 28367 15347 28373
rect 15657 28407 15715 28413
rect 15657 28373 15669 28407
rect 15703 28404 15715 28407
rect 15746 28404 15752 28416
rect 15703 28376 15752 28404
rect 15703 28373 15715 28376
rect 15657 28367 15715 28373
rect 15746 28364 15752 28376
rect 15804 28364 15810 28416
rect 16942 28364 16948 28416
rect 17000 28404 17006 28416
rect 17221 28407 17279 28413
rect 17221 28404 17233 28407
rect 17000 28376 17233 28404
rect 17000 28364 17006 28376
rect 17221 28373 17233 28376
rect 17267 28373 17279 28407
rect 17221 28367 17279 28373
rect 18414 28364 18420 28416
rect 18472 28404 18478 28416
rect 23845 28407 23903 28413
rect 23845 28404 23857 28407
rect 18472 28376 23857 28404
rect 18472 28364 18478 28376
rect 23845 28373 23857 28376
rect 23891 28373 23903 28407
rect 23845 28367 23903 28373
rect 24578 28364 24584 28416
rect 24636 28364 24642 28416
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 1946 28160 1952 28212
rect 2004 28200 2010 28212
rect 3786 28209 3792 28212
rect 2041 28203 2099 28209
rect 2041 28200 2053 28203
rect 2004 28172 2053 28200
rect 2004 28160 2010 28172
rect 2041 28169 2053 28172
rect 2087 28169 2099 28203
rect 2041 28163 2099 28169
rect 3743 28203 3792 28209
rect 3743 28169 3755 28203
rect 3789 28169 3792 28203
rect 3743 28163 3792 28169
rect 3786 28160 3792 28163
rect 3844 28160 3850 28212
rect 5902 28160 5908 28212
rect 5960 28200 5966 28212
rect 12621 28203 12679 28209
rect 5960 28172 12434 28200
rect 5960 28160 5966 28172
rect 9030 28092 9036 28144
rect 9088 28092 9094 28144
rect 12406 28132 12434 28172
rect 12621 28169 12633 28203
rect 12667 28200 12679 28203
rect 13170 28200 13176 28212
rect 12667 28172 13176 28200
rect 12667 28169 12679 28172
rect 12621 28163 12679 28169
rect 13170 28160 13176 28172
rect 13228 28160 13234 28212
rect 15654 28160 15660 28212
rect 15712 28200 15718 28212
rect 15930 28200 15936 28212
rect 15712 28172 15936 28200
rect 15712 28160 15718 28172
rect 15930 28160 15936 28172
rect 15988 28200 15994 28212
rect 16669 28203 16727 28209
rect 16669 28200 16681 28203
rect 15988 28172 16681 28200
rect 15988 28160 15994 28172
rect 16669 28169 16681 28172
rect 16715 28169 16727 28203
rect 16669 28163 16727 28169
rect 18322 28160 18328 28212
rect 18380 28160 18386 28212
rect 19521 28203 19579 28209
rect 19521 28169 19533 28203
rect 19567 28200 19579 28203
rect 20165 28203 20223 28209
rect 20165 28200 20177 28203
rect 19567 28172 20177 28200
rect 19567 28169 19579 28172
rect 19521 28163 19579 28169
rect 20165 28169 20177 28172
rect 20211 28200 20223 28203
rect 20254 28200 20260 28212
rect 20211 28172 20260 28200
rect 20211 28169 20223 28172
rect 20165 28163 20223 28169
rect 20254 28160 20260 28172
rect 20312 28160 20318 28212
rect 23753 28203 23811 28209
rect 23753 28200 23765 28203
rect 22066 28172 23765 28200
rect 16114 28132 16120 28144
rect 12406 28104 16120 28132
rect 16114 28092 16120 28104
rect 16172 28092 16178 28144
rect 18506 28132 18512 28144
rect 16224 28104 18512 28132
rect 2225 28067 2283 28073
rect 2225 28033 2237 28067
rect 2271 28064 2283 28067
rect 3418 28064 3424 28076
rect 2271 28036 3424 28064
rect 2271 28033 2283 28036
rect 2225 28027 2283 28033
rect 3418 28024 3424 28036
rect 3476 28024 3482 28076
rect 3602 28024 3608 28076
rect 3660 28073 3666 28076
rect 3660 28067 3698 28073
rect 3686 28033 3698 28067
rect 3660 28027 3698 28033
rect 3660 28024 3666 28027
rect 9582 28024 9588 28076
rect 9640 28064 9646 28076
rect 10321 28067 10379 28073
rect 10321 28064 10333 28067
rect 9640 28036 10333 28064
rect 9640 28024 9646 28036
rect 10321 28033 10333 28036
rect 10367 28064 10379 28067
rect 12526 28064 12532 28076
rect 10367 28036 12532 28064
rect 10367 28033 10379 28036
rect 10321 28027 10379 28033
rect 12526 28024 12532 28036
rect 12584 28064 12590 28076
rect 13354 28064 13360 28076
rect 12584 28036 13360 28064
rect 12584 28024 12590 28036
rect 13354 28024 13360 28036
rect 13412 28024 13418 28076
rect 15194 28024 15200 28076
rect 15252 28064 15258 28076
rect 15838 28064 15844 28076
rect 15252 28036 15844 28064
rect 15252 28024 15258 28036
rect 15838 28024 15844 28036
rect 15896 28024 15902 28076
rect 15930 28024 15936 28076
rect 15988 28064 15994 28076
rect 16224 28064 16252 28104
rect 18506 28092 18512 28104
rect 18564 28092 18570 28144
rect 18782 28092 18788 28144
rect 18840 28132 18846 28144
rect 22066 28132 22094 28172
rect 23753 28169 23765 28172
rect 23799 28169 23811 28203
rect 23753 28163 23811 28169
rect 24213 28203 24271 28209
rect 24213 28169 24225 28203
rect 24259 28200 24271 28203
rect 24302 28200 24308 28212
rect 24259 28172 24308 28200
rect 24259 28169 24271 28172
rect 24213 28163 24271 28169
rect 24228 28132 24256 28163
rect 24302 28160 24308 28172
rect 24360 28160 24366 28212
rect 18840 28104 22094 28132
rect 23506 28104 24256 28132
rect 18840 28092 18846 28104
rect 24670 28092 24676 28144
rect 24728 28092 24734 28144
rect 18233 28067 18291 28073
rect 18233 28064 18245 28067
rect 15988 28036 16252 28064
rect 15988 28024 15994 28036
rect 8297 27999 8355 28005
rect 8297 27965 8309 27999
rect 8343 27965 8355 27999
rect 8297 27959 8355 27965
rect 8312 27860 8340 27959
rect 8570 27956 8576 28008
rect 8628 27956 8634 28008
rect 8662 27956 8668 28008
rect 8720 27996 8726 28008
rect 8720 27968 10088 27996
rect 8720 27956 8726 27968
rect 10060 27937 10088 27968
rect 16022 27956 16028 28008
rect 16080 27956 16086 28008
rect 16224 28005 16252 28036
rect 17512 28036 18245 28064
rect 16209 27999 16267 28005
rect 16209 27965 16221 27999
rect 16255 27965 16267 27999
rect 16209 27959 16267 27965
rect 10045 27931 10103 27937
rect 10045 27897 10057 27931
rect 10091 27928 10103 27931
rect 11790 27928 11796 27940
rect 10091 27900 11796 27928
rect 10091 27897 10103 27900
rect 10045 27891 10103 27897
rect 11790 27888 11796 27900
rect 11848 27888 11854 27940
rect 15286 27928 15292 27940
rect 15120 27900 15292 27928
rect 9950 27860 9956 27872
rect 8312 27832 9956 27860
rect 9950 27820 9956 27832
rect 10008 27820 10014 27872
rect 12618 27820 12624 27872
rect 12676 27860 12682 27872
rect 13078 27860 13084 27872
rect 12676 27832 13084 27860
rect 12676 27820 12682 27832
rect 13078 27820 13084 27832
rect 13136 27820 13142 27872
rect 13354 27820 13360 27872
rect 13412 27820 13418 27872
rect 14734 27820 14740 27872
rect 14792 27860 14798 27872
rect 15120 27869 15148 27900
rect 15286 27888 15292 27900
rect 15344 27928 15350 27940
rect 17512 27937 17540 28036
rect 18233 28033 18245 28036
rect 18279 28033 18291 28067
rect 18233 28027 18291 28033
rect 19429 28067 19487 28073
rect 19429 28033 19441 28067
rect 19475 28064 19487 28067
rect 19518 28064 19524 28076
rect 19475 28036 19524 28064
rect 19475 28033 19487 28036
rect 19429 28027 19487 28033
rect 19518 28024 19524 28036
rect 19576 28024 19582 28076
rect 22002 28024 22008 28076
rect 22060 28024 22066 28076
rect 18506 27956 18512 28008
rect 18564 27996 18570 28008
rect 18966 27996 18972 28008
rect 18564 27968 18972 27996
rect 18564 27956 18570 27968
rect 18966 27956 18972 27968
rect 19024 27956 19030 28008
rect 19058 27956 19064 28008
rect 19116 27996 19122 28008
rect 19610 27996 19616 28008
rect 19116 27968 19616 27996
rect 19116 27956 19122 27968
rect 19610 27956 19616 27968
rect 19668 27956 19674 28008
rect 19705 27999 19763 28005
rect 19705 27965 19717 27999
rect 19751 27996 19763 27999
rect 19978 27996 19984 28008
rect 19751 27968 19984 27996
rect 19751 27965 19763 27968
rect 19705 27959 19763 27965
rect 19978 27956 19984 27968
rect 20036 27956 20042 28008
rect 22281 27999 22339 28005
rect 22281 27965 22293 27999
rect 22327 27996 22339 27999
rect 24670 27996 24676 28008
rect 22327 27968 24676 27996
rect 22327 27965 22339 27968
rect 22281 27959 22339 27965
rect 24670 27956 24676 27968
rect 24728 27956 24734 28008
rect 17497 27931 17555 27937
rect 17497 27928 17509 27931
rect 15344 27900 17509 27928
rect 15344 27888 15350 27900
rect 17497 27897 17509 27900
rect 17543 27897 17555 27931
rect 21358 27928 21364 27940
rect 17497 27891 17555 27897
rect 17696 27900 21364 27928
rect 15105 27863 15163 27869
rect 15105 27860 15117 27863
rect 14792 27832 15117 27860
rect 14792 27820 14798 27832
rect 15105 27829 15117 27832
rect 15151 27829 15163 27863
rect 15105 27823 15163 27829
rect 15562 27820 15568 27872
rect 15620 27820 15626 27872
rect 16022 27820 16028 27872
rect 16080 27860 16086 27872
rect 16390 27860 16396 27872
rect 16080 27832 16396 27860
rect 16080 27820 16086 27832
rect 16390 27820 16396 27832
rect 16448 27860 16454 27872
rect 16945 27863 17003 27869
rect 16945 27860 16957 27863
rect 16448 27832 16957 27860
rect 16448 27820 16454 27832
rect 16945 27829 16957 27832
rect 16991 27860 17003 27863
rect 17696 27860 17724 27900
rect 21358 27888 21364 27900
rect 21416 27888 21422 27940
rect 24857 27931 24915 27937
rect 24857 27928 24869 27931
rect 23308 27900 24869 27928
rect 16991 27832 17724 27860
rect 17865 27863 17923 27869
rect 16991 27829 17003 27832
rect 16945 27823 17003 27829
rect 17865 27829 17877 27863
rect 17911 27860 17923 27863
rect 18966 27860 18972 27872
rect 17911 27832 18972 27860
rect 17911 27829 17923 27832
rect 17865 27823 17923 27829
rect 18966 27820 18972 27832
rect 19024 27820 19030 27872
rect 19058 27820 19064 27872
rect 19116 27820 19122 27872
rect 22094 27820 22100 27872
rect 22152 27860 22158 27872
rect 23308 27860 23336 27900
rect 24857 27897 24869 27900
rect 24903 27897 24915 27931
rect 24857 27891 24915 27897
rect 22152 27832 23336 27860
rect 22152 27820 22158 27832
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 6444 27659 6502 27665
rect 6444 27625 6456 27659
rect 6490 27656 6502 27659
rect 9858 27656 9864 27668
rect 6490 27628 9864 27656
rect 6490 27625 6502 27628
rect 6444 27619 6502 27625
rect 9858 27616 9864 27628
rect 9916 27616 9922 27668
rect 18322 27616 18328 27668
rect 18380 27656 18386 27668
rect 18693 27659 18751 27665
rect 18693 27656 18705 27659
rect 18380 27628 18705 27656
rect 18380 27616 18386 27628
rect 18693 27625 18705 27628
rect 18739 27656 18751 27659
rect 18782 27656 18788 27668
rect 18739 27628 18788 27656
rect 18739 27625 18751 27628
rect 18693 27619 18751 27625
rect 18782 27616 18788 27628
rect 18840 27616 18846 27668
rect 20990 27656 20996 27668
rect 19996 27628 20996 27656
rect 7834 27548 7840 27600
rect 7892 27588 7898 27600
rect 7929 27591 7987 27597
rect 7929 27588 7941 27591
rect 7892 27560 7941 27588
rect 7892 27548 7898 27560
rect 7929 27557 7941 27560
rect 7975 27557 7987 27591
rect 7929 27551 7987 27557
rect 14182 27548 14188 27600
rect 14240 27588 14246 27600
rect 15378 27588 15384 27600
rect 14240 27560 15384 27588
rect 14240 27548 14246 27560
rect 15378 27548 15384 27560
rect 15436 27548 15442 27600
rect 15838 27548 15844 27600
rect 15896 27588 15902 27600
rect 16206 27588 16212 27600
rect 15896 27560 16212 27588
rect 15896 27548 15902 27560
rect 16206 27548 16212 27560
rect 16264 27588 16270 27600
rect 16393 27591 16451 27597
rect 16393 27588 16405 27591
rect 16264 27560 16405 27588
rect 16264 27548 16270 27560
rect 16393 27557 16405 27560
rect 16439 27588 16451 27591
rect 19996 27588 20024 27628
rect 20990 27616 20996 27628
rect 21048 27616 21054 27668
rect 24210 27616 24216 27668
rect 24268 27616 24274 27668
rect 16439 27560 20024 27588
rect 20073 27591 20131 27597
rect 16439 27557 16451 27560
rect 16393 27551 16451 27557
rect 20073 27557 20085 27591
rect 20119 27588 20131 27591
rect 21082 27588 21088 27600
rect 20119 27560 21088 27588
rect 20119 27557 20131 27560
rect 20073 27551 20131 27557
rect 21082 27548 21088 27560
rect 21140 27548 21146 27600
rect 24302 27548 24308 27600
rect 24360 27588 24366 27600
rect 25133 27591 25191 27597
rect 25133 27588 25145 27591
rect 24360 27560 25145 27588
rect 24360 27548 24366 27560
rect 25133 27557 25145 27560
rect 25179 27557 25191 27591
rect 25133 27551 25191 27557
rect 6181 27523 6239 27529
rect 6181 27489 6193 27523
rect 6227 27520 6239 27523
rect 6546 27520 6552 27532
rect 6227 27492 6552 27520
rect 6227 27489 6239 27492
rect 6181 27483 6239 27489
rect 6546 27480 6552 27492
rect 6604 27480 6610 27532
rect 7006 27480 7012 27532
rect 7064 27520 7070 27532
rect 8297 27523 8355 27529
rect 8297 27520 8309 27523
rect 7064 27492 8309 27520
rect 7064 27480 7070 27492
rect 8297 27489 8309 27492
rect 8343 27520 8355 27523
rect 8389 27523 8447 27529
rect 8389 27520 8401 27523
rect 8343 27492 8401 27520
rect 8343 27489 8355 27492
rect 8297 27483 8355 27489
rect 8389 27489 8401 27492
rect 8435 27520 8447 27523
rect 9030 27520 9036 27532
rect 8435 27492 9036 27520
rect 8435 27489 8447 27492
rect 8389 27483 8447 27489
rect 9030 27480 9036 27492
rect 9088 27480 9094 27532
rect 12802 27480 12808 27532
rect 12860 27520 12866 27532
rect 15657 27523 15715 27529
rect 15657 27520 15669 27523
rect 12860 27492 15669 27520
rect 12860 27480 12866 27492
rect 15657 27489 15669 27492
rect 15703 27489 15715 27523
rect 15657 27483 15715 27489
rect 17862 27480 17868 27532
rect 17920 27520 17926 27532
rect 17920 27492 19840 27520
rect 17920 27480 17926 27492
rect 9950 27412 9956 27464
rect 10008 27452 10014 27464
rect 10962 27452 10968 27464
rect 10008 27424 10968 27452
rect 10008 27412 10014 27424
rect 10962 27412 10968 27424
rect 11020 27452 11026 27464
rect 11149 27455 11207 27461
rect 11149 27452 11161 27455
rect 11020 27424 11161 27452
rect 11020 27412 11026 27424
rect 11149 27421 11161 27424
rect 11195 27421 11207 27455
rect 11149 27415 11207 27421
rect 13354 27412 13360 27464
rect 13412 27412 13418 27464
rect 14550 27412 14556 27464
rect 14608 27452 14614 27464
rect 18325 27455 18383 27461
rect 18325 27452 18337 27455
rect 14608 27424 18337 27452
rect 14608 27412 14614 27424
rect 18325 27421 18337 27424
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 7006 27344 7012 27396
rect 7064 27344 7070 27396
rect 11422 27344 11428 27396
rect 11480 27344 11486 27396
rect 13078 27384 13084 27396
rect 12650 27356 13084 27384
rect 13078 27344 13084 27356
rect 13136 27384 13142 27396
rect 13265 27387 13323 27393
rect 13265 27384 13277 27387
rect 13136 27356 13277 27384
rect 13136 27344 13142 27356
rect 13265 27353 13277 27356
rect 13311 27384 13323 27387
rect 13372 27384 13400 27412
rect 13906 27384 13912 27396
rect 13311 27356 13912 27384
rect 13311 27353 13323 27356
rect 13265 27347 13323 27353
rect 13906 27344 13912 27356
rect 13964 27384 13970 27396
rect 15194 27384 15200 27396
rect 13964 27356 15200 27384
rect 13964 27344 13970 27356
rect 15194 27344 15200 27356
rect 15252 27344 15258 27396
rect 15378 27344 15384 27396
rect 15436 27384 15442 27396
rect 15565 27387 15623 27393
rect 15565 27384 15577 27387
rect 15436 27356 15577 27384
rect 15436 27344 15442 27356
rect 15565 27353 15577 27356
rect 15611 27384 15623 27387
rect 16117 27387 16175 27393
rect 16117 27384 16129 27387
rect 15611 27356 16129 27384
rect 15611 27353 15623 27356
rect 15565 27347 15623 27353
rect 16117 27353 16129 27356
rect 16163 27384 16175 27387
rect 17218 27384 17224 27396
rect 16163 27356 17224 27384
rect 16163 27353 16175 27356
rect 16117 27347 16175 27353
rect 17218 27344 17224 27356
rect 17276 27384 17282 27396
rect 18877 27387 18935 27393
rect 18877 27384 18889 27387
rect 17276 27356 18889 27384
rect 17276 27344 17282 27356
rect 18877 27353 18889 27356
rect 18923 27384 18935 27387
rect 19518 27384 19524 27396
rect 18923 27356 19524 27384
rect 18923 27353 18935 27356
rect 18877 27347 18935 27353
rect 19518 27344 19524 27356
rect 19576 27344 19582 27396
rect 11698 27276 11704 27328
rect 11756 27316 11762 27328
rect 12894 27316 12900 27328
rect 11756 27288 12900 27316
rect 11756 27276 11762 27288
rect 12894 27276 12900 27288
rect 12952 27276 12958 27328
rect 13354 27276 13360 27328
rect 13412 27316 13418 27328
rect 13538 27316 13544 27328
rect 13412 27288 13544 27316
rect 13412 27276 13418 27288
rect 13538 27276 13544 27288
rect 13596 27276 13602 27328
rect 15010 27276 15016 27328
rect 15068 27316 15074 27328
rect 15105 27319 15163 27325
rect 15105 27316 15117 27319
rect 15068 27288 15117 27316
rect 15068 27276 15074 27288
rect 15105 27285 15117 27288
rect 15151 27285 15163 27319
rect 15105 27279 15163 27285
rect 15473 27319 15531 27325
rect 15473 27285 15485 27319
rect 15519 27316 15531 27319
rect 15838 27316 15844 27328
rect 15519 27288 15844 27316
rect 15519 27285 15531 27288
rect 15473 27279 15531 27285
rect 15838 27276 15844 27288
rect 15896 27276 15902 27328
rect 18141 27319 18199 27325
rect 18141 27285 18153 27319
rect 18187 27316 18199 27319
rect 18598 27316 18604 27328
rect 18187 27288 18604 27316
rect 18187 27285 18199 27288
rect 18141 27279 18199 27285
rect 18598 27276 18604 27288
rect 18656 27276 18662 27328
rect 19812 27325 19840 27492
rect 20530 27480 20536 27532
rect 20588 27520 20594 27532
rect 20625 27523 20683 27529
rect 20625 27520 20637 27523
rect 20588 27492 20637 27520
rect 20588 27480 20594 27492
rect 20625 27489 20637 27492
rect 20671 27489 20683 27523
rect 20625 27483 20683 27489
rect 21910 27480 21916 27532
rect 21968 27480 21974 27532
rect 23382 27480 23388 27532
rect 23440 27480 23446 27532
rect 20438 27412 20444 27464
rect 20496 27412 20502 27464
rect 23400 27452 23428 27480
rect 24320 27452 24348 27548
rect 23322 27424 24348 27452
rect 24486 27412 24492 27464
rect 24544 27452 24550 27464
rect 24673 27455 24731 27461
rect 24673 27452 24685 27455
rect 24544 27424 24685 27452
rect 24544 27412 24550 27424
rect 24673 27421 24685 27424
rect 24719 27421 24731 27455
rect 24673 27415 24731 27421
rect 20456 27384 20484 27412
rect 20533 27387 20591 27393
rect 20533 27384 20545 27387
rect 20456 27356 20545 27384
rect 20533 27353 20545 27356
rect 20579 27353 20591 27387
rect 20533 27347 20591 27353
rect 22186 27344 22192 27396
rect 22244 27344 22250 27396
rect 24857 27387 24915 27393
rect 24857 27353 24869 27387
rect 24903 27384 24915 27387
rect 25222 27384 25228 27396
rect 24903 27356 25228 27384
rect 24903 27353 24915 27356
rect 24857 27347 24915 27353
rect 25222 27344 25228 27356
rect 25280 27344 25286 27396
rect 19797 27319 19855 27325
rect 19797 27285 19809 27319
rect 19843 27316 19855 27319
rect 20441 27319 20499 27325
rect 20441 27316 20453 27319
rect 19843 27288 20453 27316
rect 19843 27285 19855 27288
rect 19797 27279 19855 27285
rect 20441 27285 20453 27288
rect 20487 27285 20499 27319
rect 20441 27279 20499 27285
rect 23106 27276 23112 27328
rect 23164 27316 23170 27328
rect 23661 27319 23719 27325
rect 23661 27316 23673 27319
rect 23164 27288 23673 27316
rect 23164 27276 23170 27288
rect 23661 27285 23673 27288
rect 23707 27285 23719 27319
rect 23661 27279 23719 27285
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 3191 27115 3249 27121
rect 3191 27081 3203 27115
rect 3237 27112 3249 27115
rect 3878 27112 3884 27124
rect 3237 27084 3884 27112
rect 3237 27081 3249 27084
rect 3191 27075 3249 27081
rect 3878 27072 3884 27084
rect 3936 27072 3942 27124
rect 6472 27084 10916 27112
rect 3120 26979 3178 26985
rect 3120 26945 3132 26979
rect 3166 26976 3178 26979
rect 3326 26976 3332 26988
rect 3166 26948 3332 26976
rect 3166 26945 3178 26948
rect 3120 26939 3178 26945
rect 3326 26936 3332 26948
rect 3384 26936 3390 26988
rect 3510 26936 3516 26988
rect 3568 26976 3574 26988
rect 3697 26979 3755 26985
rect 3697 26976 3709 26979
rect 3568 26948 3709 26976
rect 3568 26936 3574 26948
rect 3697 26945 3709 26948
rect 3743 26945 3755 26979
rect 3697 26939 3755 26945
rect 3881 26911 3939 26917
rect 3881 26877 3893 26911
rect 3927 26908 3939 26911
rect 4338 26908 4344 26920
rect 3927 26880 4344 26908
rect 3927 26877 3939 26880
rect 3881 26871 3939 26877
rect 4338 26868 4344 26880
rect 4396 26868 4402 26920
rect 4433 26911 4491 26917
rect 4433 26877 4445 26911
rect 4479 26908 4491 26911
rect 6472 26908 6500 27084
rect 7098 27004 7104 27056
rect 7156 27044 7162 27056
rect 7156 27016 7314 27044
rect 7156 27004 7162 27016
rect 10502 27004 10508 27056
rect 10560 27004 10566 27056
rect 6546 26936 6552 26988
rect 6604 26936 6610 26988
rect 9122 26936 9128 26988
rect 9180 26936 9186 26988
rect 4479 26880 6500 26908
rect 6825 26911 6883 26917
rect 4479 26877 4491 26880
rect 4433 26871 4491 26877
rect 6825 26877 6837 26911
rect 6871 26908 6883 26911
rect 7834 26908 7840 26920
rect 6871 26880 7840 26908
rect 6871 26877 6883 26880
rect 6825 26871 6883 26877
rect 4448 26840 4476 26871
rect 7834 26868 7840 26880
rect 7892 26868 7898 26920
rect 8938 26868 8944 26920
rect 8996 26908 9002 26920
rect 9217 26911 9275 26917
rect 9217 26908 9229 26911
rect 8996 26880 9229 26908
rect 8996 26868 9002 26880
rect 9217 26877 9229 26880
rect 9263 26877 9275 26911
rect 9217 26871 9275 26877
rect 9398 26868 9404 26920
rect 9456 26868 9462 26920
rect 10888 26908 10916 27084
rect 11054 27072 11060 27124
rect 11112 27112 11118 27124
rect 11514 27112 11520 27124
rect 11112 27084 11520 27112
rect 11112 27072 11118 27084
rect 11514 27072 11520 27084
rect 11572 27072 11578 27124
rect 11606 27072 11612 27124
rect 11664 27112 11670 27124
rect 12526 27112 12532 27124
rect 11664 27084 12532 27112
rect 11664 27072 11670 27084
rect 12526 27072 12532 27084
rect 12584 27072 12590 27124
rect 12894 27072 12900 27124
rect 12952 27112 12958 27124
rect 12952 27084 14136 27112
rect 12952 27072 12958 27084
rect 11330 27004 11336 27056
rect 11388 27044 11394 27056
rect 13078 27044 13084 27056
rect 11388 27016 13084 27044
rect 11388 27004 11394 27016
rect 13078 27004 13084 27016
rect 13136 27004 13142 27056
rect 14108 27044 14136 27084
rect 15102 27072 15108 27124
rect 15160 27112 15166 27124
rect 15197 27115 15255 27121
rect 15197 27112 15209 27115
rect 15160 27084 15209 27112
rect 15160 27072 15166 27084
rect 15197 27081 15209 27084
rect 15243 27081 15255 27115
rect 15197 27075 15255 27081
rect 17589 27115 17647 27121
rect 17589 27081 17601 27115
rect 17635 27112 17647 27115
rect 19981 27115 20039 27121
rect 19981 27112 19993 27115
rect 17635 27084 19993 27112
rect 17635 27081 17647 27084
rect 17589 27075 17647 27081
rect 19981 27081 19993 27084
rect 20027 27081 20039 27115
rect 24578 27112 24584 27124
rect 19981 27075 20039 27081
rect 22848 27084 24584 27112
rect 18049 27047 18107 27053
rect 14108 27016 15332 27044
rect 10962 26936 10968 26988
rect 11020 26976 11026 26988
rect 12529 26979 12587 26985
rect 12529 26976 12541 26979
rect 11020 26948 12541 26976
rect 11020 26936 11026 26948
rect 12529 26945 12541 26948
rect 12575 26945 12587 26979
rect 12529 26939 12587 26945
rect 13906 26936 13912 26988
rect 13964 26976 13970 26988
rect 14550 26976 14556 26988
rect 13964 26948 14556 26976
rect 13964 26936 13970 26948
rect 14550 26936 14556 26948
rect 14608 26936 14614 26988
rect 15105 26979 15163 26985
rect 15105 26945 15117 26979
rect 15151 26945 15163 26979
rect 15105 26939 15163 26945
rect 11606 26908 11612 26920
rect 10888 26880 11612 26908
rect 11606 26868 11612 26880
rect 11664 26868 11670 26920
rect 12802 26868 12808 26920
rect 12860 26868 12866 26920
rect 13538 26868 13544 26920
rect 13596 26908 13602 26920
rect 15120 26908 15148 26939
rect 15304 26917 15332 27016
rect 18049 27013 18061 27047
rect 18095 27044 18107 27047
rect 18414 27044 18420 27056
rect 18095 27016 18420 27044
rect 18095 27013 18107 27016
rect 18049 27007 18107 27013
rect 18414 27004 18420 27016
rect 18472 27004 18478 27056
rect 18598 27004 18604 27056
rect 18656 27044 18662 27056
rect 21726 27044 21732 27056
rect 18656 27016 21732 27044
rect 18656 27004 18662 27016
rect 21726 27004 21732 27016
rect 21784 27004 21790 27056
rect 17218 26936 17224 26988
rect 17276 26976 17282 26988
rect 17957 26979 18015 26985
rect 17957 26976 17969 26979
rect 17276 26948 17969 26976
rect 17276 26936 17282 26948
rect 17957 26945 17969 26948
rect 18003 26945 18015 26979
rect 17957 26939 18015 26945
rect 19889 26979 19947 26985
rect 19889 26945 19901 26979
rect 19935 26976 19947 26979
rect 20717 26979 20775 26985
rect 20717 26976 20729 26979
rect 19935 26948 20729 26976
rect 19935 26945 19947 26948
rect 19889 26939 19947 26945
rect 20717 26945 20729 26948
rect 20763 26945 20775 26979
rect 20717 26939 20775 26945
rect 22373 26979 22431 26985
rect 22373 26945 22385 26979
rect 22419 26976 22431 26979
rect 22848 26976 22876 27084
rect 24578 27072 24584 27084
rect 24636 27072 24642 27124
rect 23106 27004 23112 27056
rect 23164 27004 23170 27056
rect 23382 27004 23388 27056
rect 23440 27044 23446 27056
rect 23440 27016 23598 27044
rect 23440 27004 23446 27016
rect 25038 27004 25044 27056
rect 25096 27044 25102 27056
rect 25133 27047 25191 27053
rect 25133 27044 25145 27047
rect 25096 27016 25145 27044
rect 25096 27004 25102 27016
rect 25133 27013 25145 27016
rect 25179 27013 25191 27047
rect 25133 27007 25191 27013
rect 22419 26948 22876 26976
rect 22419 26945 22431 26948
rect 22373 26939 22431 26945
rect 13596 26880 15148 26908
rect 15289 26911 15347 26917
rect 13596 26868 13602 26880
rect 15289 26877 15301 26911
rect 15335 26877 15347 26911
rect 15289 26871 15347 26877
rect 18233 26911 18291 26917
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 19334 26908 19340 26920
rect 18279 26880 19340 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 19334 26868 19340 26880
rect 19392 26908 19398 26920
rect 19794 26908 19800 26920
rect 19392 26880 19800 26908
rect 19392 26868 19398 26880
rect 19794 26868 19800 26880
rect 19852 26868 19858 26920
rect 20165 26911 20223 26917
rect 20165 26877 20177 26911
rect 20211 26908 20223 26911
rect 21174 26908 21180 26920
rect 20211 26880 21180 26908
rect 20211 26877 20223 26880
rect 20165 26871 20223 26877
rect 21174 26868 21180 26880
rect 21232 26868 21238 26920
rect 22002 26868 22008 26920
rect 22060 26908 22066 26920
rect 22833 26911 22891 26917
rect 22833 26908 22845 26911
rect 22060 26880 22845 26908
rect 22060 26868 22066 26880
rect 22833 26877 22845 26880
rect 22879 26877 22891 26911
rect 23106 26908 23112 26920
rect 22833 26871 22891 26877
rect 22940 26880 23112 26908
rect 3896 26812 4476 26840
rect 3896 26784 3924 26812
rect 8294 26800 8300 26852
rect 8352 26840 8358 26852
rect 9674 26840 9680 26852
rect 8352 26812 9680 26840
rect 8352 26800 8358 26812
rect 9674 26800 9680 26812
rect 9732 26800 9738 26852
rect 10226 26800 10232 26852
rect 10284 26840 10290 26852
rect 10689 26843 10747 26849
rect 10689 26840 10701 26843
rect 10284 26812 10701 26840
rect 10284 26800 10290 26812
rect 10689 26809 10701 26812
rect 10735 26809 10747 26843
rect 10689 26803 10747 26809
rect 14737 26843 14795 26849
rect 14737 26809 14749 26843
rect 14783 26840 14795 26843
rect 17402 26840 17408 26852
rect 14783 26812 17408 26840
rect 14783 26809 14795 26812
rect 14737 26803 14795 26809
rect 17402 26800 17408 26812
rect 17460 26800 17466 26852
rect 20530 26800 20536 26852
rect 20588 26840 20594 26852
rect 22940 26840 22968 26880
rect 23106 26868 23112 26880
rect 23164 26868 23170 26920
rect 23198 26868 23204 26920
rect 23256 26908 23262 26920
rect 25317 26911 25375 26917
rect 25317 26908 25329 26911
rect 23256 26880 25329 26908
rect 23256 26868 23262 26880
rect 25317 26877 25329 26880
rect 25363 26877 25375 26911
rect 25317 26871 25375 26877
rect 20588 26812 22968 26840
rect 20588 26800 20594 26812
rect 3878 26732 3884 26784
rect 3936 26732 3942 26784
rect 8757 26775 8815 26781
rect 8757 26741 8769 26775
rect 8803 26772 8815 26775
rect 10502 26772 10508 26784
rect 8803 26744 10508 26772
rect 8803 26741 8815 26744
rect 8757 26735 8815 26741
rect 10502 26732 10508 26744
rect 10560 26732 10566 26784
rect 11330 26732 11336 26784
rect 11388 26772 11394 26784
rect 11793 26775 11851 26781
rect 11793 26772 11805 26775
rect 11388 26744 11805 26772
rect 11388 26732 11394 26744
rect 11793 26741 11805 26744
rect 11839 26741 11851 26775
rect 11793 26735 11851 26741
rect 14277 26775 14335 26781
rect 14277 26741 14289 26775
rect 14323 26772 14335 26775
rect 14366 26772 14372 26784
rect 14323 26744 14372 26772
rect 14323 26741 14335 26744
rect 14277 26735 14335 26741
rect 14366 26732 14372 26744
rect 14424 26732 14430 26784
rect 17218 26732 17224 26784
rect 17276 26732 17282 26784
rect 19518 26732 19524 26784
rect 19576 26732 19582 26784
rect 22189 26775 22247 26781
rect 22189 26741 22201 26775
rect 22235 26772 22247 26775
rect 23842 26772 23848 26784
rect 22235 26744 23848 26772
rect 22235 26741 22247 26744
rect 22189 26735 22247 26741
rect 23842 26732 23848 26744
rect 23900 26732 23906 26784
rect 24578 26732 24584 26784
rect 24636 26732 24642 26784
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 4062 26528 4068 26580
rect 4120 26528 4126 26580
rect 8570 26528 8576 26580
rect 8628 26568 8634 26580
rect 11701 26571 11759 26577
rect 11701 26568 11713 26571
rect 8628 26540 11713 26568
rect 8628 26528 8634 26540
rect 11701 26537 11713 26540
rect 11747 26568 11759 26571
rect 13630 26568 13636 26580
rect 11747 26540 13636 26568
rect 11747 26537 11759 26540
rect 11701 26531 11759 26537
rect 13630 26528 13636 26540
rect 13688 26528 13694 26580
rect 16666 26528 16672 26580
rect 16724 26568 16730 26580
rect 17129 26571 17187 26577
rect 17129 26568 17141 26571
rect 16724 26540 17141 26568
rect 16724 26528 16730 26540
rect 17129 26537 17141 26540
rect 17175 26568 17187 26571
rect 17770 26568 17776 26580
rect 17175 26540 17776 26568
rect 17175 26537 17187 26540
rect 17129 26531 17187 26537
rect 17770 26528 17776 26540
rect 17828 26528 17834 26580
rect 22186 26528 22192 26580
rect 22244 26568 22250 26580
rect 22373 26571 22431 26577
rect 22373 26568 22385 26571
rect 22244 26540 22385 26568
rect 22244 26528 22250 26540
rect 22373 26537 22385 26540
rect 22419 26537 22431 26571
rect 22373 26531 22431 26537
rect 22646 26528 22652 26580
rect 22704 26568 22710 26580
rect 24578 26568 24584 26580
rect 22704 26540 24584 26568
rect 22704 26528 22710 26540
rect 24578 26528 24584 26540
rect 24636 26528 24642 26580
rect 16758 26460 16764 26512
rect 16816 26500 16822 26512
rect 18414 26500 18420 26512
rect 16816 26472 18420 26500
rect 16816 26460 16822 26472
rect 18414 26460 18420 26472
rect 18472 26460 18478 26512
rect 19429 26503 19487 26509
rect 19429 26469 19441 26503
rect 19475 26500 19487 26503
rect 19702 26500 19708 26512
rect 19475 26472 19708 26500
rect 19475 26469 19487 26472
rect 19429 26463 19487 26469
rect 19702 26460 19708 26472
rect 19760 26460 19766 26512
rect 22002 26500 22008 26512
rect 21928 26472 22008 26500
rect 6454 26392 6460 26444
rect 6512 26392 6518 26444
rect 6733 26435 6791 26441
rect 6733 26401 6745 26435
rect 6779 26432 6791 26435
rect 8294 26432 8300 26444
rect 6779 26404 8300 26432
rect 6779 26401 6791 26404
rect 6733 26395 6791 26401
rect 8294 26392 8300 26404
rect 8352 26392 8358 26444
rect 9122 26392 9128 26444
rect 9180 26392 9186 26444
rect 10229 26435 10287 26441
rect 10229 26401 10241 26435
rect 10275 26432 10287 26435
rect 11698 26432 11704 26444
rect 10275 26404 11704 26432
rect 10275 26401 10287 26404
rect 10229 26395 10287 26401
rect 11698 26392 11704 26404
rect 11756 26392 11762 26444
rect 11790 26392 11796 26444
rect 11848 26432 11854 26444
rect 12713 26435 12771 26441
rect 12713 26432 12725 26435
rect 11848 26404 12725 26432
rect 11848 26392 11854 26404
rect 12713 26401 12725 26404
rect 12759 26401 12771 26435
rect 12713 26395 12771 26401
rect 15657 26435 15715 26441
rect 15657 26401 15669 26435
rect 15703 26432 15715 26435
rect 17586 26432 17592 26444
rect 15703 26404 17592 26432
rect 15703 26401 15715 26404
rect 15657 26395 15715 26401
rect 17586 26392 17592 26404
rect 17644 26392 17650 26444
rect 18966 26392 18972 26444
rect 19024 26432 19030 26444
rect 19889 26435 19947 26441
rect 19889 26432 19901 26435
rect 19024 26404 19901 26432
rect 19024 26392 19030 26404
rect 19889 26401 19901 26404
rect 19935 26401 19947 26435
rect 19889 26395 19947 26401
rect 20073 26435 20131 26441
rect 20073 26401 20085 26435
rect 20119 26432 20131 26435
rect 20254 26432 20260 26444
rect 20119 26404 20260 26432
rect 20119 26401 20131 26404
rect 20073 26395 20131 26401
rect 20254 26392 20260 26404
rect 20312 26392 20318 26444
rect 20625 26435 20683 26441
rect 20625 26401 20637 26435
rect 20671 26432 20683 26435
rect 21928 26432 21956 26472
rect 22002 26460 22008 26472
rect 22060 26460 22066 26512
rect 22554 26460 22560 26512
rect 22612 26500 22618 26512
rect 22833 26503 22891 26509
rect 22833 26500 22845 26503
rect 22612 26472 22845 26500
rect 22612 26460 22618 26472
rect 22833 26469 22845 26472
rect 22879 26469 22891 26503
rect 22833 26463 22891 26469
rect 23382 26460 23388 26512
rect 23440 26500 23446 26512
rect 23845 26503 23903 26509
rect 23845 26500 23857 26503
rect 23440 26472 23857 26500
rect 23440 26460 23446 26472
rect 23845 26469 23857 26472
rect 23891 26500 23903 26503
rect 24946 26500 24952 26512
rect 23891 26472 24952 26500
rect 23891 26469 23903 26472
rect 23845 26463 23903 26469
rect 24946 26460 24952 26472
rect 25004 26500 25010 26512
rect 25133 26503 25191 26509
rect 25133 26500 25145 26503
rect 25004 26472 25145 26500
rect 25004 26460 25010 26472
rect 25133 26469 25145 26472
rect 25179 26469 25191 26503
rect 25133 26463 25191 26469
rect 20671 26404 21956 26432
rect 20671 26401 20683 26404
rect 20625 26395 20683 26401
rect 22462 26392 22468 26444
rect 22520 26432 22526 26444
rect 23293 26435 23351 26441
rect 23293 26432 23305 26435
rect 22520 26404 23305 26432
rect 22520 26392 22526 26404
rect 23293 26401 23305 26404
rect 23339 26401 23351 26435
rect 23293 26395 23351 26401
rect 23477 26435 23535 26441
rect 23477 26401 23489 26435
rect 23523 26432 23535 26435
rect 24578 26432 24584 26444
rect 23523 26404 24584 26432
rect 23523 26401 23535 26404
rect 23477 26395 23535 26401
rect 24578 26392 24584 26404
rect 24636 26392 24642 26444
rect 1765 26367 1823 26373
rect 1765 26333 1777 26367
rect 1811 26364 1823 26367
rect 2038 26364 2044 26376
rect 1811 26336 2044 26364
rect 1811 26333 1823 26336
rect 1765 26327 1823 26333
rect 2038 26324 2044 26336
rect 2096 26324 2102 26376
rect 9950 26324 9956 26376
rect 10008 26324 10014 26376
rect 11330 26324 11336 26376
rect 11388 26324 11394 26376
rect 12621 26367 12679 26373
rect 12621 26333 12633 26367
rect 12667 26364 12679 26367
rect 14274 26364 14280 26376
rect 12667 26336 14280 26364
rect 12667 26333 12679 26336
rect 12621 26327 12679 26333
rect 14274 26324 14280 26336
rect 14332 26324 14338 26376
rect 15378 26324 15384 26376
rect 15436 26324 15442 26376
rect 22034 26336 22094 26364
rect 2774 26256 2780 26308
rect 2832 26256 2838 26308
rect 8665 26299 8723 26305
rect 7116 26268 7222 26296
rect 7116 26240 7144 26268
rect 8665 26265 8677 26299
rect 8711 26296 8723 26299
rect 8938 26296 8944 26308
rect 8711 26268 8944 26296
rect 8711 26265 8723 26268
rect 8665 26259 8723 26265
rect 8938 26256 8944 26268
rect 8996 26256 9002 26308
rect 13722 26296 13728 26308
rect 12176 26268 13728 26296
rect 7098 26188 7104 26240
rect 7156 26188 7162 26240
rect 7650 26188 7656 26240
rect 7708 26228 7714 26240
rect 12176 26237 12204 26268
rect 13722 26256 13728 26268
rect 13780 26256 13786 26308
rect 17405 26299 17463 26305
rect 17405 26296 17417 26299
rect 16882 26268 17417 26296
rect 17405 26265 17417 26268
rect 17451 26265 17463 26299
rect 17405 26259 17463 26265
rect 19797 26299 19855 26305
rect 19797 26265 19809 26299
rect 19843 26296 19855 26299
rect 20622 26296 20628 26308
rect 19843 26268 20628 26296
rect 19843 26265 19855 26268
rect 19797 26259 19855 26265
rect 8205 26231 8263 26237
rect 8205 26228 8217 26231
rect 7708 26200 8217 26228
rect 7708 26188 7714 26200
rect 8205 26197 8217 26200
rect 8251 26197 8263 26231
rect 8205 26191 8263 26197
rect 12161 26231 12219 26237
rect 12161 26197 12173 26231
rect 12207 26197 12219 26231
rect 12161 26191 12219 26197
rect 12526 26188 12532 26240
rect 12584 26188 12590 26240
rect 14461 26231 14519 26237
rect 14461 26197 14473 26231
rect 14507 26228 14519 26231
rect 14550 26228 14556 26240
rect 14507 26200 14556 26228
rect 14507 26197 14519 26200
rect 14461 26191 14519 26197
rect 14550 26188 14556 26200
rect 14608 26188 14614 26240
rect 17218 26188 17224 26240
rect 17276 26228 17282 26240
rect 17420 26228 17448 26259
rect 20622 26256 20628 26268
rect 20680 26256 20686 26308
rect 20901 26299 20959 26305
rect 20901 26265 20913 26299
rect 20947 26296 20959 26299
rect 21174 26296 21180 26308
rect 20947 26268 21180 26296
rect 20947 26265 20959 26268
rect 20901 26259 20959 26265
rect 21174 26256 21180 26268
rect 21232 26256 21238 26308
rect 22066 26296 22094 26336
rect 22278 26324 22284 26376
rect 22336 26364 22342 26376
rect 23201 26367 23259 26373
rect 23201 26364 23213 26367
rect 22336 26336 23213 26364
rect 22336 26324 22342 26336
rect 23201 26333 23213 26336
rect 23247 26333 23259 26367
rect 23201 26327 23259 26333
rect 24394 26324 24400 26376
rect 24452 26364 24458 26376
rect 24673 26367 24731 26373
rect 24673 26364 24685 26367
rect 24452 26336 24685 26364
rect 24452 26324 24458 26336
rect 24673 26333 24685 26336
rect 24719 26333 24731 26367
rect 24673 26327 24731 26333
rect 23382 26296 23388 26308
rect 22066 26268 23388 26296
rect 17276 26200 17448 26228
rect 17276 26188 17282 26200
rect 20990 26188 20996 26240
rect 21048 26228 21054 26240
rect 22066 26228 22094 26268
rect 23382 26256 23388 26268
rect 23440 26256 23446 26308
rect 24857 26299 24915 26305
rect 24857 26265 24869 26299
rect 24903 26296 24915 26299
rect 25222 26296 25228 26308
rect 24903 26268 25228 26296
rect 24903 26265 24915 26268
rect 24857 26259 24915 26265
rect 25038 26256 25044 26268
rect 25096 26256 25102 26308
rect 21048 26200 22094 26228
rect 21048 26188 21054 26200
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 1762 25984 1768 26036
rect 1820 26024 1826 26036
rect 2133 26027 2191 26033
rect 2133 26024 2145 26027
rect 1820 25996 2145 26024
rect 1820 25984 1826 25996
rect 2133 25993 2145 25996
rect 2179 25993 2191 26027
rect 2133 25987 2191 25993
rect 7098 25984 7104 26036
rect 7156 26024 7162 26036
rect 8481 26027 8539 26033
rect 8481 26024 8493 26027
rect 7156 25996 8493 26024
rect 7156 25984 7162 25996
rect 8481 25993 8493 25996
rect 8527 26024 8539 26027
rect 8846 26024 8852 26036
rect 8527 25996 8852 26024
rect 8527 25993 8539 25996
rect 8481 25987 8539 25993
rect 8846 25984 8852 25996
rect 8904 25984 8910 26036
rect 9217 26027 9275 26033
rect 9217 25993 9229 26027
rect 9263 25993 9275 26027
rect 9217 25987 9275 25993
rect 3510 25916 3516 25968
rect 3568 25956 3574 25968
rect 4062 25956 4068 25968
rect 3568 25928 4068 25956
rect 3568 25916 3574 25928
rect 4062 25916 4068 25928
rect 4120 25956 4126 25968
rect 9232 25956 9260 25987
rect 10502 25984 10508 26036
rect 10560 26024 10566 26036
rect 10781 26027 10839 26033
rect 10781 26024 10793 26027
rect 10560 25996 10793 26024
rect 10560 25984 10566 25996
rect 10781 25993 10793 25996
rect 10827 25993 10839 26027
rect 10781 25987 10839 25993
rect 10870 25984 10876 26036
rect 10928 25984 10934 26036
rect 15378 26024 15384 26036
rect 12728 25996 15384 26024
rect 12526 25956 12532 25968
rect 4120 25928 4200 25956
rect 9232 25928 12532 25956
rect 4120 25916 4126 25928
rect 2317 25891 2375 25897
rect 2317 25857 2329 25891
rect 2363 25888 2375 25891
rect 2866 25888 2872 25900
rect 2363 25860 2872 25888
rect 2363 25857 2375 25860
rect 2317 25851 2375 25857
rect 2866 25848 2872 25860
rect 2924 25848 2930 25900
rect 4172 25897 4200 25928
rect 12526 25916 12532 25928
rect 12584 25916 12590 25968
rect 3053 25891 3111 25897
rect 3053 25857 3065 25891
rect 3099 25888 3111 25891
rect 4157 25891 4215 25897
rect 3099 25860 4108 25888
rect 3099 25857 3111 25860
rect 3053 25851 3111 25857
rect 2774 25780 2780 25832
rect 2832 25820 2838 25832
rect 3237 25823 3295 25829
rect 3237 25820 3249 25823
rect 2832 25792 3249 25820
rect 2832 25780 2838 25792
rect 3237 25789 3249 25792
rect 3283 25820 3295 25823
rect 3602 25820 3608 25832
rect 3283 25792 3608 25820
rect 3283 25789 3295 25792
rect 3237 25783 3295 25789
rect 3602 25780 3608 25792
rect 3660 25780 3666 25832
rect 4080 25820 4108 25860
rect 4157 25857 4169 25891
rect 4203 25857 4215 25891
rect 4157 25851 4215 25857
rect 4798 25848 4804 25900
rect 4856 25888 4862 25900
rect 8478 25888 8484 25900
rect 4856 25860 8484 25888
rect 4856 25848 4862 25860
rect 8478 25848 8484 25860
rect 8536 25888 8542 25900
rect 8849 25891 8907 25897
rect 8849 25888 8861 25891
rect 8536 25860 8861 25888
rect 8536 25848 8542 25860
rect 8849 25857 8861 25860
rect 8895 25857 8907 25891
rect 8849 25851 8907 25857
rect 6178 25820 6184 25832
rect 4080 25792 6184 25820
rect 6178 25780 6184 25792
rect 6236 25780 6242 25832
rect 7834 25780 7840 25832
rect 7892 25820 7898 25832
rect 8021 25823 8079 25829
rect 8021 25820 8033 25823
rect 7892 25792 8033 25820
rect 7892 25780 7898 25792
rect 8021 25789 8033 25792
rect 8067 25789 8079 25823
rect 8864 25820 8892 25851
rect 9398 25848 9404 25900
rect 9456 25888 9462 25900
rect 12728 25897 12756 25996
rect 15378 25984 15384 25996
rect 15436 25984 15442 26036
rect 15562 25984 15568 26036
rect 15620 26024 15626 26036
rect 15841 26027 15899 26033
rect 15841 26024 15853 26027
rect 15620 25996 15853 26024
rect 15620 25984 15626 25996
rect 15841 25993 15853 25996
rect 15887 25993 15899 26027
rect 15841 25987 15899 25993
rect 19334 25984 19340 26036
rect 19392 25984 19398 26036
rect 19518 25984 19524 26036
rect 19576 26024 19582 26036
rect 20257 26027 20315 26033
rect 20257 26024 20269 26027
rect 19576 25996 20269 26024
rect 19576 25984 19582 25996
rect 20257 25993 20269 25996
rect 20303 25993 20315 26027
rect 20257 25987 20315 25993
rect 20346 25984 20352 26036
rect 20404 25984 20410 26036
rect 22370 25984 22376 26036
rect 22428 25984 22434 26036
rect 22465 26027 22523 26033
rect 22465 25993 22477 26027
rect 22511 26024 22523 26027
rect 22738 26024 22744 26036
rect 22511 25996 22744 26024
rect 22511 25993 22523 25996
rect 22465 25987 22523 25993
rect 22738 25984 22744 25996
rect 22796 25984 22802 26036
rect 14550 25956 14556 25968
rect 14214 25928 14556 25956
rect 14550 25916 14556 25928
rect 14608 25916 14614 25968
rect 15396 25956 15424 25984
rect 15396 25928 17632 25956
rect 9585 25891 9643 25897
rect 9585 25888 9597 25891
rect 9456 25860 9597 25888
rect 9456 25848 9462 25860
rect 9585 25857 9597 25860
rect 9631 25857 9643 25891
rect 9585 25851 9643 25857
rect 12713 25891 12771 25897
rect 12713 25857 12725 25891
rect 12759 25857 12771 25891
rect 12713 25851 12771 25857
rect 15749 25891 15807 25897
rect 15749 25857 15761 25891
rect 15795 25888 15807 25891
rect 17494 25888 17500 25900
rect 15795 25860 17500 25888
rect 15795 25857 15807 25860
rect 15749 25851 15807 25857
rect 17494 25848 17500 25860
rect 17552 25848 17558 25900
rect 17604 25897 17632 25928
rect 20070 25916 20076 25968
rect 20128 25956 20134 25968
rect 23293 25959 23351 25965
rect 23293 25956 23305 25959
rect 20128 25928 23305 25956
rect 20128 25916 20134 25928
rect 23293 25925 23305 25928
rect 23339 25925 23351 25959
rect 23293 25919 23351 25925
rect 17589 25891 17647 25897
rect 17589 25857 17601 25891
rect 17635 25857 17647 25891
rect 22186 25888 22192 25900
rect 18998 25874 20024 25888
rect 17589 25851 17647 25857
rect 18984 25860 20024 25874
rect 9677 25823 9735 25829
rect 9677 25820 9689 25823
rect 8864 25792 9689 25820
rect 8021 25783 8079 25789
rect 9677 25789 9689 25792
rect 9723 25789 9735 25823
rect 9677 25783 9735 25789
rect 9769 25823 9827 25829
rect 9769 25789 9781 25823
rect 9815 25789 9827 25823
rect 9769 25783 9827 25789
rect 3418 25712 3424 25764
rect 3476 25712 3482 25764
rect 3620 25752 3648 25780
rect 4617 25755 4675 25761
rect 4617 25752 4629 25755
rect 3620 25724 4629 25752
rect 4617 25721 4629 25724
rect 4663 25721 4675 25755
rect 4617 25715 4675 25721
rect 8570 25712 8576 25764
rect 8628 25752 8634 25764
rect 9784 25752 9812 25783
rect 9858 25780 9864 25832
rect 9916 25820 9922 25832
rect 10965 25823 11023 25829
rect 10965 25820 10977 25823
rect 9916 25792 10977 25820
rect 9916 25780 9922 25792
rect 10965 25789 10977 25792
rect 11011 25789 11023 25823
rect 10965 25783 11023 25789
rect 11790 25780 11796 25832
rect 11848 25820 11854 25832
rect 11977 25823 12035 25829
rect 11977 25820 11989 25823
rect 11848 25792 11989 25820
rect 11848 25780 11854 25792
rect 11977 25789 11989 25792
rect 12023 25789 12035 25823
rect 11977 25783 12035 25789
rect 12342 25780 12348 25832
rect 12400 25820 12406 25832
rect 12526 25820 12532 25832
rect 12400 25792 12532 25820
rect 12400 25780 12406 25792
rect 12526 25780 12532 25792
rect 12584 25780 12590 25832
rect 12989 25823 13047 25829
rect 12989 25789 13001 25823
rect 13035 25820 13047 25823
rect 14366 25820 14372 25832
rect 13035 25792 14372 25820
rect 13035 25789 13047 25792
rect 12989 25783 13047 25789
rect 14366 25780 14372 25792
rect 14424 25780 14430 25832
rect 14461 25823 14519 25829
rect 14461 25789 14473 25823
rect 14507 25820 14519 25823
rect 14918 25820 14924 25832
rect 14507 25792 14924 25820
rect 14507 25789 14519 25792
rect 14461 25783 14519 25789
rect 8628 25724 9812 25752
rect 10413 25755 10471 25761
rect 8628 25712 8634 25724
rect 10413 25721 10425 25755
rect 10459 25752 10471 25755
rect 12250 25752 12256 25764
rect 10459 25724 12256 25752
rect 10459 25721 10471 25724
rect 10413 25715 10471 25721
rect 12250 25712 12256 25724
rect 12308 25712 12314 25764
rect 4246 25644 4252 25696
rect 4304 25644 4310 25696
rect 11422 25644 11428 25696
rect 11480 25684 11486 25696
rect 14476 25684 14504 25783
rect 14918 25780 14924 25792
rect 14976 25780 14982 25832
rect 16022 25780 16028 25832
rect 16080 25780 16086 25832
rect 17862 25780 17868 25832
rect 17920 25780 17926 25832
rect 18230 25780 18236 25832
rect 18288 25820 18294 25832
rect 18984 25820 19012 25860
rect 18288 25792 19012 25820
rect 18288 25780 18294 25792
rect 14550 25712 14556 25764
rect 14608 25752 14614 25764
rect 14829 25755 14887 25761
rect 14829 25752 14841 25755
rect 14608 25724 14841 25752
rect 14608 25712 14614 25724
rect 14829 25721 14841 25724
rect 14875 25752 14887 25755
rect 17218 25752 17224 25764
rect 14875 25724 17224 25752
rect 14875 25721 14887 25724
rect 14829 25715 14887 25721
rect 17218 25712 17224 25724
rect 17276 25712 17282 25764
rect 19889 25755 19947 25761
rect 19889 25752 19901 25755
rect 18892 25724 19901 25752
rect 18892 25696 18920 25724
rect 19889 25721 19901 25724
rect 19935 25721 19947 25755
rect 19996 25752 20024 25860
rect 20548 25860 22192 25888
rect 20548 25829 20576 25860
rect 22186 25848 22192 25860
rect 22244 25848 22250 25900
rect 23842 25848 23848 25900
rect 23900 25888 23906 25900
rect 23937 25891 23995 25897
rect 23937 25888 23949 25891
rect 23900 25860 23949 25888
rect 23900 25848 23906 25860
rect 23937 25857 23949 25860
rect 23983 25857 23995 25891
rect 23937 25851 23995 25857
rect 20533 25823 20591 25829
rect 20533 25789 20545 25823
rect 20579 25789 20591 25823
rect 20533 25783 20591 25789
rect 21269 25823 21327 25829
rect 21269 25789 21281 25823
rect 21315 25820 21327 25823
rect 21634 25820 21640 25832
rect 21315 25792 21640 25820
rect 21315 25789 21327 25792
rect 21269 25783 21327 25789
rect 21634 25780 21640 25792
rect 21692 25780 21698 25832
rect 22649 25823 22707 25829
rect 22649 25789 22661 25823
rect 22695 25820 22707 25823
rect 22738 25820 22744 25832
rect 22695 25792 22744 25820
rect 22695 25789 22707 25792
rect 22649 25783 22707 25789
rect 22738 25780 22744 25792
rect 22796 25780 22802 25832
rect 25130 25780 25136 25832
rect 25188 25780 25194 25832
rect 23477 25755 23535 25761
rect 19996 25724 21036 25752
rect 19889 25715 19947 25721
rect 21008 25696 21036 25724
rect 23477 25721 23489 25755
rect 23523 25752 23535 25755
rect 23750 25752 23756 25764
rect 23523 25724 23756 25752
rect 23523 25721 23535 25724
rect 23477 25715 23535 25721
rect 23750 25712 23756 25724
rect 23808 25712 23814 25764
rect 11480 25656 14504 25684
rect 11480 25644 11486 25656
rect 14918 25644 14924 25696
rect 14976 25684 14982 25696
rect 15381 25687 15439 25693
rect 15381 25684 15393 25687
rect 14976 25656 15393 25684
rect 14976 25644 14982 25656
rect 15381 25653 15393 25656
rect 15427 25653 15439 25687
rect 15381 25647 15439 25653
rect 18874 25644 18880 25696
rect 18932 25644 18938 25696
rect 20990 25644 20996 25696
rect 21048 25644 21054 25696
rect 21174 25644 21180 25696
rect 21232 25684 21238 25696
rect 22005 25687 22063 25693
rect 22005 25684 22017 25687
rect 21232 25656 22017 25684
rect 21232 25644 21238 25656
rect 22005 25653 22017 25656
rect 22051 25653 22063 25687
rect 22005 25647 22063 25653
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 7088 25483 7146 25489
rect 7088 25449 7100 25483
rect 7134 25480 7146 25483
rect 7466 25480 7472 25492
rect 7134 25452 7472 25480
rect 7134 25449 7146 25452
rect 7088 25443 7146 25449
rect 7466 25440 7472 25452
rect 7524 25480 7530 25492
rect 7650 25480 7656 25492
rect 7524 25452 7656 25480
rect 7524 25440 7530 25452
rect 7650 25440 7656 25452
rect 7708 25440 7714 25492
rect 8846 25440 8852 25492
rect 8904 25480 8910 25492
rect 8941 25483 8999 25489
rect 8941 25480 8953 25483
rect 8904 25452 8953 25480
rect 8904 25440 8910 25452
rect 8941 25449 8953 25452
rect 8987 25449 8999 25483
rect 8941 25443 8999 25449
rect 11425 25483 11483 25489
rect 11425 25449 11437 25483
rect 11471 25480 11483 25483
rect 13538 25480 13544 25492
rect 11471 25452 13544 25480
rect 11471 25449 11483 25452
rect 11425 25443 11483 25449
rect 13538 25440 13544 25452
rect 13596 25440 13602 25492
rect 14737 25483 14795 25489
rect 14737 25449 14749 25483
rect 14783 25480 14795 25483
rect 16758 25480 16764 25492
rect 14783 25452 16764 25480
rect 14783 25449 14795 25452
rect 14737 25443 14795 25449
rect 16758 25440 16764 25452
rect 16816 25440 16822 25492
rect 18049 25483 18107 25489
rect 18049 25449 18061 25483
rect 18095 25480 18107 25483
rect 18230 25480 18236 25492
rect 18095 25452 18236 25480
rect 18095 25449 18107 25452
rect 18049 25443 18107 25449
rect 10045 25415 10103 25421
rect 10045 25381 10057 25415
rect 10091 25412 10103 25415
rect 12250 25412 12256 25424
rect 10091 25384 12256 25412
rect 10091 25381 10103 25384
rect 10045 25375 10103 25381
rect 12250 25372 12256 25384
rect 12308 25372 12314 25424
rect 15304 25384 16068 25412
rect 6825 25347 6883 25353
rect 6825 25313 6837 25347
rect 6871 25344 6883 25347
rect 7650 25344 7656 25356
rect 6871 25316 7656 25344
rect 6871 25313 6883 25316
rect 6825 25307 6883 25313
rect 7650 25304 7656 25316
rect 7708 25304 7714 25356
rect 8570 25304 8576 25356
rect 8628 25304 8634 25356
rect 9398 25304 9404 25356
rect 9456 25304 9462 25356
rect 9674 25304 9680 25356
rect 9732 25344 9738 25356
rect 10597 25347 10655 25353
rect 10597 25344 10609 25347
rect 9732 25316 10609 25344
rect 9732 25304 9738 25316
rect 10597 25313 10609 25316
rect 10643 25313 10655 25347
rect 10597 25307 10655 25313
rect 11422 25304 11428 25356
rect 11480 25344 11486 25356
rect 11977 25347 12035 25353
rect 11977 25344 11989 25347
rect 11480 25316 11989 25344
rect 11480 25304 11486 25316
rect 11977 25313 11989 25316
rect 12023 25313 12035 25347
rect 11977 25307 12035 25313
rect 12802 25304 12808 25356
rect 12860 25344 12866 25356
rect 15304 25353 15332 25384
rect 13173 25347 13231 25353
rect 13173 25344 13185 25347
rect 12860 25316 13185 25344
rect 12860 25304 12866 25316
rect 13173 25313 13185 25316
rect 13219 25313 13231 25347
rect 13173 25307 13231 25313
rect 15289 25347 15347 25353
rect 15289 25313 15301 25347
rect 15335 25313 15347 25347
rect 15289 25307 15347 25313
rect 15378 25304 15384 25356
rect 15436 25344 15442 25356
rect 15933 25347 15991 25353
rect 15933 25344 15945 25347
rect 15436 25316 15945 25344
rect 15436 25304 15442 25316
rect 15933 25313 15945 25316
rect 15979 25313 15991 25347
rect 16040 25344 16068 25384
rect 16209 25347 16267 25353
rect 16209 25344 16221 25347
rect 16040 25316 16221 25344
rect 15933 25307 15991 25313
rect 16209 25313 16221 25316
rect 16255 25344 16267 25347
rect 16666 25344 16672 25356
rect 16255 25316 16672 25344
rect 16255 25313 16267 25316
rect 16209 25307 16267 25313
rect 16666 25304 16672 25316
rect 16724 25304 16730 25356
rect 4062 25285 4068 25288
rect 4040 25279 4068 25285
rect 4040 25245 4052 25279
rect 4040 25239 4068 25245
rect 4062 25236 4068 25239
rect 4120 25236 4126 25288
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25276 10563 25279
rect 10778 25276 10784 25288
rect 10551 25248 10784 25276
rect 10551 25245 10563 25248
rect 10505 25239 10563 25245
rect 10778 25236 10784 25248
rect 10836 25236 10842 25288
rect 11790 25236 11796 25288
rect 11848 25236 11854 25288
rect 17218 25236 17224 25288
rect 17276 25276 17282 25288
rect 18064 25276 18092 25443
rect 18230 25440 18236 25452
rect 18288 25440 18294 25492
rect 22830 25440 22836 25492
rect 22888 25480 22894 25492
rect 23109 25483 23167 25489
rect 23109 25480 23121 25483
rect 22888 25452 23121 25480
rect 22888 25440 22894 25452
rect 23109 25449 23121 25452
rect 23155 25449 23167 25483
rect 23109 25443 23167 25449
rect 24946 25440 24952 25492
rect 25004 25480 25010 25492
rect 25133 25483 25191 25489
rect 25133 25480 25145 25483
rect 25004 25452 25145 25480
rect 25004 25440 25010 25452
rect 25133 25449 25145 25452
rect 25179 25449 25191 25483
rect 25133 25443 25191 25449
rect 25498 25440 25504 25492
rect 25556 25440 25562 25492
rect 22097 25415 22155 25421
rect 22097 25381 22109 25415
rect 22143 25412 22155 25415
rect 24854 25412 24860 25424
rect 22143 25384 24860 25412
rect 22143 25381 22155 25384
rect 22097 25375 22155 25381
rect 24854 25372 24860 25384
rect 24912 25372 24918 25424
rect 19058 25304 19064 25356
rect 19116 25344 19122 25356
rect 19889 25347 19947 25353
rect 19889 25344 19901 25347
rect 19116 25316 19901 25344
rect 19116 25304 19122 25316
rect 19889 25313 19901 25316
rect 19935 25313 19947 25347
rect 19889 25307 19947 25313
rect 20070 25304 20076 25356
rect 20128 25304 20134 25356
rect 21082 25304 21088 25356
rect 21140 25344 21146 25356
rect 22557 25347 22615 25353
rect 22557 25344 22569 25347
rect 21140 25316 22569 25344
rect 21140 25304 21146 25316
rect 22557 25313 22569 25316
rect 22603 25313 22615 25347
rect 22557 25307 22615 25313
rect 22646 25304 22652 25356
rect 22704 25304 22710 25356
rect 24026 25304 24032 25356
rect 24084 25304 24090 25356
rect 17276 25248 18092 25276
rect 18233 25279 18291 25285
rect 17276 25236 17282 25248
rect 18233 25245 18245 25279
rect 18279 25276 18291 25279
rect 18322 25276 18328 25288
rect 18279 25248 18328 25276
rect 18279 25245 18291 25248
rect 18233 25239 18291 25245
rect 18322 25236 18328 25248
rect 18380 25236 18386 25288
rect 19426 25236 19432 25288
rect 19484 25276 19490 25288
rect 19797 25279 19855 25285
rect 19797 25276 19809 25279
rect 19484 25248 19809 25276
rect 19484 25236 19490 25248
rect 19797 25245 19809 25248
rect 19843 25245 19855 25279
rect 19797 25239 19855 25245
rect 21634 25236 21640 25288
rect 21692 25276 21698 25288
rect 22465 25279 22523 25285
rect 22465 25276 22477 25279
rect 21692 25248 22477 25276
rect 21692 25236 21698 25248
rect 22465 25245 22477 25248
rect 22511 25245 22523 25279
rect 22465 25239 22523 25245
rect 23845 25279 23903 25285
rect 23845 25245 23857 25279
rect 23891 25276 23903 25279
rect 23934 25276 23940 25288
rect 23891 25248 23940 25276
rect 23891 25245 23903 25248
rect 23845 25239 23903 25245
rect 23934 25236 23940 25248
rect 23992 25236 23998 25288
rect 24044 25276 24072 25304
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 24044 25248 24685 25276
rect 24673 25245 24685 25248
rect 24719 25245 24731 25279
rect 24673 25239 24731 25245
rect 7098 25168 7104 25220
rect 7156 25208 7162 25220
rect 7156 25180 7590 25208
rect 7156 25168 7162 25180
rect 8386 25168 8392 25220
rect 8444 25208 8450 25220
rect 10413 25211 10471 25217
rect 10413 25208 10425 25211
rect 8444 25180 10425 25208
rect 8444 25168 8450 25180
rect 10413 25177 10425 25180
rect 10459 25177 10471 25211
rect 10413 25171 10471 25177
rect 12526 25168 12532 25220
rect 12584 25208 12590 25220
rect 13081 25211 13139 25217
rect 13081 25208 13093 25211
rect 12584 25180 13093 25208
rect 12584 25168 12590 25180
rect 13081 25177 13093 25180
rect 13127 25177 13139 25211
rect 13081 25171 13139 25177
rect 22370 25168 22376 25220
rect 22428 25208 22434 25220
rect 22428 25180 23428 25208
rect 22428 25168 22434 25180
rect 3970 25100 3976 25152
rect 4028 25140 4034 25152
rect 4111 25143 4169 25149
rect 4111 25140 4123 25143
rect 4028 25112 4123 25140
rect 4028 25100 4034 25112
rect 4111 25109 4123 25112
rect 4157 25109 4169 25143
rect 4111 25103 4169 25109
rect 5534 25100 5540 25152
rect 5592 25140 5598 25152
rect 11057 25143 11115 25149
rect 11057 25140 11069 25143
rect 5592 25112 11069 25140
rect 5592 25100 5598 25112
rect 11057 25109 11069 25112
rect 11103 25140 11115 25143
rect 11885 25143 11943 25149
rect 11885 25140 11897 25143
rect 11103 25112 11897 25140
rect 11103 25109 11115 25112
rect 11057 25103 11115 25109
rect 11885 25109 11897 25112
rect 11931 25140 11943 25143
rect 11974 25140 11980 25152
rect 11931 25112 11980 25140
rect 11931 25109 11943 25112
rect 11885 25103 11943 25109
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 12618 25100 12624 25152
rect 12676 25100 12682 25152
rect 12802 25100 12808 25152
rect 12860 25140 12866 25152
rect 12989 25143 13047 25149
rect 12989 25140 13001 25143
rect 12860 25112 13001 25140
rect 12860 25100 12866 25112
rect 12989 25109 13001 25112
rect 13035 25109 13047 25143
rect 12989 25103 13047 25109
rect 15102 25100 15108 25152
rect 15160 25100 15166 25152
rect 15197 25143 15255 25149
rect 15197 25109 15209 25143
rect 15243 25140 15255 25143
rect 16850 25140 16856 25152
rect 15243 25112 16856 25140
rect 15243 25109 15255 25112
rect 15197 25103 15255 25109
rect 16850 25100 16856 25112
rect 16908 25100 16914 25152
rect 17034 25100 17040 25152
rect 17092 25140 17098 25152
rect 17681 25143 17739 25149
rect 17681 25140 17693 25143
rect 17092 25112 17693 25140
rect 17092 25100 17098 25112
rect 17681 25109 17693 25112
rect 17727 25140 17739 25143
rect 17862 25140 17868 25152
rect 17727 25112 17868 25140
rect 17727 25109 17739 25112
rect 17681 25103 17739 25109
rect 17862 25100 17868 25112
rect 17920 25100 17926 25152
rect 19429 25143 19487 25149
rect 19429 25109 19441 25143
rect 19475 25140 19487 25143
rect 19518 25140 19524 25152
rect 19475 25112 19524 25140
rect 19475 25109 19487 25112
rect 19429 25103 19487 25109
rect 19518 25100 19524 25112
rect 19576 25100 19582 25152
rect 22462 25100 22468 25152
rect 22520 25140 22526 25152
rect 23293 25143 23351 25149
rect 23293 25140 23305 25143
rect 22520 25112 23305 25140
rect 22520 25100 22526 25112
rect 23293 25109 23305 25112
rect 23339 25109 23351 25143
rect 23400 25140 23428 25180
rect 24026 25168 24032 25220
rect 24084 25168 24090 25220
rect 24765 25143 24823 25149
rect 24765 25140 24777 25143
rect 23400 25112 24777 25140
rect 23293 25103 23351 25109
rect 24765 25109 24777 25112
rect 24811 25109 24823 25143
rect 24765 25103 24823 25109
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 4246 24896 4252 24948
rect 4304 24936 4310 24948
rect 5445 24939 5503 24945
rect 5445 24936 5457 24939
rect 4304 24908 5457 24936
rect 4304 24896 4310 24908
rect 5445 24905 5457 24908
rect 5491 24905 5503 24939
rect 5445 24899 5503 24905
rect 7834 24896 7840 24948
rect 7892 24936 7898 24948
rect 8021 24939 8079 24945
rect 8021 24936 8033 24939
rect 7892 24908 8033 24936
rect 7892 24896 7898 24908
rect 8021 24905 8033 24908
rect 8067 24905 8079 24939
rect 8021 24899 8079 24905
rect 12618 24896 12624 24948
rect 12676 24936 12682 24948
rect 15197 24939 15255 24945
rect 15197 24936 15209 24939
rect 12676 24908 15209 24936
rect 12676 24896 12682 24908
rect 15197 24905 15209 24908
rect 15243 24905 15255 24939
rect 15197 24899 15255 24905
rect 16850 24896 16856 24948
rect 16908 24896 16914 24948
rect 17221 24939 17279 24945
rect 17221 24905 17233 24939
rect 17267 24936 17279 24939
rect 17770 24936 17776 24948
rect 17267 24908 17776 24936
rect 17267 24905 17279 24908
rect 17221 24899 17279 24905
rect 7098 24828 7104 24880
rect 7156 24828 7162 24880
rect 7466 24828 7472 24880
rect 7524 24868 7530 24880
rect 9217 24871 9275 24877
rect 7524 24840 8340 24868
rect 7524 24828 7530 24840
rect 4982 24760 4988 24812
rect 5040 24800 5046 24812
rect 5721 24803 5779 24809
rect 5721 24800 5733 24803
rect 5040 24772 5733 24800
rect 5040 24760 5046 24772
rect 5721 24769 5733 24772
rect 5767 24800 5779 24803
rect 7116 24800 7144 24828
rect 5767 24772 7144 24800
rect 5767 24769 5779 24772
rect 5721 24763 5779 24769
rect 7374 24760 7380 24812
rect 7432 24760 7438 24812
rect 7742 24760 7748 24812
rect 7800 24800 7806 24812
rect 8312 24800 8340 24840
rect 9217 24837 9229 24871
rect 9263 24868 9275 24871
rect 12069 24871 12127 24877
rect 9263 24840 10088 24868
rect 9263 24837 9275 24840
rect 9217 24831 9275 24837
rect 10060 24809 10088 24840
rect 12069 24837 12081 24871
rect 12115 24868 12127 24871
rect 13354 24868 13360 24880
rect 12115 24840 13360 24868
rect 12115 24837 12127 24840
rect 12069 24831 12127 24837
rect 13354 24828 13360 24840
rect 13412 24828 13418 24880
rect 10045 24803 10103 24809
rect 7800 24772 8248 24800
rect 8312 24772 9444 24800
rect 7800 24760 7806 24772
rect 3697 24735 3755 24741
rect 3697 24701 3709 24735
rect 3743 24701 3755 24735
rect 3697 24695 3755 24701
rect 3973 24735 4031 24741
rect 3973 24701 3985 24735
rect 4019 24732 4031 24735
rect 5994 24732 6000 24744
rect 4019 24704 6000 24732
rect 4019 24701 4031 24704
rect 3973 24695 4031 24701
rect 3712 24596 3740 24695
rect 5994 24692 6000 24704
rect 6052 24692 6058 24744
rect 7392 24732 7420 24760
rect 8110 24732 8116 24744
rect 7392 24704 8116 24732
rect 8110 24692 8116 24704
rect 8168 24692 8174 24744
rect 8220 24741 8248 24772
rect 8205 24735 8263 24741
rect 8205 24701 8217 24735
rect 8251 24701 8263 24735
rect 8205 24695 8263 24701
rect 9306 24692 9312 24744
rect 9364 24692 9370 24744
rect 9416 24741 9444 24772
rect 10045 24769 10057 24803
rect 10091 24769 10103 24803
rect 10045 24763 10103 24769
rect 12161 24803 12219 24809
rect 12161 24769 12173 24803
rect 12207 24800 12219 24803
rect 13630 24800 13636 24812
rect 12207 24772 12434 24800
rect 12207 24769 12219 24772
rect 12161 24763 12219 24769
rect 9401 24735 9459 24741
rect 9401 24701 9413 24735
rect 9447 24701 9459 24735
rect 9401 24695 9459 24701
rect 9674 24692 9680 24744
rect 9732 24732 9738 24744
rect 12253 24735 12311 24741
rect 12253 24732 12265 24735
rect 9732 24704 12265 24732
rect 9732 24692 9738 24704
rect 12253 24701 12265 24704
rect 12299 24701 12311 24735
rect 12406 24732 12434 24772
rect 12820 24772 13636 24800
rect 12820 24732 12848 24772
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 13814 24760 13820 24812
rect 13872 24760 13878 24812
rect 15010 24760 15016 24812
rect 15068 24800 15074 24812
rect 15289 24803 15347 24809
rect 15289 24800 15301 24803
rect 15068 24772 15301 24800
rect 15068 24760 15074 24772
rect 15289 24769 15301 24772
rect 15335 24769 15347 24803
rect 15289 24763 15347 24769
rect 16485 24803 16543 24809
rect 16485 24769 16497 24803
rect 16531 24800 16543 24803
rect 16850 24800 16856 24812
rect 16531 24772 16856 24800
rect 16531 24769 16543 24772
rect 16485 24763 16543 24769
rect 16850 24760 16856 24772
rect 16908 24800 16914 24812
rect 17236 24800 17264 24899
rect 17770 24896 17776 24908
rect 17828 24896 17834 24948
rect 18322 24896 18328 24948
rect 18380 24936 18386 24948
rect 18417 24939 18475 24945
rect 18417 24936 18429 24939
rect 18380 24908 18429 24936
rect 18380 24896 18386 24908
rect 18417 24905 18429 24908
rect 18463 24905 18475 24939
rect 18417 24899 18475 24905
rect 19334 24896 19340 24948
rect 19392 24936 19398 24948
rect 19610 24936 19616 24948
rect 19392 24908 19616 24936
rect 19392 24896 19398 24908
rect 19610 24896 19616 24908
rect 19668 24936 19674 24948
rect 19889 24939 19947 24945
rect 19889 24936 19901 24939
rect 19668 24908 19901 24936
rect 19668 24896 19674 24908
rect 19889 24905 19901 24908
rect 19935 24936 19947 24939
rect 20625 24939 20683 24945
rect 20625 24936 20637 24939
rect 19935 24908 20637 24936
rect 19935 24905 19947 24908
rect 19889 24899 19947 24905
rect 20625 24905 20637 24908
rect 20671 24905 20683 24939
rect 20625 24899 20683 24905
rect 20548 24840 20760 24868
rect 16908 24772 17264 24800
rect 16908 24760 16914 24772
rect 18414 24760 18420 24812
rect 18472 24800 18478 24812
rect 18509 24803 18567 24809
rect 18509 24800 18521 24803
rect 18472 24772 18521 24800
rect 18472 24760 18478 24772
rect 18509 24769 18521 24772
rect 18555 24800 18567 24803
rect 20548 24800 20576 24840
rect 18555 24772 20576 24800
rect 20732 24800 20760 24840
rect 22646 24828 22652 24880
rect 22704 24868 22710 24880
rect 23201 24871 23259 24877
rect 23201 24868 23213 24871
rect 22704 24840 23213 24868
rect 22704 24828 22710 24840
rect 23201 24837 23213 24840
rect 23247 24837 23259 24871
rect 24946 24868 24952 24880
rect 23201 24831 23259 24837
rect 24872 24840 24952 24868
rect 20732 24772 20944 24800
rect 18555 24769 18567 24772
rect 18509 24763 18567 24769
rect 13909 24735 13967 24741
rect 13909 24732 13921 24735
rect 12406 24704 12848 24732
rect 13096 24704 13921 24732
rect 12253 24695 12311 24701
rect 7653 24667 7711 24673
rect 7653 24633 7665 24667
rect 7699 24664 7711 24667
rect 8386 24664 8392 24676
rect 7699 24636 8392 24664
rect 7699 24633 7711 24636
rect 7653 24627 7711 24633
rect 8386 24624 8392 24636
rect 8444 24624 8450 24676
rect 11701 24667 11759 24673
rect 11701 24664 11713 24667
rect 8496 24636 11713 24664
rect 3970 24596 3976 24608
rect 3712 24568 3976 24596
rect 3970 24556 3976 24568
rect 4028 24556 4034 24608
rect 7466 24556 7472 24608
rect 7524 24596 7530 24608
rect 8496 24596 8524 24636
rect 11701 24633 11713 24636
rect 11747 24633 11759 24667
rect 11701 24627 11759 24633
rect 12452 24608 12480 24704
rect 12526 24624 12532 24676
rect 12584 24664 12590 24676
rect 13096 24673 13124 24704
rect 13909 24701 13921 24704
rect 13955 24701 13967 24735
rect 13909 24695 13967 24701
rect 14090 24692 14096 24744
rect 14148 24692 14154 24744
rect 14366 24692 14372 24744
rect 14424 24732 14430 24744
rect 15381 24735 15439 24741
rect 15381 24732 15393 24735
rect 14424 24704 15393 24732
rect 14424 24692 14430 24704
rect 15381 24701 15393 24704
rect 15427 24701 15439 24735
rect 15381 24695 15439 24701
rect 16574 24692 16580 24744
rect 16632 24732 16638 24744
rect 17313 24735 17371 24741
rect 17313 24732 17325 24735
rect 16632 24704 17325 24732
rect 16632 24692 16638 24704
rect 17313 24701 17325 24704
rect 17359 24701 17371 24735
rect 17313 24695 17371 24701
rect 17494 24692 17500 24744
rect 17552 24692 17558 24744
rect 18598 24692 18604 24744
rect 18656 24692 18662 24744
rect 18690 24692 18696 24744
rect 18748 24732 18754 24744
rect 20714 24732 20720 24744
rect 18748 24704 20720 24732
rect 18748 24692 18754 24704
rect 20714 24692 20720 24704
rect 20772 24692 20778 24744
rect 20809 24735 20867 24741
rect 20809 24701 20821 24735
rect 20855 24701 20867 24735
rect 20916 24732 20944 24772
rect 22002 24760 22008 24812
rect 22060 24800 22066 24812
rect 22094 24800 22100 24812
rect 22060 24772 22100 24800
rect 22060 24760 22066 24772
rect 22094 24760 22100 24772
rect 22152 24800 22158 24812
rect 22152 24772 22968 24800
rect 22152 24760 22158 24772
rect 22940 24741 22968 24772
rect 24302 24760 24308 24812
rect 24360 24800 24366 24812
rect 24872 24800 24900 24840
rect 24946 24828 24952 24840
rect 25004 24828 25010 24880
rect 24360 24772 24900 24800
rect 25317 24803 25375 24809
rect 24360 24760 24366 24772
rect 25317 24769 25329 24803
rect 25363 24800 25375 24803
rect 25498 24800 25504 24812
rect 25363 24772 25504 24800
rect 25363 24769 25375 24772
rect 25317 24763 25375 24769
rect 25498 24760 25504 24772
rect 25556 24760 25562 24812
rect 22925 24735 22983 24741
rect 20916 24704 22876 24732
rect 20809 24695 20867 24701
rect 13081 24667 13139 24673
rect 13081 24664 13093 24667
rect 12584 24636 13093 24664
rect 12584 24624 12590 24636
rect 13081 24633 13093 24636
rect 13127 24633 13139 24667
rect 13081 24627 13139 24633
rect 13449 24667 13507 24673
rect 13449 24633 13461 24667
rect 13495 24664 13507 24667
rect 15102 24664 15108 24676
rect 13495 24636 15108 24664
rect 13495 24633 13507 24636
rect 13449 24627 13507 24633
rect 15102 24624 15108 24636
rect 15160 24624 15166 24676
rect 17678 24664 17684 24676
rect 16316 24636 17684 24664
rect 7524 24568 8524 24596
rect 8849 24599 8907 24605
rect 7524 24556 7530 24568
rect 8849 24565 8861 24599
rect 8895 24596 8907 24599
rect 11146 24596 11152 24608
rect 8895 24568 11152 24596
rect 8895 24565 8907 24568
rect 8849 24559 8907 24565
rect 11146 24556 11152 24568
rect 11204 24556 11210 24608
rect 12434 24556 12440 24608
rect 12492 24556 12498 24608
rect 12618 24556 12624 24608
rect 12676 24596 12682 24608
rect 12713 24599 12771 24605
rect 12713 24596 12725 24599
rect 12676 24568 12725 24596
rect 12676 24556 12682 24568
rect 12713 24565 12725 24568
rect 12759 24565 12771 24599
rect 12713 24559 12771 24565
rect 12989 24599 13047 24605
rect 12989 24565 13001 24599
rect 13035 24596 13047 24599
rect 13354 24596 13360 24608
rect 13035 24568 13360 24596
rect 13035 24565 13047 24568
rect 12989 24559 13047 24565
rect 13354 24556 13360 24568
rect 13412 24556 13418 24608
rect 14829 24599 14887 24605
rect 14829 24565 14841 24599
rect 14875 24596 14887 24599
rect 16316 24596 16344 24636
rect 17678 24624 17684 24636
rect 17736 24624 17742 24676
rect 20162 24624 20168 24676
rect 20220 24664 20226 24676
rect 20622 24664 20628 24676
rect 20220 24636 20628 24664
rect 20220 24624 20226 24636
rect 20622 24624 20628 24636
rect 20680 24664 20686 24676
rect 20824 24664 20852 24695
rect 22646 24664 22652 24676
rect 20680 24636 20852 24664
rect 22066 24636 22652 24664
rect 20680 24624 20686 24636
rect 14875 24568 16344 24596
rect 18049 24599 18107 24605
rect 14875 24565 14887 24568
rect 14829 24559 14887 24565
rect 18049 24565 18061 24599
rect 18095 24596 18107 24599
rect 18506 24596 18512 24608
rect 18095 24568 18512 24596
rect 18095 24565 18107 24568
rect 18049 24559 18107 24565
rect 18506 24556 18512 24568
rect 18564 24556 18570 24608
rect 20257 24599 20315 24605
rect 20257 24565 20269 24599
rect 20303 24596 20315 24599
rect 22066 24596 22094 24636
rect 22646 24624 22652 24636
rect 22704 24624 22710 24676
rect 20303 24568 22094 24596
rect 22848 24596 22876 24704
rect 22925 24701 22937 24735
rect 22971 24701 22983 24735
rect 22925 24695 22983 24701
rect 24670 24692 24676 24744
rect 24728 24692 24734 24744
rect 25133 24667 25191 24673
rect 25133 24633 25145 24667
rect 25179 24633 25191 24667
rect 25133 24627 25191 24633
rect 25148 24596 25176 24627
rect 22848 24568 25176 24596
rect 20303 24565 20315 24568
rect 20257 24559 20315 24565
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 3237 24395 3295 24401
rect 3237 24361 3249 24395
rect 3283 24361 3295 24395
rect 3237 24355 3295 24361
rect 3252 24324 3280 24355
rect 3326 24352 3332 24404
rect 3384 24392 3390 24404
rect 3421 24395 3479 24401
rect 3421 24392 3433 24395
rect 3384 24364 3433 24392
rect 3384 24352 3390 24364
rect 3421 24361 3433 24364
rect 3467 24361 3479 24395
rect 4430 24392 4436 24404
rect 3421 24355 3479 24361
rect 3528 24364 4436 24392
rect 3528 24324 3556 24364
rect 4430 24352 4436 24364
rect 4488 24392 4494 24404
rect 5721 24395 5779 24401
rect 5721 24392 5733 24395
rect 4488 24364 5733 24392
rect 4488 24352 4494 24364
rect 5721 24361 5733 24364
rect 5767 24361 5779 24395
rect 5721 24355 5779 24361
rect 6178 24352 6184 24404
rect 6236 24352 6242 24404
rect 8662 24352 8668 24404
rect 8720 24392 8726 24404
rect 8757 24395 8815 24401
rect 8757 24392 8769 24395
rect 8720 24364 8769 24392
rect 8720 24352 8726 24364
rect 8757 24361 8769 24364
rect 8803 24392 8815 24395
rect 9306 24392 9312 24404
rect 8803 24364 9312 24392
rect 8803 24361 8815 24364
rect 8757 24355 8815 24361
rect 9306 24352 9312 24364
rect 9364 24352 9370 24404
rect 9968 24364 12434 24392
rect 3252 24296 3556 24324
rect 6086 24284 6092 24336
rect 6144 24324 6150 24336
rect 6144 24296 8524 24324
rect 6144 24284 6150 24296
rect 4246 24216 4252 24268
rect 4304 24216 4310 24268
rect 4982 24216 4988 24268
rect 5040 24256 5046 24268
rect 6641 24259 6699 24265
rect 6641 24256 6653 24259
rect 5040 24228 6653 24256
rect 5040 24216 5046 24228
rect 6641 24225 6653 24228
rect 6687 24256 6699 24259
rect 8294 24256 8300 24268
rect 6687 24228 8300 24256
rect 6687 24225 6699 24228
rect 6641 24219 6699 24225
rect 8294 24216 8300 24228
rect 8352 24216 8358 24268
rect 8496 24256 8524 24296
rect 9968 24256 9996 24364
rect 12406 24324 12434 24364
rect 13630 24352 13636 24404
rect 13688 24392 13694 24404
rect 13725 24395 13783 24401
rect 13725 24392 13737 24395
rect 13688 24364 13737 24392
rect 13688 24352 13694 24364
rect 13725 24361 13737 24364
rect 13771 24392 13783 24395
rect 15470 24392 15476 24404
rect 13771 24364 15476 24392
rect 13771 24361 13783 24364
rect 13725 24355 13783 24361
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 16850 24352 16856 24404
rect 16908 24352 16914 24404
rect 16868 24324 16896 24352
rect 10152 24296 11376 24324
rect 12406 24296 16896 24324
rect 8496 24228 9996 24256
rect 10042 24216 10048 24268
rect 10100 24216 10106 24268
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2774 24188 2780 24200
rect 2271 24160 2780 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2774 24148 2780 24160
rect 2832 24148 2838 24200
rect 2961 24191 3019 24197
rect 2961 24157 2973 24191
rect 3007 24188 3019 24191
rect 3510 24188 3516 24200
rect 3007 24160 3516 24188
rect 3007 24157 3019 24160
rect 2961 24151 3019 24157
rect 2685 24123 2743 24129
rect 2685 24089 2697 24123
rect 2731 24120 2743 24123
rect 2976 24120 3004 24151
rect 3510 24148 3516 24160
rect 3568 24148 3574 24200
rect 3970 24148 3976 24200
rect 4028 24148 4034 24200
rect 6365 24191 6423 24197
rect 6365 24157 6377 24191
rect 6411 24188 6423 24191
rect 7006 24188 7012 24200
rect 6411 24160 7012 24188
rect 6411 24157 6423 24160
rect 6365 24151 6423 24157
rect 7006 24148 7012 24160
rect 7064 24148 7070 24200
rect 8570 24148 8576 24200
rect 8628 24188 8634 24200
rect 10152 24188 10180 24296
rect 11238 24216 11244 24268
rect 11296 24216 11302 24268
rect 11348 24265 11376 24296
rect 24670 24284 24676 24336
rect 24728 24324 24734 24336
rect 24728 24296 25176 24324
rect 24728 24284 24734 24296
rect 11333 24259 11391 24265
rect 11333 24225 11345 24259
rect 11379 24225 11391 24259
rect 12529 24259 12587 24265
rect 12529 24256 12541 24259
rect 11333 24219 11391 24225
rect 12406 24228 12541 24256
rect 8628 24160 10180 24188
rect 8628 24148 8634 24160
rect 11146 24148 11152 24200
rect 11204 24148 11210 24200
rect 12406 24188 12434 24228
rect 12529 24225 12541 24228
rect 12575 24225 12587 24259
rect 12529 24219 12587 24225
rect 12802 24216 12808 24268
rect 12860 24256 12866 24268
rect 13173 24259 13231 24265
rect 13173 24256 13185 24259
rect 12860 24228 13185 24256
rect 12860 24216 12866 24228
rect 13173 24225 13185 24228
rect 13219 24225 13231 24259
rect 13173 24219 13231 24225
rect 13814 24216 13820 24268
rect 13872 24256 13878 24268
rect 14277 24259 14335 24265
rect 14277 24256 14289 24259
rect 13872 24228 14289 24256
rect 13872 24216 13878 24228
rect 14277 24225 14289 24228
rect 14323 24225 14335 24259
rect 14277 24219 14335 24225
rect 16853 24259 16911 24265
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 16942 24256 16948 24268
rect 16899 24228 16948 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 17034 24216 17040 24268
rect 17092 24216 17098 24268
rect 19705 24259 19763 24265
rect 19705 24225 19717 24259
rect 19751 24256 19763 24259
rect 22094 24256 22100 24268
rect 19751 24228 22100 24256
rect 19751 24225 19763 24228
rect 19705 24219 19763 24225
rect 22094 24216 22100 24228
rect 22152 24216 22158 24268
rect 23845 24259 23903 24265
rect 23845 24225 23857 24259
rect 23891 24256 23903 24259
rect 24946 24256 24952 24268
rect 23891 24228 24952 24256
rect 23891 24225 23903 24228
rect 23845 24219 23903 24225
rect 24946 24216 24952 24228
rect 25004 24216 25010 24268
rect 25148 24265 25176 24296
rect 25133 24259 25191 24265
rect 25133 24225 25145 24259
rect 25179 24225 25191 24259
rect 25133 24219 25191 24225
rect 11256 24160 12434 24188
rect 2731 24092 3004 24120
rect 3528 24120 3556 24148
rect 4522 24120 4528 24132
rect 3528 24092 4528 24120
rect 2731 24089 2743 24092
rect 2685 24083 2743 24089
rect 4522 24080 4528 24092
rect 4580 24080 4586 24132
rect 4982 24080 4988 24132
rect 5040 24080 5046 24132
rect 10962 24080 10968 24132
rect 11020 24120 11026 24132
rect 11256 24120 11284 24160
rect 16758 24148 16764 24200
rect 16816 24148 16822 24200
rect 17310 24148 17316 24200
rect 17368 24188 17374 24200
rect 17773 24191 17831 24197
rect 17773 24188 17785 24191
rect 17368 24160 17785 24188
rect 17368 24148 17374 24160
rect 17773 24157 17785 24160
rect 17819 24157 17831 24191
rect 17773 24151 17831 24157
rect 20990 24148 20996 24200
rect 21048 24188 21054 24200
rect 21450 24188 21456 24200
rect 21048 24160 21456 24188
rect 21048 24148 21054 24160
rect 21450 24148 21456 24160
rect 21508 24148 21514 24200
rect 21542 24148 21548 24200
rect 21600 24188 21606 24200
rect 22833 24191 22891 24197
rect 21600 24160 22600 24188
rect 21600 24148 21606 24160
rect 11020 24092 11284 24120
rect 11020 24080 11026 24092
rect 11514 24080 11520 24132
rect 11572 24120 11578 24132
rect 12158 24120 12164 24132
rect 11572 24092 12164 24120
rect 11572 24080 11578 24092
rect 12158 24080 12164 24092
rect 12216 24120 12222 24132
rect 12437 24123 12495 24129
rect 12437 24120 12449 24123
rect 12216 24092 12449 24120
rect 12216 24080 12222 24092
rect 12437 24089 12449 24092
rect 12483 24089 12495 24123
rect 12437 24083 12495 24089
rect 14090 24080 14096 24132
rect 14148 24120 14154 24132
rect 17494 24120 17500 24132
rect 14148 24092 17500 24120
rect 14148 24080 14154 24092
rect 17494 24080 17500 24092
rect 17552 24080 17558 24132
rect 18414 24080 18420 24132
rect 18472 24120 18478 24132
rect 18598 24120 18604 24132
rect 18472 24092 18604 24120
rect 18472 24080 18478 24092
rect 18598 24080 18604 24092
rect 18656 24120 18662 24132
rect 19886 24120 19892 24132
rect 18656 24092 19892 24120
rect 18656 24080 18662 24092
rect 19886 24080 19892 24092
rect 19944 24120 19950 24132
rect 19981 24123 20039 24129
rect 19981 24120 19993 24123
rect 19944 24092 19993 24120
rect 19944 24080 19950 24092
rect 19981 24089 19993 24092
rect 20027 24089 20039 24123
rect 19981 24083 20039 24089
rect 21818 24080 21824 24132
rect 21876 24120 21882 24132
rect 21969 24123 22027 24129
rect 21969 24120 21981 24123
rect 21876 24092 21981 24120
rect 21876 24080 21882 24092
rect 21969 24089 21981 24092
rect 22015 24089 22027 24123
rect 21969 24083 22027 24089
rect 22186 24080 22192 24132
rect 22244 24080 22250 24132
rect 22572 24120 22600 24160
rect 22833 24157 22845 24191
rect 22879 24188 22891 24191
rect 23474 24188 23480 24200
rect 22879 24160 23480 24188
rect 22879 24157 22891 24160
rect 22833 24151 22891 24157
rect 23474 24148 23480 24160
rect 23532 24148 23538 24200
rect 25041 24123 25099 24129
rect 25041 24120 25053 24123
rect 22572 24092 25053 24120
rect 25041 24089 25053 24092
rect 25087 24089 25099 24123
rect 25041 24083 25099 24089
rect 1854 24012 1860 24064
rect 1912 24052 1918 24064
rect 2041 24055 2099 24061
rect 2041 24052 2053 24055
rect 1912 24024 2053 24052
rect 1912 24012 1918 24024
rect 2041 24021 2053 24024
rect 2087 24021 2099 24055
rect 2041 24015 2099 24021
rect 8754 24012 8760 24064
rect 8812 24052 8818 24064
rect 9401 24055 9459 24061
rect 9401 24052 9413 24055
rect 8812 24024 9413 24052
rect 8812 24012 8818 24024
rect 9401 24021 9413 24024
rect 9447 24021 9459 24055
rect 9401 24015 9459 24021
rect 9766 24012 9772 24064
rect 9824 24012 9830 24064
rect 9861 24055 9919 24061
rect 9861 24021 9873 24055
rect 9907 24052 9919 24055
rect 10502 24052 10508 24064
rect 9907 24024 10508 24052
rect 9907 24021 9919 24024
rect 9861 24015 9919 24021
rect 10502 24012 10508 24024
rect 10560 24012 10566 24064
rect 10781 24055 10839 24061
rect 10781 24021 10793 24055
rect 10827 24052 10839 24055
rect 11146 24052 11152 24064
rect 10827 24024 11152 24052
rect 10827 24021 10839 24024
rect 10781 24015 10839 24021
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 11974 24012 11980 24064
rect 12032 24012 12038 24064
rect 12345 24055 12403 24061
rect 12345 24021 12357 24055
rect 12391 24052 12403 24055
rect 13630 24052 13636 24064
rect 12391 24024 13636 24052
rect 12391 24021 12403 24024
rect 12345 24015 12403 24021
rect 13630 24012 13636 24024
rect 13688 24012 13694 24064
rect 16393 24055 16451 24061
rect 16393 24021 16405 24055
rect 16439 24052 16451 24055
rect 16666 24052 16672 24064
rect 16439 24024 16672 24052
rect 16439 24021 16451 24024
rect 16393 24015 16451 24021
rect 16666 24012 16672 24024
rect 16724 24012 16730 24064
rect 17589 24055 17647 24061
rect 17589 24021 17601 24055
rect 17635 24052 17647 24055
rect 17862 24052 17868 24064
rect 17635 24024 17868 24052
rect 17635 24021 17647 24024
rect 17589 24015 17647 24021
rect 17862 24012 17868 24024
rect 17920 24012 17926 24064
rect 20254 24012 20260 24064
rect 20312 24052 20318 24064
rect 21453 24055 21511 24061
rect 21453 24052 21465 24055
rect 20312 24024 21465 24052
rect 20312 24012 20318 24024
rect 21453 24021 21465 24024
rect 21499 24021 21511 24055
rect 21453 24015 21511 24021
rect 22462 24012 22468 24064
rect 22520 24052 22526 24064
rect 24581 24055 24639 24061
rect 24581 24052 24593 24055
rect 22520 24024 24593 24052
rect 22520 24012 22526 24024
rect 24581 24021 24593 24024
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 24854 24012 24860 24064
rect 24912 24052 24918 24064
rect 24949 24055 25007 24061
rect 24949 24052 24961 24055
rect 24912 24024 24961 24052
rect 24912 24012 24918 24024
rect 24949 24021 24961 24024
rect 24995 24021 25007 24055
rect 24949 24015 25007 24021
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 5994 23808 6000 23860
rect 6052 23808 6058 23860
rect 6822 23808 6828 23860
rect 6880 23848 6886 23860
rect 9401 23851 9459 23857
rect 9401 23848 9413 23851
rect 6880 23820 9413 23848
rect 6880 23808 6886 23820
rect 9401 23817 9413 23820
rect 9447 23848 9459 23851
rect 9674 23848 9680 23860
rect 9447 23820 9680 23848
rect 9447 23817 9459 23820
rect 9401 23811 9459 23817
rect 9674 23808 9680 23820
rect 9732 23808 9738 23860
rect 9766 23808 9772 23860
rect 9824 23848 9830 23860
rect 9861 23851 9919 23857
rect 9861 23848 9873 23851
rect 9824 23820 9873 23848
rect 9824 23808 9830 23820
rect 9861 23817 9873 23820
rect 9907 23817 9919 23851
rect 9861 23811 9919 23817
rect 10502 23808 10508 23860
rect 10560 23848 10566 23860
rect 11238 23848 11244 23860
rect 10560 23820 11244 23848
rect 10560 23808 10566 23820
rect 11238 23808 11244 23820
rect 11296 23808 11302 23860
rect 11514 23808 11520 23860
rect 11572 23848 11578 23860
rect 11793 23851 11851 23857
rect 11793 23848 11805 23851
rect 11572 23820 11805 23848
rect 11572 23808 11578 23820
rect 11793 23817 11805 23820
rect 11839 23817 11851 23851
rect 11793 23811 11851 23817
rect 12434 23808 12440 23860
rect 12492 23848 12498 23860
rect 12529 23851 12587 23857
rect 12529 23848 12541 23851
rect 12492 23820 12541 23848
rect 12492 23808 12498 23820
rect 12529 23817 12541 23820
rect 12575 23848 12587 23851
rect 12802 23848 12808 23860
rect 12575 23820 12808 23848
rect 12575 23817 12587 23820
rect 12529 23811 12587 23817
rect 12802 23808 12808 23820
rect 12860 23808 12866 23860
rect 17494 23808 17500 23860
rect 17552 23848 17558 23860
rect 17552 23820 20392 23848
rect 17552 23808 17558 23820
rect 6365 23783 6423 23789
rect 6365 23780 6377 23783
rect 5750 23752 6377 23780
rect 6365 23749 6377 23752
rect 6411 23780 6423 23783
rect 7098 23780 7104 23792
rect 6411 23752 7104 23780
rect 6411 23749 6423 23752
rect 6365 23743 6423 23749
rect 7098 23740 7104 23752
rect 7156 23740 7162 23792
rect 8202 23740 8208 23792
rect 8260 23780 8266 23792
rect 11256 23780 11284 23808
rect 11882 23780 11888 23792
rect 8260 23752 8418 23780
rect 11256 23752 11888 23780
rect 8260 23740 8266 23752
rect 11882 23740 11888 23752
rect 11940 23740 11946 23792
rect 13906 23740 13912 23792
rect 13964 23780 13970 23792
rect 17954 23780 17960 23792
rect 13964 23752 17960 23780
rect 13964 23740 13970 23752
rect 17954 23740 17960 23752
rect 18012 23740 18018 23792
rect 1762 23672 1768 23724
rect 1820 23672 1826 23724
rect 20364 23712 20392 23820
rect 20714 23808 20720 23860
rect 20772 23848 20778 23860
rect 25133 23851 25191 23857
rect 25133 23848 25145 23851
rect 20772 23820 25145 23848
rect 20772 23808 20778 23820
rect 25133 23817 25145 23820
rect 25179 23817 25191 23851
rect 25133 23811 25191 23817
rect 20622 23740 20628 23792
rect 20680 23780 20686 23792
rect 23474 23780 23480 23792
rect 20680 23752 23480 23780
rect 20680 23740 20686 23752
rect 23474 23740 23480 23752
rect 23532 23740 23538 23792
rect 20809 23715 20867 23721
rect 20809 23712 20821 23715
rect 1302 23604 1308 23656
rect 1360 23644 1366 23656
rect 2041 23647 2099 23653
rect 2041 23644 2053 23647
rect 1360 23616 2053 23644
rect 1360 23604 1366 23616
rect 2041 23613 2053 23616
rect 2087 23613 2099 23647
rect 2041 23607 2099 23613
rect 3970 23604 3976 23656
rect 4028 23644 4034 23656
rect 4249 23647 4307 23653
rect 4249 23644 4261 23647
rect 4028 23616 4261 23644
rect 4028 23604 4034 23616
rect 4249 23613 4261 23616
rect 4295 23613 4307 23647
rect 4249 23607 4307 23613
rect 4525 23647 4583 23653
rect 4525 23613 4537 23647
rect 4571 23644 4583 23647
rect 7558 23644 7564 23656
rect 4571 23616 7564 23644
rect 4571 23613 4583 23616
rect 4525 23607 4583 23613
rect 4264 23508 4292 23607
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 7650 23604 7656 23656
rect 7708 23604 7714 23656
rect 7929 23647 7987 23653
rect 7929 23613 7941 23647
rect 7975 23644 7987 23647
rect 8570 23644 8576 23656
rect 7975 23616 8576 23644
rect 7975 23613 7987 23616
rect 7929 23607 7987 23613
rect 8570 23604 8576 23616
rect 8628 23604 8634 23656
rect 10873 23647 10931 23653
rect 10873 23613 10885 23647
rect 10919 23644 10931 23647
rect 11698 23644 11704 23656
rect 10919 23616 11704 23644
rect 10919 23613 10931 23616
rect 10873 23607 10931 23613
rect 11698 23604 11704 23616
rect 11756 23604 11762 23656
rect 12066 23604 12072 23656
rect 12124 23644 12130 23656
rect 14734 23644 14740 23656
rect 12124 23616 14740 23644
rect 12124 23604 12130 23616
rect 14734 23604 14740 23616
rect 14792 23604 14798 23656
rect 17034 23604 17040 23656
rect 17092 23604 17098 23656
rect 18598 23604 18604 23656
rect 18656 23644 18662 23656
rect 18785 23647 18843 23653
rect 18785 23644 18797 23647
rect 18656 23616 18797 23644
rect 18656 23604 18662 23616
rect 18785 23613 18797 23616
rect 18831 23613 18843 23647
rect 18785 23607 18843 23613
rect 19061 23647 19119 23653
rect 19061 23613 19073 23647
rect 19107 23644 19119 23647
rect 19794 23644 19800 23656
rect 19107 23616 19800 23644
rect 19107 23613 19119 23616
rect 19061 23607 19119 23613
rect 19794 23604 19800 23616
rect 19852 23604 19858 23656
rect 20180 23644 20208 23698
rect 20364 23684 20821 23712
rect 20809 23681 20821 23684
rect 20855 23681 20867 23715
rect 20809 23675 20867 23681
rect 22002 23672 22008 23724
rect 22060 23712 22066 23724
rect 22094 23712 22100 23724
rect 22060 23684 22100 23712
rect 22060 23672 22066 23684
rect 22094 23672 22100 23684
rect 22152 23712 22158 23724
rect 22925 23715 22983 23721
rect 22925 23712 22937 23715
rect 22152 23684 22937 23712
rect 22152 23672 22158 23684
rect 22925 23681 22937 23684
rect 22971 23681 22983 23715
rect 22925 23675 22983 23681
rect 24302 23672 24308 23724
rect 24360 23672 24366 23724
rect 25314 23672 25320 23724
rect 25372 23672 25378 23724
rect 23201 23647 23259 23653
rect 20180 23616 21220 23644
rect 5718 23508 5724 23520
rect 4264 23480 5724 23508
rect 5718 23468 5724 23480
rect 5776 23468 5782 23520
rect 7668 23508 7696 23604
rect 9950 23576 9956 23588
rect 9048 23548 9956 23576
rect 9048 23508 9076 23548
rect 9950 23536 9956 23548
rect 10008 23536 10014 23588
rect 11606 23536 11612 23588
rect 11664 23576 11670 23588
rect 16482 23576 16488 23588
rect 11664 23548 16488 23576
rect 11664 23536 11670 23548
rect 16482 23536 16488 23548
rect 16540 23536 16546 23588
rect 7668 23480 9076 23508
rect 10413 23511 10471 23517
rect 10413 23477 10425 23511
rect 10459 23508 10471 23511
rect 11330 23508 11336 23520
rect 10459 23480 11336 23508
rect 10459 23477 10471 23480
rect 10413 23471 10471 23477
rect 11330 23468 11336 23480
rect 11388 23468 11394 23520
rect 12066 23468 12072 23520
rect 12124 23508 12130 23520
rect 12161 23511 12219 23517
rect 12161 23508 12173 23511
rect 12124 23480 12173 23508
rect 12124 23468 12130 23480
rect 12161 23477 12173 23480
rect 12207 23477 12219 23511
rect 12161 23471 12219 23477
rect 12434 23468 12440 23520
rect 12492 23468 12498 23520
rect 13354 23468 13360 23520
rect 13412 23508 13418 23520
rect 20162 23508 20168 23520
rect 13412 23480 20168 23508
rect 13412 23468 13418 23480
rect 20162 23468 20168 23480
rect 20220 23468 20226 23520
rect 21192 23517 21220 23616
rect 23201 23613 23213 23647
rect 23247 23644 23259 23647
rect 23566 23644 23572 23656
rect 23247 23616 23572 23644
rect 23247 23613 23259 23616
rect 23201 23607 23259 23613
rect 23566 23604 23572 23616
rect 23624 23604 23630 23656
rect 24578 23604 24584 23656
rect 24636 23644 24642 23656
rect 24673 23647 24731 23653
rect 24673 23644 24685 23647
rect 24636 23616 24685 23644
rect 24636 23604 24642 23616
rect 24673 23613 24685 23616
rect 24719 23613 24731 23647
rect 24673 23607 24731 23613
rect 21177 23511 21235 23517
rect 21177 23477 21189 23511
rect 21223 23508 21235 23511
rect 21450 23508 21456 23520
rect 21223 23480 21456 23508
rect 21223 23477 21235 23480
rect 21177 23471 21235 23477
rect 21450 23468 21456 23480
rect 21508 23508 21514 23520
rect 21545 23511 21603 23517
rect 21545 23508 21557 23511
rect 21508 23480 21557 23508
rect 21508 23468 21514 23480
rect 21545 23477 21557 23480
rect 21591 23477 21603 23511
rect 21545 23471 21603 23477
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 2038 23264 2044 23316
rect 2096 23264 2102 23316
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 3145 23307 3203 23313
rect 3145 23304 3157 23307
rect 2924 23276 3157 23304
rect 2924 23264 2930 23276
rect 3145 23273 3157 23276
rect 3191 23273 3203 23307
rect 3145 23267 3203 23273
rect 7558 23264 7564 23316
rect 7616 23264 7622 23316
rect 10870 23264 10876 23316
rect 10928 23304 10934 23316
rect 12618 23304 12624 23316
rect 10928 23276 12624 23304
rect 10928 23264 10934 23276
rect 12618 23264 12624 23276
rect 12676 23264 12682 23316
rect 14550 23264 14556 23316
rect 14608 23304 14614 23316
rect 16022 23304 16028 23316
rect 14608 23276 16028 23304
rect 14608 23264 14614 23276
rect 16022 23264 16028 23276
rect 16080 23264 16086 23316
rect 18233 23307 18291 23313
rect 18233 23273 18245 23307
rect 18279 23304 18291 23307
rect 19426 23304 19432 23316
rect 18279 23276 19432 23304
rect 18279 23273 18291 23276
rect 18233 23267 18291 23273
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 20070 23264 20076 23316
rect 20128 23304 20134 23316
rect 20438 23304 20444 23316
rect 20128 23276 20444 23304
rect 20128 23264 20134 23276
rect 20438 23264 20444 23276
rect 20496 23304 20502 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 20496 23276 21189 23304
rect 20496 23264 20502 23276
rect 21177 23273 21189 23276
rect 21223 23273 21235 23307
rect 21177 23267 21235 23273
rect 9674 23196 9680 23248
rect 9732 23236 9738 23248
rect 11333 23239 11391 23245
rect 11333 23236 11345 23239
rect 9732 23208 11345 23236
rect 9732 23196 9738 23208
rect 11333 23205 11345 23208
rect 11379 23205 11391 23239
rect 11333 23199 11391 23205
rect 12434 23196 12440 23248
rect 12492 23236 12498 23248
rect 12989 23239 13047 23245
rect 12989 23236 13001 23239
rect 12492 23208 13001 23236
rect 12492 23196 12498 23208
rect 12989 23205 13001 23208
rect 13035 23205 13047 23239
rect 12989 23199 13047 23205
rect 23658 23196 23664 23248
rect 23716 23236 23722 23248
rect 24578 23236 24584 23248
rect 23716 23208 24584 23236
rect 23716 23196 23722 23208
rect 24578 23196 24584 23208
rect 24636 23236 24642 23248
rect 24636 23208 25176 23236
rect 24636 23196 24642 23208
rect 2866 23128 2872 23180
rect 2924 23168 2930 23180
rect 2961 23171 3019 23177
rect 2961 23168 2973 23171
rect 2924 23140 2973 23168
rect 2924 23128 2930 23140
rect 2961 23137 2973 23140
rect 3007 23168 3019 23171
rect 3326 23168 3332 23180
rect 3007 23140 3332 23168
rect 3007 23137 3019 23140
rect 2961 23131 3019 23137
rect 3326 23128 3332 23140
rect 3384 23128 3390 23180
rect 5718 23128 5724 23180
rect 5776 23168 5782 23180
rect 5813 23171 5871 23177
rect 5813 23168 5825 23171
rect 5776 23140 5825 23168
rect 5776 23128 5782 23140
rect 5813 23137 5825 23140
rect 5859 23168 5871 23171
rect 6454 23168 6460 23180
rect 5859 23140 6460 23168
rect 5859 23137 5871 23140
rect 5813 23131 5871 23137
rect 6454 23128 6460 23140
rect 6512 23128 6518 23180
rect 7098 23128 7104 23180
rect 7156 23168 7162 23180
rect 7156 23140 7236 23168
rect 7156 23128 7162 23140
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23069 2283 23103
rect 2225 23063 2283 23069
rect 2777 23103 2835 23109
rect 2777 23069 2789 23103
rect 2823 23100 2835 23103
rect 2823 23072 3924 23100
rect 2823 23069 2835 23072
rect 2777 23063 2835 23069
rect 2240 23032 2268 23063
rect 3786 23032 3792 23044
rect 2240 23004 3792 23032
rect 3786 22992 3792 23004
rect 3844 22992 3850 23044
rect 3896 23032 3924 23072
rect 3970 23060 3976 23112
rect 4028 23100 4034 23112
rect 4100 23103 4158 23109
rect 4100 23100 4112 23103
rect 4028 23072 4112 23100
rect 4028 23060 4034 23072
rect 4100 23069 4112 23072
rect 4146 23069 4158 23103
rect 4100 23063 4158 23069
rect 4203 23103 4261 23109
rect 4203 23069 4215 23103
rect 4249 23100 4261 23103
rect 4338 23100 4344 23112
rect 4249 23072 4344 23100
rect 4249 23069 4261 23072
rect 4203 23063 4261 23069
rect 4338 23060 4344 23072
rect 4396 23060 4402 23112
rect 7208 23100 7236 23140
rect 11882 23128 11888 23180
rect 11940 23128 11946 23180
rect 12713 23171 12771 23177
rect 12713 23137 12725 23171
rect 12759 23168 12771 23171
rect 13538 23168 13544 23180
rect 12759 23140 13544 23168
rect 12759 23137 12771 23140
rect 12713 23131 12771 23137
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 14274 23128 14280 23180
rect 14332 23168 14338 23180
rect 15286 23168 15292 23180
rect 14332 23140 15292 23168
rect 14332 23128 14338 23140
rect 15286 23128 15292 23140
rect 15344 23168 15350 23180
rect 16485 23171 16543 23177
rect 16485 23168 16497 23171
rect 15344 23140 16497 23168
rect 15344 23128 15350 23140
rect 16485 23137 16497 23140
rect 16531 23168 16543 23171
rect 18598 23168 18604 23180
rect 16531 23140 18604 23168
rect 16531 23137 16543 23140
rect 16485 23131 16543 23137
rect 18598 23128 18604 23140
rect 18656 23168 18662 23180
rect 25148 23177 25176 23208
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 18656 23140 19441 23168
rect 18656 23128 18662 23140
rect 19429 23137 19441 23140
rect 19475 23137 19487 23171
rect 19429 23131 19487 23137
rect 22005 23171 22063 23177
rect 22005 23137 22017 23171
rect 22051 23168 22063 23171
rect 25133 23171 25191 23177
rect 22051 23140 24992 23168
rect 22051 23137 22063 23140
rect 22005 23131 22063 23137
rect 7650 23100 7656 23112
rect 7208 23086 7656 23100
rect 7222 23072 7656 23086
rect 7650 23060 7656 23072
rect 7708 23100 7714 23112
rect 7837 23103 7895 23109
rect 7837 23100 7849 23103
rect 7708 23072 7849 23100
rect 7708 23060 7714 23072
rect 7837 23069 7849 23072
rect 7883 23069 7895 23103
rect 7837 23063 7895 23069
rect 9306 23060 9312 23112
rect 9364 23100 9370 23112
rect 9953 23103 10011 23109
rect 9953 23100 9965 23103
rect 9364 23072 9965 23100
rect 9364 23060 9370 23072
rect 9953 23069 9965 23072
rect 9999 23100 10011 23103
rect 11606 23100 11612 23112
rect 9999 23072 11612 23100
rect 9999 23069 10011 23072
rect 9953 23063 10011 23069
rect 11606 23060 11612 23072
rect 11664 23060 11670 23112
rect 11698 23060 11704 23112
rect 11756 23060 11762 23112
rect 13357 23103 13415 23109
rect 13357 23069 13369 23103
rect 13403 23100 13415 23103
rect 13906 23100 13912 23112
rect 13403 23072 13912 23100
rect 13403 23069 13415 23072
rect 13357 23063 13415 23069
rect 13906 23060 13912 23072
rect 13964 23060 13970 23112
rect 16390 23100 16396 23112
rect 15686 23072 16396 23100
rect 16390 23060 16396 23072
rect 16448 23060 16454 23112
rect 22833 23103 22891 23109
rect 22833 23069 22845 23103
rect 22879 23100 22891 23103
rect 23290 23100 23296 23112
rect 22879 23072 23296 23100
rect 22879 23069 22891 23072
rect 22833 23063 22891 23069
rect 23290 23060 23296 23072
rect 23348 23060 23354 23112
rect 23842 23060 23848 23112
rect 23900 23060 23906 23112
rect 24964 23109 24992 23140
rect 25133 23137 25145 23171
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23069 25007 23103
rect 24949 23063 25007 23069
rect 5074 23032 5080 23044
rect 3896 23004 5080 23032
rect 5074 22992 5080 23004
rect 5132 22992 5138 23044
rect 6089 23035 6147 23041
rect 6089 23001 6101 23035
rect 6135 23001 6147 23035
rect 7742 23032 7748 23044
rect 6089 22995 6147 23001
rect 7484 23004 7748 23032
rect 6104 22964 6132 22995
rect 7484 22964 7512 23004
rect 7742 22992 7748 23004
rect 7800 22992 7806 23044
rect 10689 23035 10747 23041
rect 10689 23001 10701 23035
rect 10735 23001 10747 23035
rect 10689 22995 10747 23001
rect 6104 22936 7512 22964
rect 9950 22924 9956 22976
rect 10008 22964 10014 22976
rect 10704 22964 10732 22995
rect 10778 22992 10784 23044
rect 10836 23032 10842 23044
rect 12529 23035 12587 23041
rect 12529 23032 12541 23035
rect 10836 23004 12541 23032
rect 10836 22992 10842 23004
rect 12529 23001 12541 23004
rect 12575 23032 12587 23035
rect 13449 23035 13507 23041
rect 13449 23032 13461 23035
rect 12575 23004 13461 23032
rect 12575 23001 12587 23004
rect 12529 22995 12587 23001
rect 13449 23001 13461 23004
rect 13495 23001 13507 23035
rect 13449 22995 13507 23001
rect 14553 23035 14611 23041
rect 14553 23001 14565 23035
rect 14599 23001 14611 23035
rect 14553 22995 14611 23001
rect 10008 22936 10732 22964
rect 11793 22967 11851 22973
rect 10008 22924 10014 22936
rect 11793 22933 11805 22967
rect 11839 22964 11851 22967
rect 12066 22964 12072 22976
rect 11839 22936 12072 22964
rect 11839 22933 11851 22936
rect 11793 22927 11851 22933
rect 12066 22924 12072 22936
rect 12124 22924 12130 22976
rect 14568 22964 14596 22995
rect 15930 22992 15936 23044
rect 15988 23032 15994 23044
rect 16761 23035 16819 23041
rect 16761 23032 16773 23035
rect 15988 23004 16773 23032
rect 15988 22992 15994 23004
rect 16761 23001 16773 23004
rect 16807 23001 16819 23035
rect 17986 23004 18092 23032
rect 16761 22995 16819 23001
rect 15838 22964 15844 22976
rect 14568 22936 15844 22964
rect 15838 22924 15844 22936
rect 15896 22924 15902 22976
rect 16390 22924 16396 22976
rect 16448 22964 16454 22976
rect 18064 22964 18092 23004
rect 19426 22992 19432 23044
rect 19484 23032 19490 23044
rect 19705 23035 19763 23041
rect 19705 23032 19717 23035
rect 19484 23004 19717 23032
rect 19484 22992 19490 23004
rect 19705 23001 19717 23004
rect 19751 23032 19763 23035
rect 19978 23032 19984 23044
rect 19751 23004 19984 23032
rect 19751 23001 19763 23004
rect 19705 22995 19763 23001
rect 19978 22992 19984 23004
rect 20036 22992 20042 23044
rect 20930 23004 21496 23032
rect 18601 22967 18659 22973
rect 18601 22964 18613 22967
rect 16448 22936 18613 22964
rect 16448 22924 16454 22936
rect 18601 22933 18613 22936
rect 18647 22964 18659 22967
rect 21008 22964 21036 23004
rect 21468 22976 21496 23004
rect 22646 22992 22652 23044
rect 22704 23032 22710 23044
rect 25041 23035 25099 23041
rect 25041 23032 25053 23035
rect 22704 23004 25053 23032
rect 22704 22992 22710 23004
rect 25041 23001 25053 23004
rect 25087 23001 25099 23035
rect 25041 22995 25099 23001
rect 18647 22936 21036 22964
rect 18647 22933 18659 22936
rect 18601 22927 18659 22933
rect 21450 22924 21456 22976
rect 21508 22924 21514 22976
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 23532 22936 24593 22964
rect 23532 22924 23538 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 1762 22720 1768 22772
rect 1820 22760 1826 22772
rect 2041 22763 2099 22769
rect 2041 22760 2053 22763
rect 1820 22732 2053 22760
rect 1820 22720 1826 22732
rect 2041 22729 2053 22732
rect 2087 22729 2099 22763
rect 2041 22723 2099 22729
rect 5629 22763 5687 22769
rect 5629 22729 5641 22763
rect 5675 22760 5687 22763
rect 6825 22763 6883 22769
rect 6825 22760 6837 22763
rect 5675 22732 6837 22760
rect 5675 22729 5687 22732
rect 5629 22723 5687 22729
rect 6825 22729 6837 22732
rect 6871 22729 6883 22763
rect 6825 22723 6883 22729
rect 7193 22763 7251 22769
rect 7193 22729 7205 22763
rect 7239 22760 7251 22763
rect 8754 22760 8760 22772
rect 7239 22732 8760 22760
rect 7239 22729 7251 22732
rect 7193 22723 7251 22729
rect 8754 22720 8760 22732
rect 8812 22720 8818 22772
rect 9306 22720 9312 22772
rect 9364 22720 9370 22772
rect 9858 22720 9864 22772
rect 9916 22760 9922 22772
rect 10137 22763 10195 22769
rect 10137 22760 10149 22763
rect 9916 22732 10149 22760
rect 9916 22720 9922 22732
rect 10137 22729 10149 22732
rect 10183 22760 10195 22763
rect 10870 22760 10876 22772
rect 10183 22732 10876 22760
rect 10183 22729 10195 22732
rect 10137 22723 10195 22729
rect 10870 22720 10876 22732
rect 10928 22720 10934 22772
rect 12345 22763 12403 22769
rect 12345 22729 12357 22763
rect 12391 22760 12403 22763
rect 12526 22760 12532 22772
rect 12391 22732 12532 22760
rect 12391 22729 12403 22732
rect 12345 22723 12403 22729
rect 12526 22720 12532 22732
rect 12584 22720 12590 22772
rect 14918 22720 14924 22772
rect 14976 22760 14982 22772
rect 15197 22763 15255 22769
rect 15197 22760 15209 22763
rect 14976 22732 15209 22760
rect 14976 22720 14982 22732
rect 15197 22729 15209 22732
rect 15243 22729 15255 22763
rect 15197 22723 15255 22729
rect 16209 22763 16267 22769
rect 16209 22729 16221 22763
rect 16255 22760 16267 22763
rect 16390 22760 16396 22772
rect 16255 22732 16396 22760
rect 16255 22729 16267 22732
rect 16209 22723 16267 22729
rect 16390 22720 16396 22732
rect 16448 22720 16454 22772
rect 16574 22720 16580 22772
rect 16632 22760 16638 22772
rect 17494 22760 17500 22772
rect 16632 22732 17500 22760
rect 16632 22720 16638 22732
rect 17494 22720 17500 22732
rect 17552 22760 17558 22772
rect 20346 22760 20352 22772
rect 17552 22732 20352 22760
rect 17552 22720 17558 22732
rect 8021 22695 8079 22701
rect 8021 22661 8033 22695
rect 8067 22692 8079 22695
rect 9324 22692 9352 22720
rect 8067 22664 9352 22692
rect 8067 22661 8079 22664
rect 8021 22655 8079 22661
rect 11606 22652 11612 22704
rect 11664 22692 11670 22704
rect 12158 22692 12164 22704
rect 11664 22664 12164 22692
rect 11664 22652 11670 22664
rect 12158 22652 12164 22664
rect 12216 22692 12222 22704
rect 12437 22695 12495 22701
rect 12437 22692 12449 22695
rect 12216 22664 12449 22692
rect 12216 22652 12222 22664
rect 12437 22661 12449 22664
rect 12483 22661 12495 22695
rect 12437 22655 12495 22661
rect 13081 22695 13139 22701
rect 13081 22661 13093 22695
rect 13127 22692 13139 22695
rect 15654 22692 15660 22704
rect 13127 22664 15660 22692
rect 13127 22661 13139 22664
rect 13081 22655 13139 22661
rect 2225 22627 2283 22633
rect 2225 22593 2237 22627
rect 2271 22624 2283 22627
rect 2866 22624 2872 22636
rect 2271 22596 2872 22624
rect 2271 22593 2283 22596
rect 2225 22587 2283 22593
rect 2866 22584 2872 22596
rect 2924 22584 2930 22636
rect 5721 22627 5779 22633
rect 5721 22593 5733 22627
rect 5767 22624 5779 22627
rect 6914 22624 6920 22636
rect 5767 22596 6920 22624
rect 5767 22593 5779 22596
rect 5721 22587 5779 22593
rect 6914 22584 6920 22596
rect 6972 22584 6978 22636
rect 10781 22627 10839 22633
rect 10781 22593 10793 22627
rect 10827 22624 10839 22627
rect 13096 22624 13124 22655
rect 15654 22652 15660 22664
rect 15712 22652 15718 22704
rect 17880 22701 17908 22732
rect 20346 22720 20352 22732
rect 20404 22720 20410 22772
rect 23566 22720 23572 22772
rect 23624 22760 23630 22772
rect 23753 22763 23811 22769
rect 23753 22760 23765 22763
rect 23624 22732 23765 22760
rect 23624 22720 23630 22732
rect 23753 22729 23765 22732
rect 23799 22729 23811 22763
rect 23753 22723 23811 22729
rect 24213 22763 24271 22769
rect 24213 22729 24225 22763
rect 24259 22760 24271 22763
rect 24302 22760 24308 22772
rect 24259 22732 24308 22760
rect 24259 22729 24271 22732
rect 24213 22723 24271 22729
rect 17865 22695 17923 22701
rect 17865 22661 17877 22695
rect 17911 22661 17923 22695
rect 17865 22655 17923 22661
rect 18598 22652 18604 22704
rect 18656 22652 18662 22704
rect 19702 22652 19708 22704
rect 19760 22652 19766 22704
rect 20364 22692 20392 22720
rect 20533 22695 20591 22701
rect 20533 22692 20545 22695
rect 20364 22664 20545 22692
rect 20533 22661 20545 22664
rect 20579 22661 20591 22695
rect 24228 22692 24256 22723
rect 24302 22720 24308 22732
rect 24360 22760 24366 22772
rect 24765 22763 24823 22769
rect 24765 22760 24777 22763
rect 24360 22732 24777 22760
rect 24360 22720 24366 22732
rect 24765 22729 24777 22732
rect 24811 22729 24823 22763
rect 24765 22723 24823 22729
rect 25314 22720 25320 22772
rect 25372 22760 25378 22772
rect 25409 22763 25467 22769
rect 25409 22760 25421 22763
rect 25372 22732 25421 22760
rect 25372 22720 25378 22732
rect 25409 22729 25421 22732
rect 25455 22729 25467 22763
rect 25409 22723 25467 22729
rect 23506 22664 24256 22692
rect 20533 22655 20591 22661
rect 23584 22636 23612 22664
rect 10827 22596 12296 22624
rect 10827 22593 10839 22596
rect 10781 22587 10839 22593
rect 5905 22559 5963 22565
rect 5905 22525 5917 22559
rect 5951 22556 5963 22559
rect 5994 22556 6000 22568
rect 5951 22528 6000 22556
rect 5951 22525 5963 22528
rect 5905 22519 5963 22525
rect 5994 22516 6000 22528
rect 6052 22516 6058 22568
rect 7282 22516 7288 22568
rect 7340 22516 7346 22568
rect 7469 22559 7527 22565
rect 7469 22525 7481 22559
rect 7515 22556 7527 22559
rect 7558 22556 7564 22568
rect 7515 22528 7564 22556
rect 7515 22525 7527 22528
rect 7469 22519 7527 22525
rect 7558 22516 7564 22528
rect 7616 22516 7622 22568
rect 8846 22516 8852 22568
rect 8904 22516 8910 22568
rect 10962 22516 10968 22568
rect 11020 22516 11026 22568
rect 12268 22556 12296 22596
rect 12406 22596 13124 22624
rect 12406 22556 12434 22596
rect 13814 22584 13820 22636
rect 13872 22624 13878 22636
rect 15105 22627 15163 22633
rect 15105 22624 15117 22627
rect 13872 22596 15117 22624
rect 13872 22584 13878 22596
rect 15105 22593 15117 22596
rect 15151 22593 15163 22627
rect 15105 22587 15163 22593
rect 16574 22584 16580 22636
rect 16632 22624 16638 22636
rect 16850 22624 16856 22636
rect 16632 22596 16856 22624
rect 16632 22584 16638 22596
rect 16850 22584 16856 22596
rect 16908 22584 16914 22636
rect 19610 22584 19616 22636
rect 19668 22584 19674 22636
rect 21361 22627 21419 22633
rect 21361 22593 21373 22627
rect 21407 22624 21419 22627
rect 22002 22624 22008 22636
rect 21407 22596 22008 22624
rect 21407 22593 21419 22596
rect 21361 22587 21419 22593
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 23566 22584 23572 22636
rect 23624 22584 23630 22636
rect 12268 22528 12434 22556
rect 12621 22559 12679 22565
rect 12621 22525 12633 22559
rect 12667 22556 12679 22559
rect 12667 22528 13860 22556
rect 12667 22525 12679 22528
rect 12621 22519 12679 22525
rect 9398 22448 9404 22500
rect 9456 22488 9462 22500
rect 10413 22491 10471 22497
rect 10413 22488 10425 22491
rect 9456 22460 10425 22488
rect 9456 22448 9462 22460
rect 10413 22457 10425 22460
rect 10459 22457 10471 22491
rect 10413 22451 10471 22457
rect 11977 22491 12035 22497
rect 11977 22457 11989 22491
rect 12023 22488 12035 22491
rect 13630 22488 13636 22500
rect 12023 22460 13636 22488
rect 12023 22457 12035 22460
rect 11977 22451 12035 22457
rect 13630 22448 13636 22460
rect 13688 22448 13694 22500
rect 13832 22488 13860 22528
rect 13906 22516 13912 22568
rect 13964 22516 13970 22568
rect 15381 22559 15439 22565
rect 15381 22525 15393 22559
rect 15427 22556 15439 22559
rect 15930 22556 15936 22568
rect 15427 22528 15936 22556
rect 15427 22525 15439 22528
rect 15381 22519 15439 22525
rect 15930 22516 15936 22528
rect 15988 22516 15994 22568
rect 19794 22516 19800 22568
rect 19852 22516 19858 22568
rect 21634 22516 21640 22568
rect 21692 22556 21698 22568
rect 22281 22559 22339 22565
rect 22281 22556 22293 22559
rect 21692 22528 22293 22556
rect 21692 22516 21698 22528
rect 22281 22525 22293 22528
rect 22327 22525 22339 22559
rect 22281 22519 22339 22525
rect 15838 22488 15844 22500
rect 13832 22460 15844 22488
rect 15838 22448 15844 22460
rect 15896 22448 15902 22500
rect 4246 22380 4252 22432
rect 4304 22420 4310 22432
rect 5261 22423 5319 22429
rect 5261 22420 5273 22423
rect 4304 22392 5273 22420
rect 4304 22380 4310 22392
rect 5261 22389 5273 22392
rect 5307 22389 5319 22423
rect 5261 22383 5319 22389
rect 6270 22380 6276 22432
rect 6328 22420 6334 22432
rect 11606 22420 11612 22432
rect 6328 22392 11612 22420
rect 6328 22380 6334 22392
rect 11606 22380 11612 22392
rect 11664 22380 11670 22432
rect 12526 22380 12532 22432
rect 12584 22420 12590 22432
rect 12802 22420 12808 22432
rect 12584 22392 12808 22420
rect 12584 22380 12590 22392
rect 12802 22380 12808 22392
rect 12860 22380 12866 22432
rect 14737 22423 14795 22429
rect 14737 22389 14749 22423
rect 14783 22420 14795 22423
rect 15562 22420 15568 22432
rect 14783 22392 15568 22420
rect 14783 22389 14795 22392
rect 14737 22383 14795 22389
rect 15562 22380 15568 22392
rect 15620 22380 15626 22432
rect 19242 22380 19248 22432
rect 19300 22380 19306 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 16022 22176 16028 22228
rect 16080 22216 16086 22228
rect 16390 22216 16396 22228
rect 16080 22188 16396 22216
rect 16080 22176 16086 22188
rect 16390 22176 16396 22188
rect 16448 22176 16454 22228
rect 19686 22219 19744 22225
rect 19686 22216 19698 22219
rect 18708 22188 19698 22216
rect 18414 22148 18420 22160
rect 17512 22120 18420 22148
rect 10686 22040 10692 22092
rect 10744 22080 10750 22092
rect 11885 22083 11943 22089
rect 11885 22080 11897 22083
rect 10744 22052 11897 22080
rect 10744 22040 10750 22052
rect 11885 22049 11897 22052
rect 11931 22049 11943 22083
rect 11885 22043 11943 22049
rect 12069 22083 12127 22089
rect 12069 22049 12081 22083
rect 12115 22080 12127 22083
rect 12158 22080 12164 22092
rect 12115 22052 12164 22080
rect 12115 22049 12127 22052
rect 12069 22043 12127 22049
rect 12158 22040 12164 22052
rect 12216 22040 12222 22092
rect 14274 22040 14280 22092
rect 14332 22040 14338 22092
rect 16025 22083 16083 22089
rect 16025 22049 16037 22083
rect 16071 22080 16083 22083
rect 16114 22080 16120 22092
rect 16071 22052 16120 22080
rect 16071 22049 16083 22052
rect 16025 22043 16083 22049
rect 16114 22040 16120 22052
rect 16172 22040 16178 22092
rect 17512 22089 17540 22120
rect 18414 22108 18420 22120
rect 18472 22108 18478 22160
rect 16577 22083 16635 22089
rect 16577 22049 16589 22083
rect 16623 22080 16635 22083
rect 17497 22083 17555 22089
rect 16623 22052 17356 22080
rect 16623 22049 16635 22052
rect 16577 22043 16635 22049
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 22012 11851 22015
rect 13265 22015 13323 22021
rect 11839 21984 12572 22012
rect 11839 21981 11851 21984
rect 11793 21975 11851 21981
rect 10594 21904 10600 21956
rect 10652 21944 10658 21956
rect 12544 21953 12572 21984
rect 13265 21981 13277 22015
rect 13311 22012 13323 22015
rect 13354 22012 13360 22024
rect 13311 21984 13360 22012
rect 13311 21981 13323 21984
rect 13265 21975 13323 21981
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 17034 21972 17040 22024
rect 17092 22012 17098 22024
rect 17328 22021 17356 22052
rect 17497 22049 17509 22083
rect 17543 22080 17555 22083
rect 17543 22052 17577 22080
rect 17543 22049 17555 22052
rect 17497 22043 17555 22049
rect 18506 22040 18512 22092
rect 18564 22040 18570 22092
rect 18708 22089 18736 22188
rect 19686 22185 19698 22188
rect 19732 22216 19744 22219
rect 20254 22216 20260 22228
rect 19732 22188 20260 22216
rect 19732 22185 19744 22188
rect 19686 22179 19744 22185
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 21450 22108 21456 22160
rect 21508 22108 21514 22160
rect 18693 22083 18751 22089
rect 18693 22049 18705 22083
rect 18739 22049 18751 22083
rect 22002 22080 22008 22092
rect 18693 22043 18751 22049
rect 19444 22052 22008 22080
rect 19444 22024 19472 22052
rect 22002 22040 22008 22052
rect 22060 22040 22066 22092
rect 22281 22083 22339 22089
rect 22281 22049 22293 22083
rect 22327 22080 22339 22083
rect 22646 22080 22652 22092
rect 22327 22052 22652 22080
rect 22327 22049 22339 22052
rect 22281 22043 22339 22049
rect 22646 22040 22652 22052
rect 22704 22040 22710 22092
rect 22830 22040 22836 22092
rect 22888 22080 22894 22092
rect 24029 22083 24087 22089
rect 24029 22080 24041 22083
rect 22888 22052 24041 22080
rect 22888 22040 22894 22052
rect 24029 22049 24041 22052
rect 24075 22049 24087 22083
rect 24029 22043 24087 22049
rect 17221 22015 17279 22021
rect 17221 22012 17233 22015
rect 17092 21984 17233 22012
rect 17092 21972 17098 21984
rect 17221 21981 17233 21984
rect 17267 21981 17279 22015
rect 17221 21975 17279 21981
rect 17313 22015 17371 22021
rect 17313 21981 17325 22015
rect 17359 22012 17371 22015
rect 19334 22012 19340 22024
rect 17359 21984 19340 22012
rect 17359 21981 17371 21984
rect 17313 21975 17371 21981
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 19426 21972 19432 22024
rect 19484 21972 19490 22024
rect 23566 22012 23572 22024
rect 23414 21984 23572 22012
rect 23566 21972 23572 21984
rect 23624 21972 23630 22024
rect 12529 21947 12587 21953
rect 10652 21916 11468 21944
rect 10652 21904 10658 21916
rect 4433 21879 4491 21885
rect 4433 21845 4445 21879
rect 4479 21876 4491 21879
rect 4522 21876 4528 21888
rect 4479 21848 4528 21876
rect 4479 21845 4491 21848
rect 4433 21839 4491 21845
rect 4522 21836 4528 21848
rect 4580 21836 4586 21888
rect 10686 21836 10692 21888
rect 10744 21876 10750 21888
rect 11440 21885 11468 21916
rect 12529 21913 12541 21947
rect 12575 21944 12587 21947
rect 12575 21916 14136 21944
rect 12575 21913 12587 21916
rect 12529 21907 12587 21913
rect 11057 21879 11115 21885
rect 11057 21876 11069 21879
rect 10744 21848 11069 21876
rect 10744 21836 10750 21848
rect 11057 21845 11069 21848
rect 11103 21845 11115 21879
rect 11057 21839 11115 21845
rect 11425 21879 11483 21885
rect 11425 21845 11437 21879
rect 11471 21845 11483 21879
rect 11425 21839 11483 21845
rect 13081 21879 13139 21885
rect 13081 21845 13093 21879
rect 13127 21876 13139 21879
rect 13354 21876 13360 21888
rect 13127 21848 13360 21876
rect 13127 21845 13139 21848
rect 13081 21839 13139 21845
rect 13354 21836 13360 21848
rect 13412 21836 13418 21888
rect 14108 21876 14136 21916
rect 14182 21904 14188 21956
rect 14240 21944 14246 21956
rect 14550 21944 14556 21956
rect 14240 21916 14556 21944
rect 14240 21904 14246 21916
rect 14550 21904 14556 21916
rect 14608 21904 14614 21956
rect 16022 21944 16028 21956
rect 15778 21916 16028 21944
rect 16022 21904 16028 21916
rect 16080 21904 16086 21956
rect 18417 21947 18475 21953
rect 18417 21944 18429 21947
rect 16868 21916 18429 21944
rect 15930 21876 15936 21888
rect 14108 21848 15936 21876
rect 15930 21836 15936 21848
rect 15988 21836 15994 21888
rect 16868 21885 16896 21916
rect 18417 21913 18429 21916
rect 18463 21913 18475 21947
rect 21450 21944 21456 21956
rect 20930 21916 21456 21944
rect 18417 21907 18475 21913
rect 21450 21904 21456 21916
rect 21508 21904 21514 21956
rect 24673 21947 24731 21953
rect 24673 21944 24685 21947
rect 24136 21916 24685 21944
rect 16853 21879 16911 21885
rect 16853 21845 16865 21879
rect 16899 21845 16911 21879
rect 16853 21839 16911 21845
rect 18049 21879 18107 21885
rect 18049 21845 18061 21879
rect 18095 21876 18107 21879
rect 19610 21876 19616 21888
rect 18095 21848 19616 21876
rect 18095 21845 18107 21848
rect 18049 21839 18107 21845
rect 19610 21836 19616 21848
rect 19668 21836 19674 21888
rect 19886 21836 19892 21888
rect 19944 21876 19950 21888
rect 21177 21879 21235 21885
rect 21177 21876 21189 21879
rect 19944 21848 21189 21876
rect 19944 21836 19950 21848
rect 21177 21845 21189 21848
rect 21223 21845 21235 21879
rect 21177 21839 21235 21845
rect 21726 21836 21732 21888
rect 21784 21876 21790 21888
rect 24136 21876 24164 21916
rect 24673 21913 24685 21916
rect 24719 21913 24731 21947
rect 24673 21907 24731 21913
rect 21784 21848 24164 21876
rect 21784 21836 21790 21848
rect 24210 21836 24216 21888
rect 24268 21876 24274 21888
rect 24765 21879 24823 21885
rect 24765 21876 24777 21879
rect 24268 21848 24777 21876
rect 24268 21836 24274 21848
rect 24765 21845 24777 21848
rect 24811 21845 24823 21879
rect 24765 21839 24823 21845
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 7006 21632 7012 21684
rect 7064 21672 7070 21684
rect 7101 21675 7159 21681
rect 7101 21672 7113 21675
rect 7064 21644 7113 21672
rect 7064 21632 7070 21644
rect 7101 21641 7113 21644
rect 7147 21641 7159 21675
rect 7101 21635 7159 21641
rect 7469 21675 7527 21681
rect 7469 21641 7481 21675
rect 7515 21672 7527 21675
rect 8297 21675 8355 21681
rect 8297 21672 8309 21675
rect 7515 21644 8309 21672
rect 7515 21641 7527 21644
rect 7469 21635 7527 21641
rect 8297 21641 8309 21644
rect 8343 21641 8355 21675
rect 8297 21635 8355 21641
rect 8665 21675 8723 21681
rect 8665 21641 8677 21675
rect 8711 21672 8723 21675
rect 9674 21672 9680 21684
rect 8711 21644 9680 21672
rect 8711 21641 8723 21644
rect 8665 21635 8723 21641
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 9861 21675 9919 21681
rect 9861 21641 9873 21675
rect 9907 21672 9919 21675
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 9907 21644 11713 21672
rect 9907 21641 9919 21644
rect 9861 21635 9919 21641
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 11701 21635 11759 21641
rect 11974 21632 11980 21684
rect 12032 21672 12038 21684
rect 12069 21675 12127 21681
rect 12069 21672 12081 21675
rect 12032 21644 12081 21672
rect 12032 21632 12038 21644
rect 12069 21641 12081 21644
rect 12115 21641 12127 21675
rect 12069 21635 12127 21641
rect 13541 21675 13599 21681
rect 13541 21641 13553 21675
rect 13587 21672 13599 21675
rect 13814 21672 13820 21684
rect 13587 21644 13820 21672
rect 13587 21641 13599 21644
rect 13541 21635 13599 21641
rect 13814 21632 13820 21644
rect 13872 21632 13878 21684
rect 13906 21632 13912 21684
rect 13964 21632 13970 21684
rect 16025 21675 16083 21681
rect 16025 21641 16037 21675
rect 16071 21672 16083 21675
rect 21082 21672 21088 21684
rect 16071 21644 21088 21672
rect 16071 21641 16083 21644
rect 16025 21635 16083 21641
rect 21082 21632 21088 21644
rect 21140 21632 21146 21684
rect 22465 21675 22523 21681
rect 22465 21641 22477 21675
rect 22511 21672 22523 21675
rect 23474 21672 23480 21684
rect 22511 21644 23480 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 23474 21632 23480 21644
rect 23532 21632 23538 21684
rect 23566 21632 23572 21684
rect 23624 21672 23630 21684
rect 25409 21675 25467 21681
rect 25409 21672 25421 21675
rect 23624 21644 25421 21672
rect 23624 21632 23630 21644
rect 7650 21564 7656 21616
rect 7708 21604 7714 21616
rect 7708 21576 10088 21604
rect 7708 21564 7714 21576
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21536 1823 21539
rect 1854 21536 1860 21548
rect 1811 21508 1860 21536
rect 1811 21505 1823 21508
rect 1765 21499 1823 21505
rect 1854 21496 1860 21508
rect 1912 21496 1918 21548
rect 3421 21539 3479 21545
rect 3421 21505 3433 21539
rect 3467 21536 3479 21539
rect 4154 21536 4160 21548
rect 3467 21508 4160 21536
rect 3467 21505 3479 21508
rect 3421 21499 3479 21505
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 4522 21496 4528 21548
rect 4580 21496 4586 21548
rect 7561 21539 7619 21545
rect 7561 21505 7573 21539
rect 7607 21536 7619 21539
rect 8938 21536 8944 21548
rect 7607 21508 8944 21536
rect 7607 21505 7619 21508
rect 7561 21499 7619 21505
rect 8938 21496 8944 21508
rect 8996 21496 9002 21548
rect 1302 21428 1308 21480
rect 1360 21468 1366 21480
rect 2041 21471 2099 21477
rect 2041 21468 2053 21471
rect 1360 21440 2053 21468
rect 1360 21428 1366 21440
rect 2041 21437 2053 21440
rect 2087 21437 2099 21471
rect 2041 21431 2099 21437
rect 3602 21428 3608 21480
rect 3660 21468 3666 21480
rect 4062 21468 4068 21480
rect 3660 21440 4068 21468
rect 3660 21428 3666 21440
rect 4062 21428 4068 21440
rect 4120 21468 4126 21480
rect 4985 21471 5043 21477
rect 4985 21468 4997 21471
rect 4120 21440 4997 21468
rect 4120 21428 4126 21440
rect 4985 21437 4997 21440
rect 5031 21437 5043 21471
rect 4985 21431 5043 21437
rect 7650 21428 7656 21480
rect 7708 21428 7714 21480
rect 8754 21428 8760 21480
rect 8812 21428 8818 21480
rect 8849 21471 8907 21477
rect 8849 21437 8861 21471
rect 8895 21468 8907 21471
rect 9122 21468 9128 21480
rect 8895 21440 9128 21468
rect 8895 21437 8907 21440
rect 8849 21431 8907 21437
rect 9122 21428 9128 21440
rect 9180 21428 9186 21480
rect 10060 21477 10088 21576
rect 13630 21564 13636 21616
rect 13688 21604 13694 21616
rect 14001 21607 14059 21613
rect 14001 21604 14013 21607
rect 13688 21576 14013 21604
rect 13688 21564 13694 21576
rect 14001 21573 14013 21576
rect 14047 21573 14059 21607
rect 14001 21567 14059 21573
rect 14108 21576 17080 21604
rect 12161 21539 12219 21545
rect 12161 21505 12173 21539
rect 12207 21536 12219 21539
rect 13814 21536 13820 21548
rect 12207 21508 13820 21536
rect 12207 21505 12219 21508
rect 12161 21499 12219 21505
rect 13814 21496 13820 21508
rect 13872 21496 13878 21548
rect 9953 21471 10011 21477
rect 9953 21437 9965 21471
rect 9999 21437 10011 21471
rect 9953 21431 10011 21437
rect 10045 21471 10103 21477
rect 10045 21437 10057 21471
rect 10091 21437 10103 21471
rect 10045 21431 10103 21437
rect 3786 21360 3792 21412
rect 3844 21360 3850 21412
rect 6914 21360 6920 21412
rect 6972 21400 6978 21412
rect 9493 21403 9551 21409
rect 9493 21400 9505 21403
rect 6972 21372 9505 21400
rect 6972 21360 6978 21372
rect 9493 21369 9505 21372
rect 9539 21369 9551 21403
rect 9968 21400 9996 21431
rect 11882 21428 11888 21480
rect 11940 21468 11946 21480
rect 12253 21471 12311 21477
rect 12253 21468 12265 21471
rect 11940 21440 12265 21468
rect 11940 21428 11946 21440
rect 12253 21437 12265 21440
rect 12299 21437 12311 21471
rect 12253 21431 12311 21437
rect 13722 21428 13728 21480
rect 13780 21468 13786 21480
rect 14108 21468 14136 21576
rect 15194 21496 15200 21548
rect 15252 21496 15258 21548
rect 17052 21545 17080 21576
rect 22002 21564 22008 21616
rect 22060 21604 22066 21616
rect 22060 21576 23428 21604
rect 22060 21564 22066 21576
rect 16209 21539 16267 21545
rect 16209 21505 16221 21539
rect 16255 21505 16267 21539
rect 16209 21499 16267 21505
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21505 17095 21539
rect 17037 21499 17095 21505
rect 13780 21440 14136 21468
rect 13780 21428 13786 21440
rect 14182 21428 14188 21480
rect 14240 21428 14246 21480
rect 14458 21428 14464 21480
rect 14516 21468 14522 21480
rect 15102 21468 15108 21480
rect 14516 21440 15108 21468
rect 14516 21428 14522 21440
rect 15102 21428 15108 21440
rect 15160 21468 15166 21480
rect 15289 21471 15347 21477
rect 15289 21468 15301 21471
rect 15160 21440 15301 21468
rect 15160 21428 15166 21440
rect 15289 21437 15301 21440
rect 15335 21437 15347 21471
rect 15289 21431 15347 21437
rect 15470 21428 15476 21480
rect 15528 21428 15534 21480
rect 11514 21400 11520 21412
rect 9968 21372 11520 21400
rect 9493 21363 9551 21369
rect 11514 21360 11520 21372
rect 11572 21360 11578 21412
rect 12342 21360 12348 21412
rect 12400 21400 12406 21412
rect 16224 21400 16252 21499
rect 17402 21496 17408 21548
rect 17460 21536 17466 21548
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 17460 21508 18705 21536
rect 17460 21496 17466 21508
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 19978 21496 19984 21548
rect 20036 21536 20042 21548
rect 22830 21536 22836 21548
rect 20036 21508 22836 21536
rect 20036 21496 20042 21508
rect 22830 21496 22836 21508
rect 22888 21496 22894 21548
rect 23400 21545 23428 21576
rect 23658 21564 23664 21616
rect 23716 21564 23722 21616
rect 24044 21604 24072 21644
rect 25409 21641 25421 21644
rect 25455 21641 25467 21675
rect 25409 21635 25467 21641
rect 24044 21576 24150 21604
rect 23385 21539 23443 21545
rect 23385 21505 23397 21539
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 17586 21428 17592 21480
rect 17644 21468 17650 21480
rect 17681 21471 17739 21477
rect 17681 21468 17693 21471
rect 17644 21440 17693 21468
rect 17644 21428 17650 21440
rect 17681 21437 17693 21440
rect 17727 21437 17739 21471
rect 17681 21431 17739 21437
rect 17770 21428 17776 21480
rect 17828 21468 17834 21480
rect 17828 21440 18828 21468
rect 17828 21428 17834 21440
rect 12400 21372 16252 21400
rect 16853 21403 16911 21409
rect 12400 21360 12406 21372
rect 16853 21369 16865 21403
rect 16899 21400 16911 21403
rect 18690 21400 18696 21412
rect 16899 21372 18696 21400
rect 16899 21369 16911 21372
rect 16853 21363 16911 21369
rect 18690 21360 18696 21372
rect 18748 21360 18754 21412
rect 18800 21400 18828 21440
rect 20162 21428 20168 21480
rect 20220 21468 20226 21480
rect 20438 21468 20444 21480
rect 20220 21440 20444 21468
rect 20220 21428 20226 21440
rect 20438 21428 20444 21440
rect 20496 21428 20502 21480
rect 22554 21428 22560 21480
rect 22612 21428 22618 21480
rect 22646 21428 22652 21480
rect 22704 21468 22710 21480
rect 22741 21471 22799 21477
rect 22741 21468 22753 21471
rect 22704 21440 22753 21468
rect 22704 21428 22710 21440
rect 22741 21437 22753 21440
rect 22787 21468 22799 21471
rect 22787 21440 23520 21468
rect 22787 21437 22799 21440
rect 22741 21431 22799 21437
rect 20254 21400 20260 21412
rect 18800 21372 20260 21400
rect 20254 21360 20260 21372
rect 20312 21400 20318 21412
rect 20898 21400 20904 21412
rect 20312 21372 20904 21400
rect 20312 21360 20318 21372
rect 20898 21360 20904 21372
rect 20956 21360 20962 21412
rect 4801 21335 4859 21341
rect 4801 21301 4813 21335
rect 4847 21332 4859 21335
rect 5810 21332 5816 21344
rect 4847 21304 5816 21332
rect 4847 21301 4859 21304
rect 4801 21295 4859 21301
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 10318 21292 10324 21344
rect 10376 21332 10382 21344
rect 10870 21332 10876 21344
rect 10376 21304 10876 21332
rect 10376 21292 10382 21304
rect 10870 21292 10876 21304
rect 10928 21292 10934 21344
rect 13446 21292 13452 21344
rect 13504 21332 13510 21344
rect 14829 21335 14887 21341
rect 14829 21332 14841 21335
rect 13504 21304 14841 21332
rect 13504 21292 13510 21304
rect 14829 21301 14841 21304
rect 14875 21301 14887 21335
rect 14829 21295 14887 21301
rect 15286 21292 15292 21344
rect 15344 21332 15350 21344
rect 15470 21332 15476 21344
rect 15344 21304 15476 21332
rect 15344 21292 15350 21304
rect 15470 21292 15476 21304
rect 15528 21292 15534 21344
rect 18509 21335 18567 21341
rect 18509 21301 18521 21335
rect 18555 21332 18567 21335
rect 19058 21332 19064 21344
rect 18555 21304 19064 21332
rect 18555 21301 18567 21304
rect 18509 21295 18567 21301
rect 19058 21292 19064 21304
rect 19116 21292 19122 21344
rect 20438 21292 20444 21344
rect 20496 21292 20502 21344
rect 22097 21335 22155 21341
rect 22097 21301 22109 21335
rect 22143 21332 22155 21335
rect 22278 21332 22284 21344
rect 22143 21304 22284 21332
rect 22143 21301 22155 21304
rect 22097 21295 22155 21301
rect 22278 21292 22284 21304
rect 22336 21292 22342 21344
rect 23492 21332 23520 21440
rect 25133 21335 25191 21341
rect 25133 21332 25145 21335
rect 23492 21304 25145 21332
rect 25133 21301 25145 21304
rect 25179 21301 25191 21335
rect 25133 21295 25191 21301
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 2866 21088 2872 21140
rect 2924 21128 2930 21140
rect 3145 21131 3203 21137
rect 3145 21128 3157 21131
rect 2924 21100 3157 21128
rect 2924 21088 2930 21100
rect 3145 21097 3157 21100
rect 3191 21097 3203 21131
rect 3145 21091 3203 21097
rect 7282 21088 7288 21140
rect 7340 21128 7346 21140
rect 7837 21131 7895 21137
rect 7837 21128 7849 21131
rect 7340 21100 7849 21128
rect 7340 21088 7346 21100
rect 7837 21097 7849 21100
rect 7883 21097 7895 21131
rect 7837 21091 7895 21097
rect 12066 21088 12072 21140
rect 12124 21128 12130 21140
rect 14458 21128 14464 21140
rect 12124 21100 14464 21128
rect 12124 21088 12130 21100
rect 14458 21088 14464 21100
rect 14516 21088 14522 21140
rect 16574 21088 16580 21140
rect 16632 21128 16638 21140
rect 16853 21131 16911 21137
rect 16853 21128 16865 21131
rect 16632 21100 16865 21128
rect 16632 21088 16638 21100
rect 16853 21097 16865 21100
rect 16899 21097 16911 21131
rect 19978 21128 19984 21140
rect 16853 21091 16911 21097
rect 17144 21100 19984 21128
rect 4065 21063 4123 21069
rect 4065 21029 4077 21063
rect 4111 21029 4123 21063
rect 4065 21023 4123 21029
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20992 2835 20995
rect 4080 20992 4108 21023
rect 15194 21020 15200 21072
rect 15252 21060 15258 21072
rect 16117 21063 16175 21069
rect 16117 21060 16129 21063
rect 15252 21032 16129 21060
rect 15252 21020 15258 21032
rect 16117 21029 16129 21032
rect 16163 21060 16175 21063
rect 17144 21060 17172 21100
rect 19978 21088 19984 21100
rect 20036 21128 20042 21140
rect 21542 21128 21548 21140
rect 20036 21100 21548 21128
rect 20036 21088 20042 21100
rect 21542 21088 21548 21100
rect 21600 21088 21606 21140
rect 16163 21032 17172 21060
rect 17221 21063 17279 21069
rect 16163 21029 16175 21032
rect 16117 21023 16175 21029
rect 17221 21029 17233 21063
rect 17267 21060 17279 21063
rect 19334 21060 19340 21072
rect 17267 21032 19340 21060
rect 17267 21029 17279 21032
rect 17221 21023 17279 21029
rect 19334 21020 19340 21032
rect 19392 21020 19398 21072
rect 21450 21020 21456 21072
rect 21508 21060 21514 21072
rect 21913 21063 21971 21069
rect 21913 21060 21925 21063
rect 21508 21032 21925 21060
rect 21508 21020 21514 21032
rect 21913 21029 21925 21032
rect 21959 21060 21971 21063
rect 22554 21060 22560 21072
rect 21959 21032 22560 21060
rect 21959 21029 21971 21032
rect 21913 21023 21971 21029
rect 22554 21020 22560 21032
rect 22612 21020 22618 21072
rect 2823 20964 4108 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 7834 20952 7840 21004
rect 7892 20992 7898 21004
rect 8481 20995 8539 21001
rect 8481 20992 8493 20995
rect 7892 20964 8493 20992
rect 7892 20952 7898 20964
rect 8481 20961 8493 20964
rect 8527 20992 8539 20995
rect 10042 20992 10048 21004
rect 8527 20964 10048 20992
rect 8527 20961 8539 20964
rect 8481 20955 8539 20961
rect 10042 20952 10048 20964
rect 10100 20992 10106 21004
rect 11517 20995 11575 21001
rect 11517 20992 11529 20995
rect 10100 20964 11529 20992
rect 10100 20952 10106 20964
rect 11517 20961 11529 20964
rect 11563 20992 11575 20995
rect 11882 20992 11888 21004
rect 11563 20964 11888 20992
rect 11563 20961 11575 20964
rect 11517 20955 11575 20961
rect 11882 20952 11888 20964
rect 11940 20952 11946 21004
rect 14921 20995 14979 21001
rect 14921 20992 14933 20995
rect 14292 20964 14933 20992
rect 14292 20936 14320 20964
rect 14921 20961 14933 20964
rect 14967 20961 14979 20995
rect 16301 20995 16359 21001
rect 16301 20992 16313 20995
rect 14921 20955 14979 20961
rect 15672 20964 16313 20992
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20893 2283 20927
rect 2225 20887 2283 20893
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20924 3019 20927
rect 4062 20924 4068 20936
rect 3007 20896 4068 20924
rect 3007 20893 3019 20896
rect 2961 20887 3019 20893
rect 2240 20856 2268 20887
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 4246 20884 4252 20936
rect 4304 20884 4310 20936
rect 9769 20927 9827 20933
rect 9769 20893 9781 20927
rect 9815 20893 9827 20927
rect 11330 20924 11336 20936
rect 11178 20896 11336 20924
rect 9769 20887 9827 20893
rect 8662 20856 8668 20868
rect 2240 20828 2774 20856
rect 2746 20800 2774 20828
rect 8220 20828 8668 20856
rect 1762 20748 1768 20800
rect 1820 20788 1826 20800
rect 2041 20791 2099 20797
rect 2041 20788 2053 20791
rect 1820 20760 2053 20788
rect 1820 20748 1826 20760
rect 2041 20757 2053 20760
rect 2087 20757 2099 20791
rect 2746 20760 2780 20800
rect 2041 20751 2099 20757
rect 2774 20748 2780 20760
rect 2832 20748 2838 20800
rect 5442 20748 5448 20800
rect 5500 20788 5506 20800
rect 8220 20797 8248 20828
rect 8662 20816 8668 20828
rect 8720 20816 8726 20868
rect 9784 20856 9812 20887
rect 11330 20884 11336 20896
rect 11388 20924 11394 20936
rect 11977 20927 12035 20933
rect 11977 20924 11989 20927
rect 11388 20896 11989 20924
rect 11388 20884 11394 20896
rect 11977 20893 11989 20896
rect 12023 20893 12035 20927
rect 14274 20924 14280 20936
rect 11977 20887 12035 20893
rect 13832 20896 14280 20924
rect 9950 20856 9956 20868
rect 9784 20828 9956 20856
rect 9950 20816 9956 20828
rect 10008 20816 10014 20868
rect 10045 20859 10103 20865
rect 10045 20825 10057 20859
rect 10091 20856 10103 20859
rect 10318 20856 10324 20868
rect 10091 20828 10324 20856
rect 10091 20825 10103 20828
rect 10045 20819 10103 20825
rect 10318 20816 10324 20828
rect 10376 20816 10382 20868
rect 13832 20856 13860 20896
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 14737 20927 14795 20933
rect 14737 20893 14749 20927
rect 14783 20924 14795 20927
rect 15672 20924 15700 20964
rect 16301 20961 16313 20964
rect 16347 20992 16359 20995
rect 17770 20992 17776 21004
rect 16347 20964 17776 20992
rect 16347 20961 16359 20964
rect 16301 20955 16359 20961
rect 17770 20952 17776 20964
rect 17828 20952 17834 21004
rect 17865 20995 17923 21001
rect 17865 20961 17877 20995
rect 17911 20992 17923 20995
rect 17911 20964 19380 20992
rect 17911 20961 17923 20964
rect 17865 20955 17923 20961
rect 14783 20896 15700 20924
rect 14783 20893 14795 20896
rect 14737 20887 14795 20893
rect 15746 20884 15752 20936
rect 15804 20884 15810 20936
rect 17586 20884 17592 20936
rect 17644 20884 17650 20936
rect 17678 20884 17684 20936
rect 17736 20924 17742 20936
rect 18877 20927 18935 20933
rect 18877 20924 18889 20927
rect 17736 20896 18889 20924
rect 17736 20884 17742 20896
rect 18877 20893 18889 20896
rect 18923 20893 18935 20927
rect 18877 20887 18935 20893
rect 14826 20856 14832 20868
rect 11348 20828 13860 20856
rect 13924 20828 14832 20856
rect 7469 20791 7527 20797
rect 7469 20788 7481 20791
rect 5500 20760 7481 20788
rect 5500 20748 5506 20760
rect 7469 20757 7481 20760
rect 7515 20788 7527 20791
rect 8205 20791 8263 20797
rect 8205 20788 8217 20791
rect 7515 20760 8217 20788
rect 7515 20757 7527 20760
rect 7469 20751 7527 20757
rect 8205 20757 8217 20760
rect 8251 20757 8263 20791
rect 8205 20751 8263 20757
rect 8297 20791 8355 20797
rect 8297 20757 8309 20791
rect 8343 20788 8355 20791
rect 10410 20788 10416 20800
rect 8343 20760 10416 20788
rect 8343 20757 8355 20760
rect 8297 20751 8355 20757
rect 10410 20748 10416 20760
rect 10468 20748 10474 20800
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 11348 20788 11376 20828
rect 13924 20800 13952 20828
rect 14826 20816 14832 20828
rect 14884 20816 14890 20868
rect 15378 20816 15384 20868
rect 15436 20856 15442 20868
rect 16758 20856 16764 20868
rect 15436 20828 16764 20856
rect 15436 20816 15442 20828
rect 16758 20816 16764 20828
rect 16816 20816 16822 20868
rect 19352 20856 19380 20964
rect 19426 20952 19432 21004
rect 19484 20992 19490 21004
rect 19889 20995 19947 21001
rect 19889 20992 19901 20995
rect 19484 20964 19901 20992
rect 19484 20952 19490 20964
rect 19889 20961 19901 20964
rect 19935 20961 19947 20995
rect 19889 20955 19947 20961
rect 20714 20952 20720 21004
rect 20772 20992 20778 21004
rect 23845 20995 23903 21001
rect 20772 20964 21312 20992
rect 20772 20952 20778 20964
rect 21284 20924 21312 20964
rect 23845 20961 23857 20995
rect 23891 20992 23903 20995
rect 24854 20992 24860 21004
rect 23891 20964 24860 20992
rect 23891 20961 23903 20964
rect 23845 20955 23903 20961
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 21450 20924 21456 20936
rect 21284 20910 21456 20924
rect 21298 20896 21456 20910
rect 21450 20884 21456 20896
rect 21508 20884 21514 20936
rect 22186 20884 22192 20936
rect 22244 20924 22250 20936
rect 22649 20927 22707 20933
rect 22649 20924 22661 20927
rect 22244 20896 22661 20924
rect 22244 20884 22250 20896
rect 22649 20893 22661 20896
rect 22695 20893 22707 20927
rect 22649 20887 22707 20893
rect 20162 20856 20168 20868
rect 19352 20828 20168 20856
rect 20162 20816 20168 20828
rect 20220 20816 20226 20868
rect 24854 20856 24860 20868
rect 21468 20828 24860 20856
rect 11020 20760 11376 20788
rect 11020 20748 11026 20760
rect 13906 20748 13912 20800
rect 13964 20748 13970 20800
rect 14366 20748 14372 20800
rect 14424 20748 14430 20800
rect 15470 20748 15476 20800
rect 15528 20788 15534 20800
rect 15565 20791 15623 20797
rect 15565 20788 15577 20791
rect 15528 20760 15577 20788
rect 15528 20748 15534 20760
rect 15565 20757 15577 20760
rect 15611 20757 15623 20791
rect 15565 20751 15623 20757
rect 16574 20748 16580 20800
rect 16632 20788 16638 20800
rect 17681 20791 17739 20797
rect 17681 20788 17693 20791
rect 16632 20760 17693 20788
rect 16632 20748 16638 20760
rect 17681 20757 17693 20760
rect 17727 20757 17739 20791
rect 17681 20751 17739 20757
rect 18693 20791 18751 20797
rect 18693 20757 18705 20791
rect 18739 20788 18751 20791
rect 21468 20788 21496 20828
rect 24854 20816 24860 20828
rect 24912 20816 24918 20868
rect 18739 20760 21496 20788
rect 18739 20757 18751 20760
rect 18693 20751 18751 20757
rect 21634 20748 21640 20800
rect 21692 20748 21698 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 6546 20544 6552 20596
rect 6604 20584 6610 20596
rect 8846 20584 8852 20596
rect 6604 20556 8852 20584
rect 6604 20544 6610 20556
rect 8846 20544 8852 20556
rect 8904 20544 8910 20596
rect 8938 20544 8944 20596
rect 8996 20584 9002 20596
rect 9953 20587 10011 20593
rect 9953 20584 9965 20587
rect 8996 20556 9965 20584
rect 8996 20544 9002 20556
rect 9953 20553 9965 20556
rect 9999 20553 10011 20587
rect 11974 20584 11980 20596
rect 9953 20547 10011 20553
rect 10060 20556 11980 20584
rect 4249 20519 4307 20525
rect 4249 20485 4261 20519
rect 4295 20516 4307 20519
rect 4338 20516 4344 20528
rect 4295 20488 4344 20516
rect 4295 20485 4307 20488
rect 4249 20479 4307 20485
rect 4338 20476 4344 20488
rect 4396 20476 4402 20528
rect 5997 20519 6055 20525
rect 5997 20516 6009 20519
rect 5474 20488 6009 20516
rect 5997 20485 6009 20488
rect 6043 20516 6055 20519
rect 7098 20516 7104 20528
rect 6043 20488 7104 20516
rect 6043 20485 6055 20488
rect 5997 20479 6055 20485
rect 7098 20476 7104 20488
rect 7156 20516 7162 20528
rect 7156 20488 7314 20516
rect 8864 20488 9444 20516
rect 7156 20476 7162 20488
rect 3973 20451 4031 20457
rect 3973 20417 3985 20451
rect 4019 20417 4031 20451
rect 3973 20411 4031 20417
rect 3988 20380 4016 20411
rect 6546 20408 6552 20460
rect 6604 20408 6610 20460
rect 5718 20380 5724 20392
rect 3988 20352 5724 20380
rect 5718 20340 5724 20352
rect 5776 20340 5782 20392
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 8864 20380 8892 20488
rect 8938 20408 8944 20460
rect 8996 20448 9002 20460
rect 9125 20451 9183 20457
rect 9125 20448 9137 20451
rect 8996 20420 9137 20448
rect 8996 20408 9002 20420
rect 9125 20417 9137 20420
rect 9171 20417 9183 20451
rect 9125 20411 9183 20417
rect 9416 20448 9444 20488
rect 10060 20448 10088 20556
rect 11974 20544 11980 20556
rect 12032 20544 12038 20596
rect 12529 20587 12587 20593
rect 12529 20553 12541 20587
rect 12575 20584 12587 20587
rect 13630 20584 13636 20596
rect 12575 20556 13636 20584
rect 12575 20553 12587 20556
rect 12529 20547 12587 20553
rect 13630 20544 13636 20556
rect 13688 20584 13694 20596
rect 13998 20584 14004 20596
rect 13688 20556 14004 20584
rect 13688 20544 13694 20556
rect 13998 20544 14004 20556
rect 14056 20544 14062 20596
rect 17310 20544 17316 20596
rect 17368 20584 17374 20596
rect 17368 20556 17724 20584
rect 17368 20544 17374 20556
rect 10413 20519 10471 20525
rect 10413 20485 10425 20519
rect 10459 20516 10471 20519
rect 10962 20516 10968 20528
rect 10459 20488 10968 20516
rect 10459 20485 10471 20488
rect 10413 20479 10471 20485
rect 10962 20476 10968 20488
rect 11020 20476 11026 20528
rect 12250 20476 12256 20528
rect 12308 20516 12314 20528
rect 17696 20525 17724 20556
rect 19334 20544 19340 20596
rect 19392 20544 19398 20596
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 19518 20584 19524 20596
rect 19475 20556 19524 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 17681 20519 17739 20525
rect 12308 20488 15700 20516
rect 12308 20476 12314 20488
rect 9416 20420 10088 20448
rect 10321 20451 10379 20457
rect 9416 20389 9444 20420
rect 10321 20417 10333 20451
rect 10367 20448 10379 20451
rect 11698 20448 11704 20460
rect 10367 20420 11704 20448
rect 10367 20417 10379 20420
rect 10321 20411 10379 20417
rect 11698 20408 11704 20420
rect 11756 20408 11762 20460
rect 15672 20457 15700 20488
rect 17681 20485 17693 20519
rect 17727 20485 17739 20519
rect 17681 20479 17739 20485
rect 23293 20519 23351 20525
rect 23293 20485 23305 20519
rect 23339 20516 23351 20519
rect 23382 20516 23388 20528
rect 23339 20488 23388 20516
rect 23339 20485 23351 20488
rect 23293 20479 23351 20485
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 12437 20451 12495 20457
rect 12437 20417 12449 20451
rect 12483 20448 12495 20451
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 12483 20420 13277 20448
rect 12483 20417 12495 20420
rect 12437 20411 12495 20417
rect 13265 20417 13277 20420
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 15657 20451 15715 20457
rect 15657 20417 15669 20451
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 18509 20451 18567 20457
rect 18509 20417 18521 20451
rect 18555 20448 18567 20451
rect 19150 20448 19156 20460
rect 18555 20420 19156 20448
rect 18555 20417 18567 20420
rect 18509 20411 18567 20417
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 22281 20451 22339 20457
rect 22281 20417 22293 20451
rect 22327 20448 22339 20451
rect 22370 20448 22376 20460
rect 22327 20420 22376 20448
rect 22327 20417 22339 20420
rect 22281 20411 22339 20417
rect 22370 20408 22376 20420
rect 22428 20408 22434 20460
rect 24121 20451 24179 20457
rect 24121 20417 24133 20451
rect 24167 20448 24179 20451
rect 25038 20448 25044 20460
rect 24167 20420 25044 20448
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 25038 20408 25044 20420
rect 25096 20408 25102 20460
rect 6871 20352 8892 20380
rect 9217 20383 9275 20389
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 9217 20349 9229 20383
rect 9263 20349 9275 20383
rect 9217 20343 9275 20349
rect 9401 20383 9459 20389
rect 9401 20349 9413 20383
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 8754 20272 8760 20324
rect 8812 20272 8818 20324
rect 9232 20312 9260 20343
rect 9582 20340 9588 20392
rect 9640 20380 9646 20392
rect 10505 20383 10563 20389
rect 10505 20380 10517 20383
rect 9640 20352 10517 20380
rect 9640 20340 9646 20352
rect 10505 20349 10517 20352
rect 10551 20349 10563 20383
rect 10505 20343 10563 20349
rect 11146 20340 11152 20392
rect 11204 20380 11210 20392
rect 11204 20352 12434 20380
rect 11204 20340 11210 20352
rect 11606 20312 11612 20324
rect 9232 20284 11612 20312
rect 11606 20272 11612 20284
rect 11664 20272 11670 20324
rect 12406 20312 12434 20352
rect 12710 20340 12716 20392
rect 12768 20340 12774 20392
rect 19613 20383 19671 20389
rect 19613 20349 19625 20383
rect 19659 20380 19671 20383
rect 21634 20380 21640 20392
rect 19659 20352 21640 20380
rect 19659 20349 19671 20352
rect 19613 20343 19671 20349
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 24397 20383 24455 20389
rect 24397 20380 24409 20383
rect 23348 20352 24409 20380
rect 23348 20340 23354 20352
rect 24397 20349 24409 20352
rect 24443 20349 24455 20383
rect 24397 20343 24455 20349
rect 17034 20312 17040 20324
rect 12406 20284 17040 20312
rect 17034 20272 17040 20284
rect 17092 20272 17098 20324
rect 5721 20247 5779 20253
rect 5721 20213 5733 20247
rect 5767 20244 5779 20247
rect 5810 20244 5816 20256
rect 5767 20216 5816 20244
rect 5767 20213 5779 20216
rect 5721 20207 5779 20213
rect 5810 20204 5816 20216
rect 5868 20204 5874 20256
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 9122 20244 9128 20256
rect 8352 20216 9128 20244
rect 8352 20204 8358 20216
rect 9122 20204 9128 20216
rect 9180 20244 9186 20256
rect 9582 20244 9588 20256
rect 9180 20216 9588 20244
rect 9180 20204 9186 20216
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 12066 20204 12072 20256
rect 12124 20204 12130 20256
rect 13630 20204 13636 20256
rect 13688 20244 13694 20256
rect 13725 20247 13783 20253
rect 13725 20244 13737 20247
rect 13688 20216 13737 20244
rect 13688 20204 13694 20216
rect 13725 20213 13737 20216
rect 13771 20213 13783 20247
rect 13725 20207 13783 20213
rect 14737 20247 14795 20253
rect 14737 20213 14749 20247
rect 14783 20244 14795 20247
rect 15102 20244 15108 20256
rect 14783 20216 15108 20244
rect 14783 20213 14795 20216
rect 14737 20207 14795 20213
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 15470 20204 15476 20256
rect 15528 20204 15534 20256
rect 16850 20204 16856 20256
rect 16908 20244 16914 20256
rect 17773 20247 17831 20253
rect 17773 20244 17785 20247
rect 16908 20216 17785 20244
rect 16908 20204 16914 20216
rect 17773 20213 17785 20216
rect 17819 20213 17831 20247
rect 17773 20207 17831 20213
rect 18325 20247 18383 20253
rect 18325 20213 18337 20247
rect 18371 20244 18383 20247
rect 18414 20244 18420 20256
rect 18371 20216 18420 20244
rect 18371 20213 18383 20216
rect 18325 20207 18383 20213
rect 18414 20204 18420 20216
rect 18472 20204 18478 20256
rect 18969 20247 19027 20253
rect 18969 20213 18981 20247
rect 19015 20244 19027 20247
rect 19794 20244 19800 20256
rect 19015 20216 19800 20244
rect 19015 20213 19027 20216
rect 18969 20207 19027 20213
rect 19794 20204 19800 20216
rect 19852 20204 19858 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 5074 20000 5080 20052
rect 5132 20000 5138 20052
rect 5718 20000 5724 20052
rect 5776 20040 5782 20052
rect 6546 20040 6552 20052
rect 5776 20012 6552 20040
rect 5776 20000 5782 20012
rect 6546 20000 6552 20012
rect 6604 20000 6610 20052
rect 11698 20000 11704 20052
rect 11756 20000 11762 20052
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 12250 20040 12256 20052
rect 12032 20012 12256 20040
rect 12032 20000 12038 20012
rect 12250 20000 12256 20012
rect 12308 20000 12314 20052
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 13872 20012 14289 20040
rect 13872 20000 13878 20012
rect 14277 20009 14289 20012
rect 14323 20009 14335 20043
rect 14277 20003 14335 20009
rect 20349 20043 20407 20049
rect 20349 20009 20361 20043
rect 20395 20040 20407 20043
rect 20806 20040 20812 20052
rect 20395 20012 20812 20040
rect 20395 20009 20407 20012
rect 20349 20003 20407 20009
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 5736 19913 5764 20000
rect 12158 19932 12164 19984
rect 12216 19972 12222 19984
rect 12618 19972 12624 19984
rect 12216 19944 12624 19972
rect 12216 19932 12222 19944
rect 12618 19932 12624 19944
rect 12676 19932 12682 19984
rect 15381 19975 15439 19981
rect 15381 19941 15393 19975
rect 15427 19972 15439 19975
rect 18782 19972 18788 19984
rect 15427 19944 18788 19972
rect 15427 19941 15439 19944
rect 15381 19935 15439 19941
rect 5721 19907 5779 19913
rect 5721 19873 5733 19907
rect 5767 19873 5779 19907
rect 5721 19867 5779 19873
rect 5997 19907 6055 19913
rect 5997 19873 6009 19907
rect 6043 19904 6055 19907
rect 8294 19904 8300 19916
rect 6043 19876 8300 19904
rect 6043 19873 6055 19876
rect 5997 19867 6055 19873
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 8846 19864 8852 19916
rect 8904 19904 8910 19916
rect 9125 19907 9183 19913
rect 9125 19904 9137 19907
rect 8904 19876 9137 19904
rect 8904 19864 8910 19876
rect 9125 19873 9137 19876
rect 9171 19873 9183 19907
rect 9125 19867 9183 19873
rect 11149 19907 11207 19913
rect 11149 19873 11161 19907
rect 11195 19904 11207 19907
rect 12176 19904 12204 19932
rect 11195 19876 12204 19904
rect 11195 19873 11207 19876
rect 11149 19867 11207 19873
rect 12250 19864 12256 19916
rect 12308 19864 12314 19916
rect 14182 19864 14188 19916
rect 14240 19904 14246 19916
rect 14829 19907 14887 19913
rect 14829 19904 14841 19907
rect 14240 19876 14841 19904
rect 14240 19864 14246 19876
rect 14829 19873 14841 19876
rect 14875 19873 14887 19907
rect 14829 19867 14887 19873
rect 5261 19839 5319 19845
rect 5261 19805 5273 19839
rect 5307 19805 5319 19839
rect 5261 19799 5319 19805
rect 5276 19700 5304 19799
rect 7098 19796 7104 19848
rect 7156 19836 7162 19848
rect 7742 19836 7748 19848
rect 7156 19808 7748 19836
rect 7156 19796 7162 19808
rect 7742 19796 7748 19808
rect 7800 19836 7806 19848
rect 8202 19836 8208 19848
rect 7800 19808 8208 19836
rect 7800 19796 7806 19808
rect 8202 19796 8208 19808
rect 8260 19836 8266 19848
rect 8389 19839 8447 19845
rect 8389 19836 8401 19839
rect 8260 19808 8401 19836
rect 8260 19796 8266 19808
rect 8389 19805 8401 19808
rect 8435 19836 8447 19839
rect 9030 19836 9036 19848
rect 8435 19808 9036 19836
rect 8435 19805 8447 19808
rect 8389 19799 8447 19805
rect 9030 19796 9036 19808
rect 9088 19796 9094 19848
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19836 12127 19839
rect 12434 19836 12440 19848
rect 12115 19808 12440 19836
rect 12115 19805 12127 19808
rect 12069 19799 12127 19805
rect 12434 19796 12440 19808
rect 12492 19796 12498 19848
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19836 14703 19839
rect 15396 19836 15424 19935
rect 18782 19932 18788 19944
rect 18840 19972 18846 19984
rect 20254 19972 20260 19984
rect 18840 19944 20260 19972
rect 18840 19932 18846 19944
rect 20254 19932 20260 19944
rect 20312 19932 20318 19984
rect 17862 19864 17868 19916
rect 17920 19904 17926 19916
rect 23845 19907 23903 19913
rect 17920 19876 22048 19904
rect 17920 19864 17926 19876
rect 14691 19808 15424 19836
rect 17221 19839 17279 19845
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 17221 19805 17233 19839
rect 17267 19836 17279 19839
rect 17770 19836 17776 19848
rect 17267 19808 17776 19836
rect 17267 19805 17279 19808
rect 17221 19799 17279 19805
rect 17770 19796 17776 19808
rect 17828 19796 17834 19848
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19836 18751 19839
rect 18874 19836 18880 19848
rect 18739 19808 18880 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 18874 19796 18880 19808
rect 18932 19796 18938 19848
rect 22020 19845 22048 19876
rect 23845 19873 23857 19907
rect 23891 19904 23903 19907
rect 24946 19904 24952 19916
rect 23891 19876 24952 19904
rect 23891 19873 23903 19876
rect 23845 19867 23903 19873
rect 24946 19864 24952 19876
rect 25004 19864 25010 19916
rect 22005 19839 22063 19845
rect 22005 19805 22017 19839
rect 22051 19805 22063 19839
rect 22005 19799 22063 19805
rect 22833 19839 22891 19845
rect 22833 19805 22845 19839
rect 22879 19836 22891 19839
rect 25222 19836 25228 19848
rect 22879 19808 25228 19836
rect 22879 19805 22891 19808
rect 22833 19799 22891 19805
rect 25222 19796 25228 19808
rect 25280 19796 25286 19848
rect 7650 19768 7656 19780
rect 7484 19740 7656 19768
rect 7282 19700 7288 19712
rect 5276 19672 7288 19700
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 7484 19709 7512 19740
rect 7650 19728 7656 19740
rect 7708 19768 7714 19780
rect 9401 19771 9459 19777
rect 9401 19768 9413 19771
rect 7708 19740 9413 19768
rect 7708 19728 7714 19740
rect 9401 19737 9413 19740
rect 9447 19737 9459 19771
rect 9401 19731 9459 19737
rect 9508 19740 9890 19768
rect 7469 19703 7527 19709
rect 7469 19669 7481 19703
rect 7515 19669 7527 19703
rect 7469 19663 7527 19669
rect 8665 19703 8723 19709
rect 8665 19669 8677 19703
rect 8711 19700 8723 19703
rect 8846 19700 8852 19712
rect 8711 19672 8852 19700
rect 8711 19669 8723 19672
rect 8665 19663 8723 19669
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 9030 19660 9036 19712
rect 9088 19700 9094 19712
rect 9508 19700 9536 19740
rect 11422 19728 11428 19780
rect 11480 19768 11486 19780
rect 13817 19771 13875 19777
rect 13817 19768 13829 19771
rect 11480 19740 13829 19768
rect 11480 19728 11486 19740
rect 13817 19737 13829 19740
rect 13863 19768 13875 19771
rect 14737 19771 14795 19777
rect 14737 19768 14749 19771
rect 13863 19740 14749 19768
rect 13863 19737 13875 19740
rect 13817 19731 13875 19737
rect 14737 19737 14749 19740
rect 14783 19768 14795 19771
rect 17310 19768 17316 19780
rect 14783 19740 17316 19768
rect 14783 19737 14795 19740
rect 14737 19731 14795 19737
rect 17310 19728 17316 19740
rect 17368 19728 17374 19780
rect 17957 19771 18015 19777
rect 17957 19737 17969 19771
rect 18003 19768 18015 19771
rect 18782 19768 18788 19780
rect 18003 19740 18788 19768
rect 18003 19737 18015 19740
rect 17957 19731 18015 19737
rect 18782 19728 18788 19740
rect 18840 19728 18846 19780
rect 22189 19771 22247 19777
rect 22189 19737 22201 19771
rect 22235 19768 22247 19771
rect 23842 19768 23848 19780
rect 22235 19740 23848 19768
rect 22235 19737 22247 19740
rect 22189 19731 22247 19737
rect 23842 19728 23848 19740
rect 23900 19728 23906 19780
rect 9088 19672 9536 19700
rect 12161 19703 12219 19709
rect 9088 19660 9094 19672
rect 12161 19669 12173 19703
rect 12207 19700 12219 19703
rect 13722 19700 13728 19712
rect 12207 19672 13728 19700
rect 12207 19669 12219 19672
rect 12161 19663 12219 19669
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 18506 19660 18512 19712
rect 18564 19660 18570 19712
rect 19334 19660 19340 19712
rect 19392 19660 19398 19712
rect 19426 19660 19432 19712
rect 19484 19700 19490 19712
rect 21542 19700 21548 19712
rect 19484 19672 21548 19700
rect 19484 19660 19490 19672
rect 21542 19660 21548 19672
rect 21600 19660 21606 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 1486 19456 1492 19508
rect 1544 19496 1550 19508
rect 2041 19499 2099 19505
rect 2041 19496 2053 19499
rect 1544 19468 2053 19496
rect 1544 19456 1550 19468
rect 2041 19465 2053 19468
rect 2087 19465 2099 19499
rect 2041 19459 2099 19465
rect 4154 19456 4160 19508
rect 4212 19496 4218 19508
rect 4249 19499 4307 19505
rect 4249 19496 4261 19499
rect 4212 19468 4261 19496
rect 4212 19456 4218 19468
rect 4249 19465 4261 19468
rect 4295 19465 4307 19499
rect 4249 19459 4307 19465
rect 7834 19456 7840 19508
rect 7892 19496 7898 19508
rect 8757 19499 8815 19505
rect 8757 19496 8769 19499
rect 7892 19468 8769 19496
rect 7892 19456 7898 19468
rect 8757 19465 8769 19468
rect 8803 19465 8815 19499
rect 8757 19459 8815 19465
rect 9217 19499 9275 19505
rect 9217 19465 9229 19499
rect 9263 19496 9275 19499
rect 9398 19496 9404 19508
rect 9263 19468 9404 19496
rect 9263 19465 9275 19468
rect 9217 19459 9275 19465
rect 9398 19456 9404 19468
rect 9456 19456 9462 19508
rect 11606 19456 11612 19508
rect 11664 19496 11670 19508
rect 11701 19499 11759 19505
rect 11701 19496 11713 19499
rect 11664 19468 11713 19496
rect 11664 19456 11670 19468
rect 11701 19465 11713 19468
rect 11747 19465 11759 19499
rect 11701 19459 11759 19465
rect 13909 19499 13967 19505
rect 13909 19465 13921 19499
rect 13955 19465 13967 19499
rect 13909 19459 13967 19465
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19496 16911 19499
rect 17218 19496 17224 19508
rect 16899 19468 17224 19496
rect 16899 19465 16911 19468
rect 16853 19459 16911 19465
rect 7098 19388 7104 19440
rect 7156 19428 7162 19440
rect 13924 19428 13952 19459
rect 17218 19456 17224 19468
rect 17276 19456 17282 19508
rect 17310 19456 17316 19508
rect 17368 19496 17374 19508
rect 17865 19499 17923 19505
rect 17865 19496 17877 19499
rect 17368 19468 17877 19496
rect 17368 19456 17374 19468
rect 17865 19465 17877 19468
rect 17911 19465 17923 19499
rect 17865 19459 17923 19465
rect 19426 19456 19432 19508
rect 19484 19456 19490 19508
rect 19518 19456 19524 19508
rect 19576 19496 19582 19508
rect 19797 19499 19855 19505
rect 19797 19496 19809 19499
rect 19576 19468 19809 19496
rect 19576 19456 19582 19468
rect 19797 19465 19809 19468
rect 19843 19465 19855 19499
rect 19797 19459 19855 19465
rect 19889 19499 19947 19505
rect 19889 19465 19901 19499
rect 19935 19496 19947 19499
rect 20806 19496 20812 19508
rect 19935 19468 20812 19496
rect 19935 19465 19947 19468
rect 19889 19459 19947 19465
rect 20806 19456 20812 19468
rect 20864 19456 20870 19508
rect 21174 19456 21180 19508
rect 21232 19456 21238 19508
rect 21818 19456 21824 19508
rect 21876 19496 21882 19508
rect 23753 19499 23811 19505
rect 23753 19496 23765 19499
rect 21876 19468 23765 19496
rect 21876 19456 21882 19468
rect 23753 19465 23765 19468
rect 23799 19465 23811 19499
rect 23753 19459 23811 19465
rect 14918 19428 14924 19440
rect 7156 19400 7314 19428
rect 13924 19400 14924 19428
rect 7156 19388 7162 19400
rect 14918 19388 14924 19400
rect 14976 19388 14982 19440
rect 18785 19431 18843 19437
rect 18785 19397 18797 19431
rect 18831 19428 18843 19431
rect 19242 19428 19248 19440
rect 18831 19400 19248 19428
rect 18831 19397 18843 19400
rect 18785 19391 18843 19397
rect 19242 19388 19248 19400
rect 19300 19388 19306 19440
rect 20530 19428 20536 19440
rect 19720 19400 20536 19428
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19360 2283 19363
rect 3602 19360 3608 19372
rect 2271 19332 3608 19360
rect 2271 19329 2283 19332
rect 2225 19323 2283 19329
rect 3602 19320 3608 19332
rect 3660 19320 3666 19372
rect 4433 19363 4491 19369
rect 4433 19329 4445 19363
rect 4479 19360 4491 19363
rect 6270 19360 6276 19372
rect 4479 19332 6276 19360
rect 4479 19329 4491 19332
rect 4433 19323 4491 19329
rect 6270 19320 6276 19332
rect 6328 19320 6334 19372
rect 6546 19320 6552 19372
rect 6604 19320 6610 19372
rect 8386 19320 8392 19372
rect 8444 19360 8450 19372
rect 8570 19360 8576 19372
rect 8444 19332 8576 19360
rect 8444 19320 8450 19332
rect 8570 19320 8576 19332
rect 8628 19360 8634 19372
rect 9125 19363 9183 19369
rect 9125 19360 9137 19363
rect 8628 19332 9137 19360
rect 8628 19320 8634 19332
rect 9125 19329 9137 19332
rect 9171 19329 9183 19363
rect 9125 19323 9183 19329
rect 12069 19363 12127 19369
rect 12069 19329 12081 19363
rect 12115 19360 12127 19363
rect 13354 19360 13360 19372
rect 12115 19332 13360 19360
rect 12115 19329 12127 19332
rect 12069 19323 12127 19329
rect 13354 19320 13360 19332
rect 13412 19320 13418 19372
rect 13538 19334 13544 19372
rect 13464 19320 13544 19334
rect 13596 19360 13602 19372
rect 14001 19364 14059 19369
rect 13924 19363 14059 19364
rect 13596 19320 13676 19360
rect 13464 19306 13676 19320
rect 13924 19336 14013 19363
rect 6822 19252 6828 19304
rect 6880 19252 6886 19304
rect 9214 19252 9220 19304
rect 9272 19292 9278 19304
rect 9309 19295 9367 19301
rect 9309 19292 9321 19295
rect 9272 19264 9321 19292
rect 9272 19252 9278 19264
rect 9309 19261 9321 19264
rect 9355 19261 9367 19295
rect 11054 19292 11060 19304
rect 9309 19255 9367 19261
rect 10888 19264 11060 19292
rect 10888 19168 10916 19264
rect 11054 19252 11060 19264
rect 11112 19292 11118 19304
rect 12161 19295 12219 19301
rect 12161 19292 12173 19295
rect 11112 19264 12173 19292
rect 11112 19252 11118 19264
rect 12161 19261 12173 19264
rect 12207 19261 12219 19295
rect 12161 19255 12219 19261
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19292 12311 19295
rect 12986 19292 12992 19304
rect 12299 19264 12992 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12268 19224 12296 19255
rect 12986 19252 12992 19264
rect 13044 19292 13050 19304
rect 13464 19292 13492 19306
rect 13924 19292 13952 19336
rect 14001 19329 14013 19336
rect 14047 19360 14059 19363
rect 14090 19360 14096 19372
rect 14047 19332 14096 19360
rect 14047 19329 14059 19332
rect 14001 19323 14059 19329
rect 14090 19320 14096 19332
rect 14148 19360 14154 19372
rect 14734 19360 14740 19372
rect 14148 19332 14740 19360
rect 14148 19320 14154 19332
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 17034 19320 17040 19372
rect 17092 19320 17098 19372
rect 19720 19360 19748 19400
rect 20530 19388 20536 19400
rect 20588 19388 20594 19440
rect 22554 19388 22560 19440
rect 22612 19428 22618 19440
rect 22612 19400 22770 19428
rect 22612 19388 22618 19400
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 17512 19332 19748 19360
rect 19904 19332 21097 19360
rect 14182 19292 14188 19304
rect 13044 19264 13492 19292
rect 13832 19264 13952 19292
rect 14016 19264 14188 19292
rect 13044 19252 13050 19264
rect 13078 19224 13084 19236
rect 11072 19196 12296 19224
rect 12360 19196 13084 19224
rect 11072 19168 11100 19196
rect 7558 19116 7564 19168
rect 7616 19156 7622 19168
rect 8297 19159 8355 19165
rect 8297 19156 8309 19159
rect 7616 19128 8309 19156
rect 7616 19116 7622 19128
rect 8297 19125 8309 19128
rect 8343 19125 8355 19159
rect 8297 19119 8355 19125
rect 10870 19116 10876 19168
rect 10928 19116 10934 19168
rect 11054 19116 11060 19168
rect 11112 19116 11118 19168
rect 11146 19116 11152 19168
rect 11204 19156 11210 19168
rect 11241 19159 11299 19165
rect 11241 19156 11253 19159
rect 11204 19128 11253 19156
rect 11204 19116 11210 19128
rect 11241 19125 11253 19128
rect 11287 19156 11299 19159
rect 11330 19156 11336 19168
rect 11287 19128 11336 19156
rect 11287 19125 11299 19128
rect 11241 19119 11299 19125
rect 11330 19116 11336 19128
rect 11388 19116 11394 19168
rect 11698 19116 11704 19168
rect 11756 19156 11762 19168
rect 12360 19156 12388 19196
rect 13078 19184 13084 19196
rect 13136 19184 13142 19236
rect 13262 19184 13268 19236
rect 13320 19224 13326 19236
rect 13541 19227 13599 19233
rect 13541 19224 13553 19227
rect 13320 19196 13553 19224
rect 13320 19184 13326 19196
rect 13541 19193 13553 19196
rect 13587 19193 13599 19227
rect 13541 19187 13599 19193
rect 11756 19128 12388 19156
rect 11756 19116 11762 19128
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 13173 19159 13231 19165
rect 13173 19156 13185 19159
rect 12492 19128 13185 19156
rect 12492 19116 12498 19128
rect 13173 19125 13185 19128
rect 13219 19156 13231 19159
rect 13832 19156 13860 19264
rect 14016 19236 14044 19264
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 14550 19252 14556 19304
rect 14608 19252 14614 19304
rect 13998 19184 14004 19236
rect 14056 19184 14062 19236
rect 17512 19233 17540 19332
rect 17957 19295 18015 19301
rect 17957 19292 17969 19295
rect 17788 19264 17969 19292
rect 17497 19227 17555 19233
rect 17497 19193 17509 19227
rect 17543 19193 17555 19227
rect 17497 19187 17555 19193
rect 17788 19168 17816 19264
rect 17957 19261 17969 19264
rect 18003 19261 18015 19295
rect 17957 19255 18015 19261
rect 18141 19295 18199 19301
rect 18141 19261 18153 19295
rect 18187 19292 18199 19295
rect 19334 19292 19340 19304
rect 18187 19264 19340 19292
rect 18187 19261 18199 19264
rect 18141 19255 18199 19261
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 19242 19184 19248 19236
rect 19300 19224 19306 19236
rect 19904 19224 19932 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 20073 19295 20131 19301
rect 20073 19261 20085 19295
rect 20119 19292 20131 19295
rect 21266 19292 21272 19304
rect 20119 19264 21272 19292
rect 20119 19261 20131 19264
rect 20073 19255 20131 19261
rect 21266 19252 21272 19264
rect 21324 19252 21330 19304
rect 21361 19295 21419 19301
rect 21361 19261 21373 19295
rect 21407 19292 21419 19295
rect 21818 19292 21824 19304
rect 21407 19264 21824 19292
rect 21407 19261 21419 19264
rect 21361 19255 21419 19261
rect 21818 19252 21824 19264
rect 21876 19252 21882 19304
rect 22002 19252 22008 19304
rect 22060 19252 22066 19304
rect 22281 19295 22339 19301
rect 22281 19261 22293 19295
rect 22327 19292 22339 19295
rect 22738 19292 22744 19304
rect 22327 19264 22744 19292
rect 22327 19261 22339 19264
rect 22281 19255 22339 19261
rect 22738 19252 22744 19264
rect 22796 19252 22802 19304
rect 19300 19196 19932 19224
rect 19300 19184 19306 19196
rect 13219 19128 13860 19156
rect 13219 19125 13231 19128
rect 13173 19119 13231 19125
rect 17126 19116 17132 19168
rect 17184 19156 17190 19168
rect 17770 19156 17776 19168
rect 17184 19128 17776 19156
rect 17184 19116 17190 19128
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 18874 19116 18880 19168
rect 18932 19116 18938 19168
rect 20714 19116 20720 19168
rect 20772 19116 20778 19168
rect 22646 19116 22652 19168
rect 22704 19156 22710 19168
rect 24029 19159 24087 19165
rect 24029 19156 24041 19159
rect 22704 19128 24041 19156
rect 22704 19116 22710 19128
rect 24029 19125 24041 19128
rect 24075 19156 24087 19159
rect 24394 19156 24400 19168
rect 24075 19128 24400 19156
rect 24075 19125 24087 19128
rect 24029 19119 24087 19125
rect 24394 19116 24400 19128
rect 24452 19116 24458 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 8389 18955 8447 18961
rect 8389 18952 8401 18955
rect 8352 18924 8401 18952
rect 8352 18912 8358 18924
rect 8389 18921 8401 18924
rect 8435 18952 8447 18955
rect 11146 18952 11152 18964
rect 8435 18924 11152 18952
rect 8435 18921 8447 18924
rect 8389 18915 8447 18921
rect 11146 18912 11152 18924
rect 11204 18912 11210 18964
rect 12158 18912 12164 18964
rect 12216 18912 12222 18964
rect 13722 18912 13728 18964
rect 13780 18952 13786 18964
rect 14277 18955 14335 18961
rect 14277 18952 14289 18955
rect 13780 18924 14289 18952
rect 13780 18912 13786 18924
rect 14277 18921 14289 18924
rect 14323 18921 14335 18955
rect 14277 18915 14335 18921
rect 15764 18924 17540 18952
rect 1302 18776 1308 18828
rect 1360 18816 1366 18828
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 1360 18788 2053 18816
rect 1360 18776 1366 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 1762 18708 1768 18760
rect 1820 18708 1826 18760
rect 6546 18708 6552 18760
rect 6604 18748 6610 18760
rect 9306 18748 9312 18760
rect 6604 18720 9312 18748
rect 6604 18708 6610 18720
rect 9306 18708 9312 18720
rect 9364 18748 9370 18760
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 9364 18720 9781 18748
rect 9364 18708 9370 18720
rect 9769 18717 9781 18720
rect 9815 18717 9827 18751
rect 11164 18748 11192 18912
rect 12710 18844 12716 18896
rect 12768 18884 12774 18896
rect 12768 18856 13584 18884
rect 12768 18844 12774 18856
rect 13446 18776 13452 18828
rect 13504 18776 13510 18828
rect 13556 18825 13584 18856
rect 13814 18844 13820 18896
rect 13872 18884 13878 18896
rect 13998 18884 14004 18896
rect 13872 18856 14004 18884
rect 13872 18844 13878 18856
rect 13998 18844 14004 18856
rect 14056 18844 14062 18896
rect 13541 18819 13599 18825
rect 13541 18785 13553 18819
rect 13587 18816 13599 18819
rect 14182 18816 14188 18828
rect 13587 18788 14188 18816
rect 13587 18785 13599 18788
rect 13541 18779 13599 18785
rect 14182 18776 14188 18788
rect 14240 18776 14246 18828
rect 14550 18776 14556 18828
rect 14608 18816 14614 18828
rect 14826 18816 14832 18828
rect 14608 18788 14832 18816
rect 14608 18776 14614 18788
rect 14826 18776 14832 18788
rect 14884 18776 14890 18828
rect 11885 18751 11943 18757
rect 11885 18748 11897 18751
rect 11164 18734 11897 18748
rect 11178 18720 11897 18734
rect 9769 18711 9827 18717
rect 11885 18717 11897 18720
rect 11931 18748 11943 18751
rect 14645 18751 14703 18757
rect 11931 18720 12434 18748
rect 11931 18717 11943 18720
rect 11885 18711 11943 18717
rect 10045 18683 10103 18689
rect 10045 18649 10057 18683
rect 10091 18649 10103 18683
rect 12250 18680 12256 18692
rect 10045 18643 10103 18649
rect 11808 18652 12256 18680
rect 8570 18572 8576 18624
rect 8628 18572 8634 18624
rect 9122 18572 9128 18624
rect 9180 18612 9186 18624
rect 9401 18615 9459 18621
rect 9401 18612 9413 18615
rect 9180 18584 9413 18612
rect 9180 18572 9186 18584
rect 9401 18581 9413 18584
rect 9447 18612 9459 18615
rect 10060 18612 10088 18643
rect 11808 18624 11836 18652
rect 12250 18640 12256 18652
rect 12308 18640 12314 18692
rect 12406 18680 12434 18720
rect 14645 18717 14657 18751
rect 14691 18748 14703 18751
rect 15764 18748 15792 18924
rect 17512 18884 17540 18924
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 18325 18955 18383 18961
rect 18325 18952 18337 18955
rect 17828 18924 18337 18952
rect 17828 18912 17834 18924
rect 18325 18921 18337 18924
rect 18371 18921 18383 18955
rect 18325 18915 18383 18921
rect 18966 18912 18972 18964
rect 19024 18912 19030 18964
rect 22738 18912 22744 18964
rect 22796 18952 22802 18964
rect 24029 18955 24087 18961
rect 24029 18952 24041 18955
rect 22796 18924 24041 18952
rect 22796 18912 22802 18924
rect 24029 18921 24041 18924
rect 24075 18921 24087 18955
rect 24029 18915 24087 18921
rect 24394 18912 24400 18964
rect 24452 18912 24458 18964
rect 18506 18884 18512 18896
rect 17512 18856 18512 18884
rect 18506 18844 18512 18856
rect 18564 18844 18570 18896
rect 18601 18887 18659 18893
rect 18601 18853 18613 18887
rect 18647 18884 18659 18887
rect 20622 18884 20628 18896
rect 18647 18856 20628 18884
rect 18647 18853 18659 18856
rect 18601 18847 18659 18853
rect 15838 18776 15844 18828
rect 15896 18816 15902 18828
rect 17957 18819 18015 18825
rect 17957 18816 17969 18819
rect 15896 18788 17969 18816
rect 15896 18776 15902 18788
rect 17957 18785 17969 18788
rect 18003 18785 18015 18819
rect 17957 18779 18015 18785
rect 14691 18720 15792 18748
rect 14691 18717 14703 18720
rect 14645 18711 14703 18717
rect 16206 18708 16212 18760
rect 16264 18708 16270 18760
rect 18616 18748 18644 18847
rect 20622 18844 20628 18856
rect 20680 18844 20686 18896
rect 17618 18720 18644 18748
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19024 18720 19625 18748
rect 19024 18708 19030 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18748 20407 18751
rect 20438 18748 20444 18760
rect 20395 18720 20444 18748
rect 20395 18717 20407 18720
rect 20349 18711 20407 18717
rect 20438 18708 20444 18720
rect 20496 18748 20502 18760
rect 21545 18751 21603 18757
rect 21545 18748 21557 18751
rect 20496 18720 21557 18748
rect 20496 18708 20502 18720
rect 21545 18717 21557 18720
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 22281 18751 22339 18757
rect 22281 18717 22293 18751
rect 22327 18717 22339 18751
rect 22281 18711 22339 18717
rect 12802 18680 12808 18692
rect 12406 18652 12808 18680
rect 12802 18640 12808 18652
rect 12860 18640 12866 18692
rect 13722 18640 13728 18692
rect 13780 18680 13786 18692
rect 14737 18683 14795 18689
rect 14737 18680 14749 18683
rect 13780 18652 14749 18680
rect 13780 18640 13786 18652
rect 14737 18649 14749 18652
rect 14783 18649 14795 18683
rect 14737 18643 14795 18649
rect 16485 18683 16543 18689
rect 16485 18649 16497 18683
rect 16531 18649 16543 18683
rect 16485 18643 16543 18649
rect 21177 18683 21235 18689
rect 21177 18649 21189 18683
rect 21223 18680 21235 18683
rect 21726 18680 21732 18692
rect 21223 18652 21732 18680
rect 21223 18649 21235 18652
rect 21177 18643 21235 18649
rect 11054 18612 11060 18624
rect 9447 18584 11060 18612
rect 9447 18581 9459 18584
rect 9401 18575 9459 18581
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 11517 18615 11575 18621
rect 11517 18581 11529 18615
rect 11563 18612 11575 18615
rect 11790 18612 11796 18624
rect 11563 18584 11796 18612
rect 11563 18581 11575 18584
rect 11517 18575 11575 18581
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 11974 18572 11980 18624
rect 12032 18612 12038 18624
rect 12989 18615 13047 18621
rect 12989 18612 13001 18615
rect 12032 18584 13001 18612
rect 12032 18572 12038 18584
rect 12989 18581 13001 18584
rect 13035 18581 13047 18615
rect 12989 18575 13047 18581
rect 13354 18572 13360 18624
rect 13412 18572 13418 18624
rect 16500 18612 16528 18643
rect 21726 18640 21732 18652
rect 21784 18680 21790 18692
rect 22002 18680 22008 18692
rect 21784 18652 22008 18680
rect 21784 18640 21790 18652
rect 22002 18640 22008 18652
rect 22060 18680 22066 18692
rect 22296 18680 22324 18711
rect 22060 18652 22324 18680
rect 22060 18640 22066 18652
rect 22554 18640 22560 18692
rect 22612 18640 22618 18692
rect 22646 18640 22652 18692
rect 22704 18680 22710 18692
rect 22704 18652 23046 18680
rect 22704 18640 22710 18652
rect 18966 18612 18972 18624
rect 16500 18584 18972 18612
rect 18966 18572 18972 18584
rect 19024 18572 19030 18624
rect 19702 18572 19708 18624
rect 19760 18572 19766 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 7745 18411 7803 18417
rect 7745 18408 7757 18411
rect 7524 18380 7757 18408
rect 7524 18368 7530 18380
rect 7745 18377 7757 18380
rect 7791 18377 7803 18411
rect 7745 18371 7803 18377
rect 10410 18368 10416 18420
rect 10468 18368 10474 18420
rect 10781 18411 10839 18417
rect 10781 18377 10793 18411
rect 10827 18408 10839 18411
rect 12158 18408 12164 18420
rect 10827 18380 12164 18408
rect 10827 18377 10839 18380
rect 10781 18371 10839 18377
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 13354 18368 13360 18420
rect 13412 18408 13418 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 13412 18380 14289 18408
rect 13412 18368 13418 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 14645 18411 14703 18417
rect 14645 18377 14657 18411
rect 14691 18408 14703 18411
rect 15381 18411 15439 18417
rect 15381 18408 15393 18411
rect 14691 18380 15393 18408
rect 14691 18377 14703 18380
rect 14645 18371 14703 18377
rect 15381 18377 15393 18380
rect 15427 18408 15439 18411
rect 18322 18408 18328 18420
rect 15427 18380 18328 18408
rect 15427 18377 15439 18380
rect 15381 18371 15439 18377
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 19334 18408 19340 18420
rect 19168 18380 19340 18408
rect 9306 18300 9312 18352
rect 9364 18300 9370 18352
rect 11698 18300 11704 18352
rect 11756 18340 11762 18352
rect 12069 18343 12127 18349
rect 12069 18340 12081 18343
rect 11756 18312 12081 18340
rect 11756 18300 11762 18312
rect 12069 18309 12081 18312
rect 12115 18309 12127 18343
rect 12069 18303 12127 18309
rect 13722 18300 13728 18352
rect 13780 18340 13786 18352
rect 13909 18343 13967 18349
rect 13909 18340 13921 18343
rect 13780 18312 13921 18340
rect 13780 18300 13786 18312
rect 13909 18309 13921 18312
rect 13955 18309 13967 18343
rect 13909 18303 13967 18309
rect 16298 18300 16304 18352
rect 16356 18340 16362 18352
rect 16482 18340 16488 18352
rect 16356 18312 16488 18340
rect 16356 18300 16362 18312
rect 16482 18300 16488 18312
rect 16540 18300 16546 18352
rect 17221 18343 17279 18349
rect 17221 18309 17233 18343
rect 17267 18340 17279 18343
rect 17494 18340 17500 18352
rect 17267 18312 17500 18340
rect 17267 18309 17279 18312
rect 17221 18303 17279 18309
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 19168 18349 19196 18380
rect 19334 18368 19340 18380
rect 19392 18368 19398 18420
rect 19153 18343 19211 18349
rect 19153 18309 19165 18343
rect 19199 18309 19211 18343
rect 20622 18340 20628 18352
rect 20378 18312 20628 18340
rect 19153 18303 19211 18309
rect 20622 18300 20628 18312
rect 20680 18300 20686 18352
rect 7653 18275 7711 18281
rect 7653 18272 7665 18275
rect 6932 18244 7665 18272
rect 4890 18096 4896 18148
rect 4948 18136 4954 18148
rect 6932 18145 6960 18244
rect 7653 18241 7665 18244
rect 7699 18241 7711 18275
rect 7653 18235 7711 18241
rect 8481 18275 8539 18281
rect 8481 18241 8493 18275
rect 8527 18272 8539 18275
rect 9766 18272 9772 18284
rect 8527 18244 9772 18272
rect 8527 18241 8539 18244
rect 8481 18235 8539 18241
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 10318 18232 10324 18284
rect 10376 18272 10382 18284
rect 10376 18244 11100 18272
rect 10376 18232 10382 18244
rect 11072 18216 11100 18244
rect 11882 18232 11888 18284
rect 11940 18272 11946 18284
rect 11940 18244 12296 18272
rect 11940 18232 11946 18244
rect 7558 18164 7564 18216
rect 7616 18204 7622 18216
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 7616 18176 7849 18204
rect 7616 18164 7622 18176
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 10873 18207 10931 18213
rect 10873 18173 10885 18207
rect 10919 18173 10931 18207
rect 10873 18167 10931 18173
rect 6917 18139 6975 18145
rect 6917 18136 6929 18139
rect 4948 18108 6929 18136
rect 4948 18096 4954 18108
rect 6917 18105 6929 18108
rect 6963 18105 6975 18139
rect 6917 18099 6975 18105
rect 4154 18028 4160 18080
rect 4212 18068 4218 18080
rect 5534 18068 5540 18080
rect 4212 18040 5540 18068
rect 4212 18028 4218 18040
rect 5534 18028 5540 18040
rect 5592 18028 5598 18080
rect 7285 18071 7343 18077
rect 7285 18037 7297 18071
rect 7331 18068 7343 18071
rect 8662 18068 8668 18080
rect 7331 18040 8668 18068
rect 7331 18037 7343 18040
rect 7285 18031 7343 18037
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 9766 18028 9772 18080
rect 9824 18028 9830 18080
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 10045 18071 10103 18077
rect 10045 18068 10057 18071
rect 9916 18040 10057 18068
rect 9916 18028 9922 18040
rect 10045 18037 10057 18040
rect 10091 18068 10103 18071
rect 10888 18068 10916 18167
rect 11054 18164 11060 18216
rect 11112 18164 11118 18216
rect 12158 18164 12164 18216
rect 12216 18164 12222 18216
rect 12268 18213 12296 18244
rect 12253 18207 12311 18213
rect 12253 18173 12265 18207
rect 12299 18173 12311 18207
rect 12253 18167 12311 18173
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 13541 18207 13599 18213
rect 13541 18204 13553 18207
rect 12492 18176 13553 18204
rect 12492 18164 12498 18176
rect 13541 18173 13553 18176
rect 13587 18173 13599 18207
rect 13541 18167 13599 18173
rect 11514 18096 11520 18148
rect 11572 18136 11578 18148
rect 11701 18139 11759 18145
rect 11701 18136 11713 18139
rect 11572 18108 11713 18136
rect 11572 18096 11578 18108
rect 11701 18105 11713 18108
rect 11747 18105 11759 18139
rect 11701 18099 11759 18105
rect 12342 18096 12348 18148
rect 12400 18136 12406 18148
rect 13740 18136 13768 18300
rect 14737 18275 14795 18281
rect 14737 18241 14749 18275
rect 14783 18272 14795 18275
rect 15010 18272 15016 18284
rect 14783 18244 15016 18272
rect 14783 18241 14795 18244
rect 14737 18235 14795 18241
rect 13817 18207 13875 18213
rect 13817 18173 13829 18207
rect 13863 18204 13875 18207
rect 14752 18204 14780 18235
rect 15010 18232 15016 18244
rect 15068 18232 15074 18284
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 14921 18207 14979 18213
rect 14921 18204 14933 18207
rect 13863 18176 14780 18204
rect 14844 18176 14933 18204
rect 13863 18173 13875 18176
rect 13817 18167 13875 18173
rect 12400 18108 13768 18136
rect 12400 18096 12406 18108
rect 10091 18040 10916 18068
rect 10091 18037 10103 18040
rect 10045 18031 10103 18037
rect 12618 18028 12624 18080
rect 12676 18068 12682 18080
rect 13262 18068 13268 18080
rect 12676 18040 13268 18068
rect 12676 18028 12682 18040
rect 13262 18028 13268 18040
rect 13320 18068 13326 18080
rect 14844 18068 14872 18176
rect 14921 18173 14933 18176
rect 14967 18204 14979 18207
rect 15286 18204 15292 18216
rect 14967 18176 15292 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 15286 18164 15292 18176
rect 15344 18204 15350 18216
rect 15930 18204 15936 18216
rect 15344 18176 15936 18204
rect 15344 18164 15350 18176
rect 15930 18164 15936 18176
rect 15988 18164 15994 18216
rect 16206 18164 16212 18216
rect 16264 18204 16270 18216
rect 16482 18204 16488 18216
rect 16264 18176 16488 18204
rect 16264 18164 16270 18176
rect 16482 18164 16488 18176
rect 16540 18204 16546 18216
rect 18325 18207 18383 18213
rect 18325 18204 18337 18207
rect 16540 18176 18337 18204
rect 16540 18164 16546 18176
rect 18325 18173 18337 18176
rect 18371 18204 18383 18207
rect 18877 18207 18935 18213
rect 18877 18204 18889 18207
rect 18371 18176 18889 18204
rect 18371 18173 18383 18176
rect 18325 18167 18383 18173
rect 18877 18173 18889 18176
rect 18923 18173 18935 18207
rect 18877 18167 18935 18173
rect 19150 18164 19156 18216
rect 19208 18204 19214 18216
rect 21284 18204 21312 18235
rect 22094 18232 22100 18284
rect 22152 18232 22158 18284
rect 24026 18232 24032 18284
rect 24084 18232 24090 18284
rect 19208 18176 21312 18204
rect 23293 18207 23351 18213
rect 19208 18164 19214 18176
rect 23293 18173 23305 18207
rect 23339 18204 23351 18207
rect 23382 18204 23388 18216
rect 23339 18176 23388 18204
rect 23339 18173 23351 18176
rect 23293 18167 23351 18173
rect 23382 18164 23388 18176
rect 23440 18164 23446 18216
rect 24762 18164 24768 18216
rect 24820 18164 24826 18216
rect 21453 18139 21511 18145
rect 21453 18105 21465 18139
rect 21499 18136 21511 18139
rect 22186 18136 22192 18148
rect 21499 18108 22192 18136
rect 21499 18105 21511 18108
rect 21453 18099 21511 18105
rect 22186 18096 22192 18108
rect 22244 18096 22250 18148
rect 13320 18040 14872 18068
rect 13320 18028 13326 18040
rect 14918 18028 14924 18080
rect 14976 18068 14982 18080
rect 18874 18068 18880 18080
rect 14976 18040 18880 18068
rect 14976 18028 14982 18040
rect 18874 18028 18880 18040
rect 18932 18028 18938 18080
rect 20162 18028 20168 18080
rect 20220 18068 20226 18080
rect 20625 18071 20683 18077
rect 20625 18068 20637 18071
rect 20220 18040 20637 18068
rect 20220 18028 20226 18040
rect 20625 18037 20637 18040
rect 20671 18037 20683 18071
rect 20625 18031 20683 18037
rect 22094 18028 22100 18080
rect 22152 18068 22158 18080
rect 22738 18068 22744 18080
rect 22152 18040 22744 18068
rect 22152 18028 22158 18040
rect 22738 18028 22744 18040
rect 22796 18028 22802 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 6270 17824 6276 17876
rect 6328 17824 6334 17876
rect 7282 17824 7288 17876
rect 7340 17864 7346 17876
rect 9125 17867 9183 17873
rect 9125 17864 9137 17867
rect 7340 17836 9137 17864
rect 7340 17824 7346 17836
rect 9125 17833 9137 17836
rect 9171 17833 9183 17867
rect 17494 17864 17500 17876
rect 9125 17827 9183 17833
rect 12636 17836 17500 17864
rect 8294 17756 8300 17808
rect 8352 17796 8358 17808
rect 8665 17799 8723 17805
rect 8665 17796 8677 17799
rect 8352 17768 8677 17796
rect 8352 17756 8358 17768
rect 8665 17765 8677 17768
rect 8711 17765 8723 17799
rect 8665 17759 8723 17765
rect 6825 17731 6883 17737
rect 6825 17697 6837 17731
rect 6871 17728 6883 17731
rect 6914 17728 6920 17740
rect 6871 17700 6920 17728
rect 6871 17697 6883 17700
rect 6825 17691 6883 17697
rect 6914 17688 6920 17700
rect 6972 17688 6978 17740
rect 7834 17688 7840 17740
rect 7892 17728 7898 17740
rect 7929 17731 7987 17737
rect 7929 17728 7941 17731
rect 7892 17700 7941 17728
rect 7892 17688 7898 17700
rect 7929 17697 7941 17700
rect 7975 17697 7987 17731
rect 7929 17691 7987 17697
rect 8113 17731 8171 17737
rect 8113 17697 8125 17731
rect 8159 17728 8171 17731
rect 8386 17728 8392 17740
rect 8159 17700 8392 17728
rect 8159 17697 8171 17700
rect 8113 17691 8171 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9456 17700 9689 17728
rect 9456 17688 9462 17700
rect 9677 17697 9689 17700
rect 9723 17697 9735 17731
rect 9677 17691 9735 17697
rect 9766 17688 9772 17740
rect 9824 17728 9830 17740
rect 12437 17731 12495 17737
rect 12437 17728 12449 17731
rect 9824 17700 12449 17728
rect 9824 17688 9830 17700
rect 10520 17669 10548 17700
rect 12437 17697 12449 17700
rect 12483 17728 12495 17731
rect 12636 17728 12664 17836
rect 17494 17824 17500 17836
rect 17552 17824 17558 17876
rect 21266 17824 21272 17876
rect 21324 17864 21330 17876
rect 21637 17867 21695 17873
rect 21637 17864 21649 17867
rect 21324 17836 21649 17864
rect 21324 17824 21330 17836
rect 21637 17833 21649 17836
rect 21683 17864 21695 17867
rect 21683 17836 22232 17864
rect 21683 17833 21695 17836
rect 21637 17827 21695 17833
rect 12710 17756 12716 17808
rect 12768 17756 12774 17808
rect 17221 17799 17279 17805
rect 17221 17796 17233 17799
rect 16684 17768 17233 17796
rect 12483 17700 12664 17728
rect 12728 17728 12756 17756
rect 13449 17731 13507 17737
rect 13449 17728 13461 17731
rect 12728 17700 13461 17728
rect 12483 17697 12495 17700
rect 12437 17691 12495 17697
rect 10505 17663 10563 17669
rect 10505 17629 10517 17663
rect 10551 17629 10563 17663
rect 10505 17623 10563 17629
rect 6641 17595 6699 17601
rect 6641 17561 6653 17595
rect 6687 17592 6699 17595
rect 6687 17564 7512 17592
rect 6687 17561 6699 17564
rect 6641 17555 6699 17561
rect 6733 17527 6791 17533
rect 6733 17493 6745 17527
rect 6779 17524 6791 17527
rect 7282 17524 7288 17536
rect 6779 17496 7288 17524
rect 6779 17493 6791 17496
rect 6733 17487 6791 17493
rect 7282 17484 7288 17496
rect 7340 17484 7346 17536
rect 7484 17533 7512 17564
rect 9306 17552 9312 17604
rect 9364 17592 9370 17604
rect 9364 17564 9720 17592
rect 9364 17552 9370 17564
rect 7469 17527 7527 17533
rect 7469 17493 7481 17527
rect 7515 17493 7527 17527
rect 7469 17487 7527 17493
rect 7834 17484 7840 17536
rect 7892 17484 7898 17536
rect 9490 17484 9496 17536
rect 9548 17484 9554 17536
rect 9582 17484 9588 17536
rect 9640 17484 9646 17536
rect 9692 17524 9720 17564
rect 11330 17552 11336 17604
rect 11388 17552 11394 17604
rect 11606 17552 11612 17604
rect 11664 17592 11670 17604
rect 12728 17592 12756 17700
rect 13449 17697 13461 17700
rect 13495 17697 13507 17731
rect 13449 17691 13507 17697
rect 13633 17731 13691 17737
rect 13633 17697 13645 17731
rect 13679 17728 13691 17731
rect 13998 17728 14004 17740
rect 13679 17700 14004 17728
rect 13679 17697 13691 17700
rect 13633 17691 13691 17697
rect 13998 17688 14004 17700
rect 14056 17728 14062 17740
rect 14274 17728 14280 17740
rect 14056 17700 14280 17728
rect 14056 17688 14062 17700
rect 14274 17688 14280 17700
rect 14332 17688 14338 17740
rect 14734 17688 14740 17740
rect 14792 17688 14798 17740
rect 14826 17688 14832 17740
rect 14884 17688 14890 17740
rect 16390 17688 16396 17740
rect 16448 17728 16454 17740
rect 16684 17737 16712 17768
rect 17221 17765 17233 17768
rect 17267 17765 17279 17799
rect 17221 17759 17279 17765
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 16448 17700 16681 17728
rect 16448 17688 16454 17700
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 16853 17731 16911 17737
rect 16853 17697 16865 17731
rect 16899 17728 16911 17731
rect 17126 17728 17132 17740
rect 16899 17700 17132 17728
rect 16899 17697 16911 17700
rect 16853 17691 16911 17697
rect 17126 17688 17132 17700
rect 17184 17688 17190 17740
rect 21726 17688 21732 17740
rect 21784 17728 21790 17740
rect 22097 17731 22155 17737
rect 22097 17728 22109 17731
rect 21784 17700 22109 17728
rect 21784 17688 21790 17700
rect 22097 17697 22109 17700
rect 22143 17697 22155 17731
rect 22204 17728 22232 17836
rect 22554 17824 22560 17876
rect 22612 17864 22618 17876
rect 22738 17864 22744 17876
rect 22612 17836 22744 17864
rect 22612 17824 22618 17836
rect 22738 17824 22744 17836
rect 22796 17864 22802 17876
rect 23845 17867 23903 17873
rect 23845 17864 23857 17867
rect 22796 17836 23857 17864
rect 22796 17824 22802 17836
rect 23845 17833 23857 17836
rect 23891 17833 23903 17867
rect 23845 17827 23903 17833
rect 22373 17731 22431 17737
rect 22373 17728 22385 17731
rect 22204 17700 22385 17728
rect 22097 17691 22155 17697
rect 22373 17697 22385 17700
rect 22419 17697 22431 17731
rect 22373 17691 22431 17697
rect 14645 17663 14703 17669
rect 14645 17629 14657 17663
rect 14691 17660 14703 17663
rect 14918 17660 14924 17672
rect 14691 17632 14924 17660
rect 14691 17629 14703 17632
rect 14645 17623 14703 17629
rect 14918 17620 14924 17632
rect 14976 17620 14982 17672
rect 15562 17620 15568 17672
rect 15620 17620 15626 17672
rect 19518 17620 19524 17672
rect 19576 17660 19582 17672
rect 19889 17663 19947 17669
rect 19889 17660 19901 17663
rect 19576 17632 19901 17660
rect 19576 17620 19582 17632
rect 19889 17629 19901 17632
rect 19935 17629 19947 17663
rect 19889 17623 19947 17629
rect 24854 17620 24860 17672
rect 24912 17620 24918 17672
rect 11664 17564 12756 17592
rect 13357 17595 13415 17601
rect 11664 17552 11670 17564
rect 13357 17561 13369 17595
rect 13403 17592 13415 17595
rect 15378 17592 15384 17604
rect 13403 17564 15384 17592
rect 13403 17561 13415 17564
rect 13357 17555 13415 17561
rect 15378 17552 15384 17564
rect 15436 17552 15442 17604
rect 18874 17592 18880 17604
rect 16224 17564 18880 17592
rect 11885 17527 11943 17533
rect 11885 17524 11897 17527
rect 9692 17496 11897 17524
rect 11885 17493 11897 17496
rect 11931 17493 11943 17527
rect 11885 17487 11943 17493
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 12989 17527 13047 17533
rect 12989 17524 13001 17527
rect 12768 17496 13001 17524
rect 12768 17484 12774 17496
rect 12989 17493 13001 17496
rect 13035 17493 13047 17527
rect 12989 17487 13047 17493
rect 14274 17484 14280 17536
rect 14332 17484 14338 17536
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 16224 17533 16252 17564
rect 18874 17552 18880 17564
rect 18932 17552 18938 17604
rect 20162 17552 20168 17604
rect 20220 17552 20226 17604
rect 20622 17552 20628 17604
rect 20680 17552 20686 17604
rect 22646 17552 22652 17604
rect 22704 17592 22710 17604
rect 22830 17592 22836 17604
rect 22704 17564 22836 17592
rect 22704 17552 22710 17564
rect 15657 17527 15715 17533
rect 15657 17524 15669 17527
rect 15620 17496 15669 17524
rect 15620 17484 15626 17496
rect 15657 17493 15669 17496
rect 15703 17493 15715 17527
rect 15657 17487 15715 17493
rect 16209 17527 16267 17533
rect 16209 17493 16221 17527
rect 16255 17493 16267 17527
rect 16209 17487 16267 17493
rect 16574 17484 16580 17536
rect 16632 17484 16638 17536
rect 22756 17524 22784 17564
rect 22830 17552 22836 17564
rect 22888 17552 22894 17604
rect 24121 17527 24179 17533
rect 24121 17524 24133 17527
rect 22756 17496 24133 17524
rect 24121 17493 24133 17496
rect 24167 17493 24179 17527
rect 24121 17487 24179 17493
rect 24302 17484 24308 17536
rect 24360 17524 24366 17536
rect 24673 17527 24731 17533
rect 24673 17524 24685 17527
rect 24360 17496 24685 17524
rect 24360 17484 24366 17496
rect 24673 17493 24685 17496
rect 24719 17493 24731 17527
rect 24673 17487 24731 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 4522 17280 4528 17332
rect 4580 17320 4586 17332
rect 4580 17292 9076 17320
rect 4580 17280 4586 17292
rect 8294 17252 8300 17264
rect 8050 17224 8300 17252
rect 8294 17212 8300 17224
rect 8352 17212 8358 17264
rect 9048 17196 9076 17292
rect 9490 17280 9496 17332
rect 9548 17320 9554 17332
rect 10045 17323 10103 17329
rect 10045 17320 10057 17323
rect 9548 17292 10057 17320
rect 9548 17280 9554 17292
rect 10045 17289 10057 17292
rect 10091 17289 10103 17323
rect 10045 17283 10103 17289
rect 10413 17323 10471 17329
rect 10413 17289 10425 17323
rect 10459 17320 10471 17323
rect 12066 17320 12072 17332
rect 10459 17292 12072 17320
rect 10459 17289 10471 17292
rect 10413 17283 10471 17289
rect 12066 17280 12072 17292
rect 12124 17280 12130 17332
rect 14182 17280 14188 17332
rect 14240 17320 14246 17332
rect 14369 17323 14427 17329
rect 14369 17320 14381 17323
rect 14240 17292 14381 17320
rect 14240 17280 14246 17292
rect 14369 17289 14381 17292
rect 14415 17289 14427 17323
rect 14369 17283 14427 17289
rect 14826 17280 14832 17332
rect 14884 17280 14890 17332
rect 19518 17320 19524 17332
rect 17788 17292 19524 17320
rect 12802 17212 12808 17264
rect 12860 17252 12866 17264
rect 13354 17252 13360 17264
rect 12860 17224 13360 17252
rect 12860 17212 12866 17224
rect 13354 17212 13360 17224
rect 13412 17212 13418 17264
rect 17788 17252 17816 17292
rect 19518 17280 19524 17292
rect 19576 17280 19582 17332
rect 17696 17224 17816 17252
rect 6546 17144 6552 17196
rect 6604 17144 6610 17196
rect 9030 17144 9036 17196
rect 9088 17144 9094 17196
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 17696 17193 17724 17224
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 18012 17224 18446 17252
rect 18012 17212 18018 17224
rect 21082 17212 21088 17264
rect 21140 17252 21146 17264
rect 22097 17255 22155 17261
rect 22097 17252 22109 17255
rect 21140 17224 22109 17252
rect 21140 17212 21146 17224
rect 22097 17221 22109 17224
rect 22143 17221 22155 17255
rect 22097 17215 22155 17221
rect 17037 17187 17095 17193
rect 17037 17184 17049 17187
rect 16724 17156 17049 17184
rect 16724 17144 16730 17156
rect 17037 17153 17049 17156
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 19797 17187 19855 17193
rect 19797 17153 19809 17187
rect 19843 17184 19855 17187
rect 20622 17184 20628 17196
rect 19843 17156 20628 17184
rect 19843 17153 19855 17156
rect 19797 17147 19855 17153
rect 20622 17144 20628 17156
rect 20680 17184 20686 17196
rect 20901 17187 20959 17193
rect 20901 17184 20913 17187
rect 20680 17156 20913 17184
rect 20680 17144 20686 17156
rect 20901 17153 20913 17156
rect 20947 17184 20959 17187
rect 21545 17187 21603 17193
rect 21545 17184 21557 17187
rect 20947 17156 21557 17184
rect 20947 17153 20959 17156
rect 20901 17147 20959 17153
rect 21545 17153 21557 17156
rect 21591 17153 21603 17187
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 21545 17147 21603 17153
rect 22204 17156 22845 17184
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 6914 17116 6920 17128
rect 6871 17088 6920 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 6914 17076 6920 17088
rect 6972 17076 6978 17128
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 10318 17116 10324 17128
rect 8619 17088 10324 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 10502 17076 10508 17128
rect 10560 17076 10566 17128
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 10870 17116 10876 17128
rect 10735 17088 10876 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 11330 17076 11336 17128
rect 11388 17116 11394 17128
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 11388 17088 12633 17116
rect 11388 17076 11394 17088
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 12897 17119 12955 17125
rect 12897 17085 12909 17119
rect 12943 17116 12955 17119
rect 13262 17116 13268 17128
rect 12943 17088 13268 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 13262 17076 13268 17088
rect 13320 17076 13326 17128
rect 13354 17076 13360 17128
rect 13412 17116 13418 17128
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 13412 17088 14933 17116
rect 13412 17076 13418 17088
rect 14921 17085 14933 17088
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 17957 17119 18015 17125
rect 17957 17085 17969 17119
rect 18003 17116 18015 17119
rect 18598 17116 18604 17128
rect 18003 17088 18604 17116
rect 18003 17085 18015 17088
rect 17957 17079 18015 17085
rect 11514 17048 11520 17060
rect 9232 17020 11520 17048
rect 9232 16989 9260 17020
rect 11514 17008 11520 17020
rect 11572 17008 11578 17060
rect 14936 17048 14964 17079
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 18690 17076 18696 17128
rect 18748 17116 18754 17128
rect 18748 17088 19288 17116
rect 18748 17076 18754 17088
rect 19260 17048 19288 17088
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 19429 17119 19487 17125
rect 19429 17116 19441 17119
rect 19392 17088 19441 17116
rect 19392 17076 19398 17088
rect 19429 17085 19441 17088
rect 19475 17085 19487 17119
rect 19429 17079 19487 17085
rect 20438 17076 20444 17128
rect 20496 17076 20502 17128
rect 22204 17048 22232 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 23750 17144 23756 17196
rect 23808 17184 23814 17196
rect 23937 17187 23995 17193
rect 23937 17184 23949 17187
rect 23808 17156 23949 17184
rect 23808 17144 23814 17156
rect 23937 17153 23949 17156
rect 23983 17153 23995 17187
rect 23937 17147 23995 17153
rect 24670 17076 24676 17128
rect 24728 17076 24734 17128
rect 14936 17020 17816 17048
rect 19260 17020 22232 17048
rect 22281 17051 22339 17057
rect 9217 16983 9275 16989
rect 9217 16949 9229 16983
rect 9263 16949 9275 16983
rect 9217 16943 9275 16949
rect 9490 16940 9496 16992
rect 9548 16940 9554 16992
rect 10318 16940 10324 16992
rect 10376 16980 10382 16992
rect 10778 16980 10784 16992
rect 10376 16952 10784 16980
rect 10376 16940 10382 16952
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 16025 16983 16083 16989
rect 16025 16980 16037 16983
rect 15068 16952 16037 16980
rect 15068 16940 15074 16952
rect 16025 16949 16037 16952
rect 16071 16980 16083 16983
rect 16574 16980 16580 16992
rect 16071 16952 16580 16980
rect 16071 16949 16083 16952
rect 16025 16943 16083 16949
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 16853 16983 16911 16989
rect 16853 16949 16865 16983
rect 16899 16980 16911 16983
rect 17310 16980 17316 16992
rect 16899 16952 17316 16980
rect 16899 16949 16911 16952
rect 16853 16943 16911 16949
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 17788 16980 17816 17020
rect 22281 17017 22293 17051
rect 22327 17048 22339 17051
rect 22646 17048 22652 17060
rect 22327 17020 22652 17048
rect 22327 17017 22339 17020
rect 22281 17011 22339 17017
rect 22646 17008 22652 17020
rect 22704 17008 22710 17060
rect 23017 17051 23075 17057
rect 23017 17017 23029 17051
rect 23063 17048 23075 17051
rect 23290 17048 23296 17060
rect 23063 17020 23296 17048
rect 23063 17017 23075 17020
rect 23017 17011 23075 17017
rect 23290 17008 23296 17020
rect 23348 17008 23354 17060
rect 17954 16980 17960 16992
rect 17788 16952 17960 16980
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 5616 16779 5674 16785
rect 5616 16745 5628 16779
rect 5662 16776 5674 16779
rect 5662 16748 6868 16776
rect 5662 16745 5674 16748
rect 5616 16739 5674 16745
rect 6840 16708 6868 16748
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7101 16779 7159 16785
rect 7101 16776 7113 16779
rect 6972 16748 7113 16776
rect 6972 16736 6978 16748
rect 7101 16745 7113 16748
rect 7147 16745 7159 16779
rect 7101 16739 7159 16745
rect 7466 16736 7472 16788
rect 7524 16776 7530 16788
rect 8294 16776 8300 16788
rect 7524 16748 8300 16776
rect 7524 16736 7530 16748
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16776 8815 16779
rect 9030 16776 9036 16788
rect 8803 16748 9036 16776
rect 8803 16745 8815 16748
rect 8757 16739 8815 16745
rect 9030 16736 9036 16748
rect 9088 16736 9094 16788
rect 12618 16776 12624 16788
rect 9692 16748 12624 16776
rect 8386 16708 8392 16720
rect 6840 16680 8392 16708
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16640 5411 16643
rect 6362 16640 6368 16652
rect 5399 16612 6368 16640
rect 5399 16609 5411 16612
rect 5353 16603 5411 16609
rect 6362 16600 6368 16612
rect 6420 16600 6426 16652
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 9214 16640 9220 16652
rect 8352 16612 9220 16640
rect 8352 16600 8358 16612
rect 9214 16600 9220 16612
rect 9272 16640 9278 16652
rect 9692 16649 9720 16748
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 21818 16736 21824 16788
rect 21876 16736 21882 16788
rect 10870 16668 10876 16720
rect 10928 16668 10934 16720
rect 14366 16708 14372 16720
rect 12268 16680 14372 16708
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 9272 16612 9689 16640
rect 9272 16600 9278 16612
rect 9677 16609 9689 16612
rect 9723 16609 9735 16643
rect 10888 16640 10916 16668
rect 12268 16649 12296 16680
rect 14366 16668 14372 16680
rect 14424 16668 14430 16720
rect 11057 16643 11115 16649
rect 11057 16640 11069 16643
rect 10888 16612 11069 16640
rect 9677 16603 9735 16609
rect 11057 16609 11069 16612
rect 11103 16609 11115 16643
rect 11057 16603 11115 16609
rect 12253 16643 12311 16649
rect 12253 16609 12265 16643
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16640 12403 16643
rect 12618 16640 12624 16652
rect 12391 16612 12624 16640
rect 12391 16609 12403 16612
rect 12345 16603 12403 16609
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 15746 16600 15752 16652
rect 15804 16600 15810 16652
rect 15930 16600 15936 16652
rect 15988 16600 15994 16652
rect 20162 16600 20168 16652
rect 20220 16640 20226 16652
rect 20625 16643 20683 16649
rect 20625 16640 20637 16643
rect 20220 16612 20637 16640
rect 20220 16600 20226 16612
rect 20625 16609 20637 16612
rect 20671 16609 20683 16643
rect 21836 16640 21864 16736
rect 22005 16643 22063 16649
rect 22005 16640 22017 16643
rect 21836 16612 22017 16640
rect 20625 16603 20683 16609
rect 22005 16609 22017 16612
rect 22051 16609 22063 16643
rect 22005 16603 22063 16609
rect 23014 16600 23020 16652
rect 23072 16640 23078 16652
rect 23382 16640 23388 16652
rect 23072 16612 23388 16640
rect 23072 16600 23078 16612
rect 1486 16532 1492 16584
rect 1544 16572 1550 16584
rect 1581 16575 1639 16581
rect 1581 16572 1593 16575
rect 1544 16544 1593 16572
rect 1544 16532 1550 16544
rect 1581 16541 1593 16544
rect 1627 16541 1639 16575
rect 1581 16535 1639 16541
rect 9306 16532 9312 16584
rect 9364 16572 9370 16584
rect 9493 16575 9551 16581
rect 9493 16572 9505 16575
rect 9364 16544 9505 16572
rect 9364 16532 9370 16544
rect 9493 16541 9505 16544
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 9582 16532 9588 16584
rect 9640 16532 9646 16584
rect 10873 16575 10931 16581
rect 10873 16541 10885 16575
rect 10919 16572 10931 16575
rect 11974 16572 11980 16584
rect 10919 16544 11980 16572
rect 10919 16541 10931 16544
rect 10873 16535 10931 16541
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16572 12219 16575
rect 12710 16572 12716 16584
rect 12207 16544 12716 16572
rect 12207 16541 12219 16544
rect 12161 16535 12219 16541
rect 12710 16532 12716 16544
rect 12768 16532 12774 16584
rect 20438 16532 20444 16584
rect 20496 16532 20502 16584
rect 20530 16532 20536 16584
rect 20588 16532 20594 16584
rect 21726 16532 21732 16584
rect 21784 16532 21790 16584
rect 23124 16546 23152 16612
rect 23382 16600 23388 16612
rect 23440 16640 23446 16652
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 23440 16612 23765 16640
rect 23440 16600 23446 16612
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 7466 16504 7472 16516
rect 6854 16476 7472 16504
rect 2501 16467 2559 16473
rect 7466 16464 7472 16476
rect 7524 16464 7530 16516
rect 7834 16464 7840 16516
rect 7892 16504 7898 16516
rect 9600 16504 9628 16532
rect 7892 16476 9168 16504
rect 9600 16476 10548 16504
rect 7892 16464 7898 16476
rect 9140 16445 9168 16476
rect 9125 16439 9183 16445
rect 9125 16405 9137 16439
rect 9171 16405 9183 16439
rect 9125 16399 9183 16405
rect 9585 16439 9643 16445
rect 9585 16405 9597 16439
rect 9631 16436 9643 16439
rect 10226 16436 10232 16448
rect 9631 16408 10232 16436
rect 9631 16405 9643 16408
rect 9585 16399 9643 16405
rect 10226 16396 10232 16408
rect 10284 16396 10290 16448
rect 10520 16445 10548 16476
rect 19518 16464 19524 16516
rect 19576 16504 19582 16516
rect 21744 16504 21772 16532
rect 19576 16476 21772 16504
rect 19576 16464 19582 16476
rect 10505 16439 10563 16445
rect 10505 16405 10517 16439
rect 10551 16405 10563 16439
rect 10505 16399 10563 16405
rect 10965 16439 11023 16445
rect 10965 16405 10977 16439
rect 11011 16436 11023 16439
rect 11698 16436 11704 16448
rect 11011 16408 11704 16436
rect 11011 16405 11023 16408
rect 10965 16399 11023 16405
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 11790 16396 11796 16448
rect 11848 16396 11854 16448
rect 14642 16396 14648 16448
rect 14700 16436 14706 16448
rect 15289 16439 15347 16445
rect 15289 16436 15301 16439
rect 14700 16408 15301 16436
rect 14700 16396 14706 16408
rect 15289 16405 15301 16408
rect 15335 16405 15347 16439
rect 15289 16399 15347 16405
rect 15657 16439 15715 16445
rect 15657 16405 15669 16439
rect 15703 16436 15715 16439
rect 16298 16436 16304 16448
rect 15703 16408 16304 16436
rect 15703 16405 15715 16408
rect 15657 16399 15715 16405
rect 16298 16396 16304 16408
rect 16356 16436 16362 16448
rect 16393 16439 16451 16445
rect 16393 16436 16405 16439
rect 16356 16408 16405 16436
rect 16356 16396 16362 16408
rect 16393 16405 16405 16408
rect 16439 16436 16451 16439
rect 17494 16436 17500 16448
rect 16439 16408 17500 16436
rect 16439 16405 16451 16408
rect 16393 16399 16451 16405
rect 17494 16396 17500 16408
rect 17552 16396 17558 16448
rect 20070 16396 20076 16448
rect 20128 16396 20134 16448
rect 21174 16396 21180 16448
rect 21232 16436 21238 16448
rect 23477 16439 23535 16445
rect 23477 16436 23489 16439
rect 21232 16408 23489 16436
rect 21232 16396 21238 16408
rect 23477 16405 23489 16408
rect 23523 16405 23535 16439
rect 23477 16399 23535 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 8941 16235 8999 16241
rect 8941 16232 8953 16235
rect 7340 16204 8953 16232
rect 7340 16192 7346 16204
rect 8941 16201 8953 16204
rect 8987 16201 8999 16235
rect 8941 16195 8999 16201
rect 10137 16235 10195 16241
rect 10137 16201 10149 16235
rect 10183 16232 10195 16235
rect 10502 16232 10508 16244
rect 10183 16204 10508 16232
rect 10183 16201 10195 16204
rect 10137 16195 10195 16201
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 10594 16192 10600 16244
rect 10652 16192 10658 16244
rect 10962 16192 10968 16244
rect 11020 16232 11026 16244
rect 11701 16235 11759 16241
rect 11701 16232 11713 16235
rect 11020 16204 11713 16232
rect 11020 16192 11026 16204
rect 11701 16201 11713 16204
rect 11747 16201 11759 16235
rect 11701 16195 11759 16201
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 13446 16232 13452 16244
rect 12584 16204 13452 16232
rect 12584 16192 12590 16204
rect 13446 16192 13452 16204
rect 13504 16232 13510 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 13504 16204 13737 16232
rect 13504 16192 13510 16204
rect 13725 16201 13737 16204
rect 13771 16201 13783 16235
rect 13725 16195 13783 16201
rect 16390 16192 16396 16244
rect 16448 16192 16454 16244
rect 16500 16204 18460 16232
rect 2498 16124 2504 16176
rect 2556 16124 2562 16176
rect 7466 16124 7472 16176
rect 7524 16124 7530 16176
rect 9309 16167 9367 16173
rect 9309 16133 9321 16167
rect 9355 16164 9367 16167
rect 11790 16164 11796 16176
rect 9355 16136 11796 16164
rect 9355 16133 9367 16136
rect 9309 16127 9367 16133
rect 11790 16124 11796 16136
rect 11848 16124 11854 16176
rect 12069 16167 12127 16173
rect 12069 16133 12081 16167
rect 12115 16164 12127 16167
rect 14274 16164 14280 16176
rect 12115 16136 14280 16164
rect 12115 16133 12127 16136
rect 12069 16127 12127 16133
rect 14274 16124 14280 16136
rect 14332 16124 14338 16176
rect 15933 16167 15991 16173
rect 15933 16133 15945 16167
rect 15979 16164 15991 16167
rect 16408 16164 16436 16192
rect 15979 16136 16436 16164
rect 15979 16133 15991 16136
rect 15933 16127 15991 16133
rect 6546 16056 6552 16108
rect 6604 16096 6610 16108
rect 6641 16099 6699 16105
rect 6641 16096 6653 16099
rect 6604 16068 6653 16096
rect 6604 16056 6610 16068
rect 6641 16065 6653 16068
rect 6687 16065 6699 16099
rect 6641 16059 6699 16065
rect 8404 16068 9536 16096
rect 8404 16040 8432 16068
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 16028 6975 16031
rect 8294 16028 8300 16040
rect 6963 16000 8300 16028
rect 6963 15997 6975 16000
rect 6917 15991 6975 15997
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 8386 15988 8392 16040
rect 8444 15988 8450 16040
rect 9508 16037 9536 16068
rect 10410 16056 10416 16108
rect 10468 16096 10474 16108
rect 10505 16099 10563 16105
rect 10505 16096 10517 16099
rect 10468 16068 10517 16096
rect 10468 16056 10474 16068
rect 10505 16065 10517 16068
rect 10551 16065 10563 16099
rect 10505 16059 10563 16065
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12802 16096 12808 16108
rect 12207 16068 12808 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 14182 16056 14188 16108
rect 14240 16096 14246 16108
rect 14645 16099 14703 16105
rect 14645 16096 14657 16099
rect 14240 16068 14657 16096
rect 14240 16056 14246 16068
rect 14645 16065 14657 16068
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 16298 16096 16304 16108
rect 15804 16068 16304 16096
rect 15804 16056 15810 16068
rect 16298 16056 16304 16068
rect 16356 16096 16362 16108
rect 16500 16096 16528 16204
rect 17126 16124 17132 16176
rect 17184 16124 17190 16176
rect 17862 16124 17868 16176
rect 17920 16124 17926 16176
rect 18432 16164 18460 16204
rect 18598 16192 18604 16244
rect 18656 16192 18662 16244
rect 19242 16192 19248 16244
rect 19300 16192 19306 16244
rect 20070 16192 20076 16244
rect 20128 16232 20134 16244
rect 22830 16232 22836 16244
rect 20128 16204 22836 16232
rect 20128 16192 20134 16204
rect 22830 16192 22836 16204
rect 22888 16192 22894 16244
rect 19705 16167 19763 16173
rect 19705 16164 19717 16167
rect 18432 16136 19717 16164
rect 19705 16133 19717 16136
rect 19751 16133 19763 16167
rect 22094 16164 22100 16176
rect 19705 16127 19763 16133
rect 20916 16136 22100 16164
rect 16356 16068 16528 16096
rect 16356 16056 16362 16068
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16632 16068 16865 16096
rect 16632 16056 16638 16068
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 18138 16056 18144 16108
rect 18196 16096 18202 16108
rect 18877 16099 18935 16105
rect 18877 16096 18889 16099
rect 18196 16068 18889 16096
rect 18196 16056 18202 16068
rect 18877 16065 18889 16068
rect 18923 16065 18935 16099
rect 18877 16059 18935 16065
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16096 19671 16099
rect 20441 16099 20499 16105
rect 20441 16096 20453 16099
rect 19659 16068 20453 16096
rect 19659 16065 19671 16068
rect 19613 16059 19671 16065
rect 20441 16065 20453 16068
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 9401 16031 9459 16037
rect 9401 15997 9413 16031
rect 9447 15997 9459 16031
rect 9401 15991 9459 15997
rect 9493 16031 9551 16037
rect 9493 15997 9505 16031
rect 9539 15997 9551 16031
rect 9493 15991 9551 15997
rect 1762 15852 1768 15904
rect 1820 15892 1826 15904
rect 2593 15895 2651 15901
rect 2593 15892 2605 15895
rect 1820 15864 2605 15892
rect 1820 15852 1826 15864
rect 2593 15861 2605 15864
rect 2639 15861 2651 15895
rect 9416 15892 9444 15991
rect 10226 15988 10232 16040
rect 10284 16028 10290 16040
rect 10689 16031 10747 16037
rect 10689 16028 10701 16031
rect 10284 16000 10701 16028
rect 10284 15988 10290 16000
rect 10689 15997 10701 16000
rect 10735 15997 10747 16031
rect 10689 15991 10747 15997
rect 11882 15988 11888 16040
rect 11940 16028 11946 16040
rect 12253 16031 12311 16037
rect 12253 16028 12265 16031
rect 11940 16000 12265 16028
rect 11940 15988 11946 16000
rect 12253 15997 12265 16000
rect 12299 15997 12311 16031
rect 12253 15991 12311 15997
rect 15470 15988 15476 16040
rect 15528 16028 15534 16040
rect 19889 16031 19947 16037
rect 15528 16000 19656 16028
rect 15528 15988 15534 16000
rect 10962 15920 10968 15972
rect 11020 15960 11026 15972
rect 13998 15960 14004 15972
rect 11020 15932 14004 15960
rect 11020 15920 11026 15932
rect 13998 15920 14004 15932
rect 14056 15920 14062 15972
rect 19628 15960 19656 16000
rect 19889 15997 19901 16031
rect 19935 16028 19947 16031
rect 20916 16028 20944 16136
rect 22094 16124 22100 16136
rect 22152 16124 22158 16176
rect 22462 16124 22468 16176
rect 22520 16124 22526 16176
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 19935 16000 20944 16028
rect 19935 15997 19947 16000
rect 19889 15991 19947 15997
rect 21284 15960 21312 16059
rect 22370 16056 22376 16108
rect 22428 16056 22434 16108
rect 22480 16096 22508 16124
rect 23385 16099 23443 16105
rect 23385 16096 23397 16099
rect 22480 16068 23397 16096
rect 23385 16065 23397 16068
rect 23431 16065 23443 16099
rect 23385 16059 23443 16065
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16096 24179 16099
rect 24210 16096 24216 16108
rect 24167 16068 24216 16096
rect 24167 16065 24179 16068
rect 24121 16059 24179 16065
rect 24210 16056 24216 16068
rect 24268 16056 24274 16108
rect 21542 15988 21548 16040
rect 21600 16028 21606 16040
rect 22465 16031 22523 16037
rect 22465 16028 22477 16031
rect 21600 16000 22477 16028
rect 21600 15988 21606 16000
rect 22465 15997 22477 16000
rect 22511 15997 22523 16031
rect 22465 15991 22523 15997
rect 22649 16031 22707 16037
rect 22649 15997 22661 16031
rect 22695 16028 22707 16031
rect 22738 16028 22744 16040
rect 22695 16000 22744 16028
rect 22695 15997 22707 16000
rect 22649 15991 22707 15997
rect 22738 15988 22744 16000
rect 22796 15988 22802 16040
rect 24762 15988 24768 16040
rect 24820 15988 24826 16040
rect 19628 15932 21312 15960
rect 21453 15963 21511 15969
rect 21453 15929 21465 15963
rect 21499 15960 21511 15963
rect 22554 15960 22560 15972
rect 21499 15932 22560 15960
rect 21499 15929 21511 15932
rect 21453 15923 21511 15929
rect 22554 15920 22560 15932
rect 22612 15920 22618 15972
rect 12342 15892 12348 15904
rect 9416 15864 12348 15892
rect 2593 15855 2651 15861
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 12618 15852 12624 15904
rect 12676 15892 12682 15904
rect 12989 15895 13047 15901
rect 12989 15892 13001 15895
rect 12676 15864 13001 15892
rect 12676 15852 12682 15864
rect 12989 15861 13001 15864
rect 13035 15861 13047 15895
rect 12989 15855 13047 15861
rect 14274 15852 14280 15904
rect 14332 15852 14338 15904
rect 15194 15852 15200 15904
rect 15252 15892 15258 15904
rect 16025 15895 16083 15901
rect 16025 15892 16037 15895
rect 15252 15864 16037 15892
rect 15252 15852 15258 15864
rect 16025 15861 16037 15864
rect 16071 15861 16083 15895
rect 16025 15855 16083 15861
rect 21910 15852 21916 15904
rect 21968 15892 21974 15904
rect 22005 15895 22063 15901
rect 22005 15892 22017 15895
rect 21968 15864 22017 15892
rect 21968 15852 21974 15864
rect 22005 15861 22017 15864
rect 22051 15861 22063 15895
rect 22005 15855 22063 15861
rect 22094 15852 22100 15904
rect 22152 15892 22158 15904
rect 23201 15895 23259 15901
rect 23201 15892 23213 15895
rect 22152 15864 23213 15892
rect 22152 15852 22158 15864
rect 23201 15861 23213 15864
rect 23247 15861 23259 15895
rect 23201 15855 23259 15861
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 7466 15648 7472 15700
rect 7524 15688 7530 15700
rect 8481 15691 8539 15697
rect 8481 15688 8493 15691
rect 7524 15660 8493 15688
rect 7524 15648 7530 15660
rect 8481 15657 8493 15660
rect 8527 15688 8539 15691
rect 9306 15688 9312 15700
rect 8527 15660 9312 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 11756 15660 14289 15688
rect 11756 15648 11762 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 17218 15648 17224 15700
rect 17276 15688 17282 15700
rect 20806 15688 20812 15700
rect 17276 15660 20812 15688
rect 17276 15648 17282 15660
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 20990 15648 20996 15700
rect 21048 15688 21054 15700
rect 22094 15688 22100 15700
rect 21048 15660 22100 15688
rect 21048 15648 21054 15660
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 12434 15580 12440 15632
rect 12492 15620 12498 15632
rect 13633 15623 13691 15629
rect 13633 15620 13645 15623
rect 12492 15592 13645 15620
rect 12492 15580 12498 15592
rect 13633 15589 13645 15592
rect 13679 15589 13691 15623
rect 13633 15583 13691 15589
rect 17313 15623 17371 15629
rect 17313 15589 17325 15623
rect 17359 15620 17371 15623
rect 19886 15620 19892 15632
rect 17359 15592 19892 15620
rect 17359 15589 17371 15592
rect 17313 15583 17371 15589
rect 19886 15580 19892 15592
rect 19944 15580 19950 15632
rect 19978 15580 19984 15632
rect 20036 15620 20042 15632
rect 21085 15623 21143 15629
rect 21085 15620 21097 15623
rect 20036 15592 21097 15620
rect 20036 15580 20042 15592
rect 21085 15589 21097 15592
rect 21131 15589 21143 15623
rect 21085 15583 21143 15589
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15552 11115 15555
rect 11330 15552 11336 15564
rect 11103 15524 11336 15552
rect 11103 15521 11115 15524
rect 11057 15515 11115 15521
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 14090 15512 14096 15564
rect 14148 15552 14154 15564
rect 14829 15555 14887 15561
rect 14829 15552 14841 15555
rect 14148 15524 14841 15552
rect 14148 15512 14154 15524
rect 14829 15521 14841 15524
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 17402 15512 17408 15564
rect 17460 15552 17466 15564
rect 17865 15555 17923 15561
rect 17865 15552 17877 15555
rect 17460 15524 17877 15552
rect 17460 15512 17466 15524
rect 17865 15521 17877 15524
rect 17911 15521 17923 15555
rect 17865 15515 17923 15521
rect 20073 15555 20131 15561
rect 20073 15521 20085 15555
rect 20119 15552 20131 15555
rect 21174 15552 21180 15564
rect 20119 15524 21180 15552
rect 20119 15521 20131 15524
rect 20073 15515 20131 15521
rect 21174 15512 21180 15524
rect 21232 15512 21238 15564
rect 12618 15484 12624 15496
rect 12466 15456 12624 15484
rect 12618 15444 12624 15456
rect 12676 15444 12682 15496
rect 13446 15444 13452 15496
rect 13504 15444 13510 15496
rect 14642 15444 14648 15496
rect 14700 15444 14706 15496
rect 16114 15444 16120 15496
rect 16172 15484 16178 15496
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 16172 15456 17785 15484
rect 16172 15444 16178 15456
rect 17773 15453 17785 15456
rect 17819 15484 17831 15487
rect 18325 15487 18383 15493
rect 18325 15484 18337 15487
rect 17819 15456 18337 15484
rect 17819 15453 17831 15456
rect 17773 15447 17831 15453
rect 18325 15453 18337 15456
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15484 19947 15487
rect 19978 15484 19984 15496
rect 19935 15456 19984 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 20809 15487 20867 15493
rect 20809 15453 20821 15487
rect 20855 15484 20867 15487
rect 22278 15484 22284 15496
rect 20855 15456 22284 15484
rect 20855 15453 20867 15456
rect 20809 15447 20867 15453
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 22833 15487 22891 15493
rect 22833 15453 22845 15487
rect 22879 15484 22891 15487
rect 24302 15484 24308 15496
rect 22879 15456 24308 15484
rect 22879 15453 22891 15456
rect 22833 15447 22891 15453
rect 24302 15444 24308 15456
rect 24360 15444 24366 15496
rect 10962 15376 10968 15428
rect 11020 15416 11026 15428
rect 11333 15419 11391 15425
rect 11333 15416 11345 15419
rect 11020 15388 11345 15416
rect 11020 15376 11026 15388
rect 11333 15385 11345 15388
rect 11379 15385 11391 15419
rect 14090 15416 14096 15428
rect 11333 15379 11391 15385
rect 12636 15388 14096 15416
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 12636 15348 12664 15388
rect 14090 15376 14096 15388
rect 14148 15376 14154 15428
rect 21266 15416 21272 15428
rect 19444 15388 21272 15416
rect 10284 15320 12664 15348
rect 10284 15308 10290 15320
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 12805 15351 12863 15357
rect 12805 15348 12817 15351
rect 12768 15320 12817 15348
rect 12768 15308 12774 15320
rect 12805 15317 12817 15320
rect 12851 15317 12863 15351
rect 12805 15311 12863 15317
rect 14737 15351 14795 15357
rect 14737 15317 14749 15351
rect 14783 15348 14795 15351
rect 15654 15348 15660 15360
rect 14783 15320 15660 15348
rect 14783 15317 14795 15320
rect 14737 15311 14795 15317
rect 15654 15308 15660 15320
rect 15712 15308 15718 15360
rect 16666 15308 16672 15360
rect 16724 15348 16730 15360
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 16724 15320 17693 15348
rect 16724 15308 16730 15320
rect 17681 15317 17693 15320
rect 17727 15317 17739 15351
rect 17681 15311 17739 15317
rect 18690 15308 18696 15360
rect 18748 15308 18754 15360
rect 19444 15357 19472 15388
rect 21266 15376 21272 15388
rect 21324 15376 21330 15428
rect 21821 15419 21879 15425
rect 21821 15416 21833 15419
rect 21376 15388 21833 15416
rect 19429 15351 19487 15357
rect 19429 15317 19441 15351
rect 19475 15317 19487 15351
rect 19429 15311 19487 15317
rect 19610 15308 19616 15360
rect 19668 15348 19674 15360
rect 19797 15351 19855 15357
rect 19797 15348 19809 15351
rect 19668 15320 19809 15348
rect 19668 15308 19674 15320
rect 19797 15317 19809 15320
rect 19843 15317 19855 15351
rect 19797 15311 19855 15317
rect 20622 15308 20628 15360
rect 20680 15308 20686 15360
rect 20806 15308 20812 15360
rect 20864 15348 20870 15360
rect 21376 15348 21404 15388
rect 21821 15385 21833 15388
rect 21867 15385 21879 15419
rect 21821 15379 21879 15385
rect 23845 15419 23903 15425
rect 23845 15385 23857 15419
rect 23891 15416 23903 15419
rect 24946 15416 24952 15428
rect 23891 15388 24952 15416
rect 23891 15385 23903 15388
rect 23845 15379 23903 15385
rect 24946 15376 24952 15388
rect 25004 15376 25010 15428
rect 20864 15320 21404 15348
rect 20864 15308 20870 15320
rect 21542 15308 21548 15360
rect 21600 15348 21606 15360
rect 21913 15351 21971 15357
rect 21913 15348 21925 15351
rect 21600 15320 21925 15348
rect 21600 15308 21606 15320
rect 21913 15317 21925 15320
rect 21959 15317 21971 15351
rect 21913 15311 21971 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 2682 15104 2688 15156
rect 2740 15144 2746 15156
rect 8570 15144 8576 15156
rect 2740 15116 8576 15144
rect 2740 15104 2746 15116
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 9306 15104 9312 15156
rect 9364 15144 9370 15156
rect 9364 15116 9536 15144
rect 9364 15104 9370 15116
rect 9398 15036 9404 15088
rect 9456 15036 9462 15088
rect 9508 15076 9536 15116
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 9824 15116 11529 15144
rect 9824 15104 9830 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 9784 15076 9812 15104
rect 9508 15048 9890 15076
rect 10962 15036 10968 15088
rect 11020 15076 11026 15088
rect 11149 15079 11207 15085
rect 11149 15076 11161 15079
rect 11020 15048 11161 15076
rect 11020 15036 11026 15048
rect 11149 15045 11161 15048
rect 11195 15045 11207 15079
rect 11532 15076 11560 15107
rect 12158 15104 12164 15156
rect 12216 15144 12222 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12216 15116 13001 15144
rect 12216 15104 12222 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 14185 15147 14243 15153
rect 14185 15113 14197 15147
rect 14231 15144 14243 15147
rect 17034 15144 17040 15156
rect 14231 15116 17040 15144
rect 14231 15113 14243 15116
rect 14185 15107 14243 15113
rect 17034 15104 17040 15116
rect 17092 15104 17098 15156
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 18748 15116 18797 15144
rect 18748 15104 18754 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 18785 15107 18843 15113
rect 18874 15104 18880 15156
rect 18932 15104 18938 15156
rect 22281 15147 22339 15153
rect 22281 15113 22293 15147
rect 22327 15144 22339 15147
rect 22370 15144 22376 15156
rect 22327 15116 22376 15144
rect 22327 15113 22339 15116
rect 22281 15107 22339 15113
rect 22370 15104 22376 15116
rect 22428 15104 22434 15156
rect 11974 15076 11980 15088
rect 11532 15048 11980 15076
rect 11149 15039 11207 15045
rect 11974 15036 11980 15048
rect 12032 15076 12038 15088
rect 12618 15076 12624 15088
rect 12032 15048 12624 15076
rect 12032 15036 12038 15048
rect 12618 15036 12624 15048
rect 12676 15036 12682 15088
rect 13446 15036 13452 15088
rect 13504 15076 13510 15088
rect 16666 15076 16672 15088
rect 13504 15048 16672 15076
rect 13504 15036 13510 15048
rect 16666 15036 16672 15048
rect 16724 15036 16730 15088
rect 16758 15036 16764 15088
rect 16816 15076 16822 15088
rect 17221 15079 17279 15085
rect 17221 15076 17233 15079
rect 16816 15048 17233 15076
rect 16816 15036 16822 15048
rect 17221 15045 17233 15048
rect 17267 15076 17279 15079
rect 17681 15079 17739 15085
rect 17681 15076 17693 15079
rect 17267 15048 17693 15076
rect 17267 15045 17279 15048
rect 17221 15039 17279 15045
rect 17681 15045 17693 15048
rect 17727 15045 17739 15079
rect 17681 15039 17739 15045
rect 13354 14968 13360 15020
rect 13412 14968 13418 15020
rect 14550 14968 14556 15020
rect 14608 14968 14614 15020
rect 14645 15011 14703 15017
rect 14645 14977 14657 15011
rect 14691 15008 14703 15011
rect 15657 15011 15715 15017
rect 14691 14980 15332 15008
rect 14691 14977 14703 14980
rect 14645 14971 14703 14977
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14909 9183 14943
rect 9125 14903 9183 14909
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13814 14940 13820 14952
rect 13679 14912 13820 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 9140 14804 9168 14903
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 14826 14900 14832 14952
rect 14884 14900 14890 14952
rect 15304 14949 15332 14980
rect 15657 14977 15669 15011
rect 15703 15008 15715 15011
rect 16022 15008 16028 15020
rect 15703 14980 16028 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 16022 14968 16028 14980
rect 16080 15008 16086 15020
rect 16209 15011 16267 15017
rect 16209 15008 16221 15011
rect 16080 14980 16221 15008
rect 16080 14968 16086 14980
rect 16209 14977 16221 14980
rect 16255 14977 16267 15011
rect 16209 14971 16267 14977
rect 18598 14968 18604 15020
rect 18656 15008 18662 15020
rect 18656 14980 19012 15008
rect 18656 14968 18662 14980
rect 15289 14943 15347 14949
rect 15289 14909 15301 14943
rect 15335 14940 15347 14943
rect 16114 14940 16120 14952
rect 15335 14912 16120 14940
rect 15335 14909 15347 14912
rect 15289 14903 15347 14909
rect 16114 14900 16120 14912
rect 16172 14900 16178 14952
rect 18984 14949 19012 14980
rect 19794 14968 19800 15020
rect 19852 14968 19858 15020
rect 23842 14968 23848 15020
rect 23900 15008 23906 15020
rect 23937 15011 23995 15017
rect 23937 15008 23949 15011
rect 23900 14980 23949 15008
rect 23900 14968 23906 14980
rect 23937 14977 23949 14980
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14909 19027 14943
rect 18969 14903 19027 14909
rect 24670 14900 24676 14952
rect 24728 14900 24734 14952
rect 15841 14875 15899 14881
rect 15841 14841 15853 14875
rect 15887 14872 15899 14875
rect 16850 14872 16856 14884
rect 15887 14844 16856 14872
rect 15887 14841 15899 14844
rect 15841 14835 15899 14841
rect 16850 14832 16856 14844
rect 16908 14832 16914 14884
rect 17494 14832 17500 14884
rect 17552 14872 17558 14884
rect 20806 14872 20812 14884
rect 17552 14844 20812 14872
rect 17552 14832 17558 14844
rect 20806 14832 20812 14844
rect 20864 14832 20870 14884
rect 9950 14804 9956 14816
rect 9140 14776 9956 14804
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 13722 14804 13728 14816
rect 13320 14776 13728 14804
rect 13320 14764 13326 14776
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 16666 14764 16672 14816
rect 16724 14804 16730 14816
rect 17313 14807 17371 14813
rect 17313 14804 17325 14807
rect 16724 14776 17325 14804
rect 16724 14764 16730 14776
rect 17313 14773 17325 14776
rect 17359 14773 17371 14807
rect 17313 14767 17371 14773
rect 18417 14807 18475 14813
rect 18417 14773 18429 14807
rect 18463 14804 18475 14807
rect 19334 14804 19340 14816
rect 18463 14776 19340 14804
rect 18463 14773 18475 14776
rect 18417 14767 18475 14773
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 19613 14807 19671 14813
rect 19613 14773 19625 14807
rect 19659 14804 19671 14807
rect 20438 14804 20444 14816
rect 19659 14776 20444 14804
rect 19659 14773 19671 14776
rect 19613 14767 19671 14773
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10778 14600 10784 14612
rect 9916 14572 10784 14600
rect 9916 14560 9922 14572
rect 10778 14560 10784 14572
rect 10836 14600 10842 14612
rect 10836 14572 12434 14600
rect 10836 14560 10842 14572
rect 11330 14492 11336 14544
rect 11388 14492 11394 14544
rect 11974 14492 11980 14544
rect 12032 14492 12038 14544
rect 12406 14532 12434 14572
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12860 14572 13001 14600
rect 12860 14560 12866 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 15344 14572 17080 14600
rect 15344 14560 15350 14572
rect 14093 14535 14151 14541
rect 14093 14532 14105 14535
rect 12406 14504 14105 14532
rect 14093 14501 14105 14504
rect 14139 14532 14151 14535
rect 14550 14532 14556 14544
rect 14139 14504 14556 14532
rect 14139 14501 14151 14504
rect 14093 14495 14151 14501
rect 14550 14492 14556 14504
rect 14608 14492 14614 14544
rect 17052 14532 17080 14572
rect 17126 14560 17132 14612
rect 17184 14560 17190 14612
rect 19426 14532 19432 14544
rect 17052 14504 19432 14532
rect 19426 14492 19432 14504
rect 19484 14492 19490 14544
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 11348 14464 11376 14492
rect 10008 14436 11376 14464
rect 10008 14424 10014 14436
rect 11992 14396 12020 14492
rect 12618 14424 12624 14476
rect 12676 14464 12682 14476
rect 13446 14464 13452 14476
rect 12676 14436 13452 14464
rect 12676 14424 12682 14436
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 14734 14464 14740 14476
rect 13587 14436 14740 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 11362 14368 12020 14396
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14396 12771 14399
rect 13556 14396 13584 14427
rect 14734 14424 14740 14436
rect 14792 14424 14798 14476
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 16390 14464 16396 14476
rect 15436 14436 16396 14464
rect 15436 14424 15442 14436
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 21174 14424 21180 14476
rect 21232 14424 21238 14476
rect 12759 14368 13584 14396
rect 18233 14399 18291 14405
rect 12759 14365 12771 14368
rect 12713 14359 12771 14365
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 18598 14396 18604 14408
rect 18279 14368 18604 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 19518 14356 19524 14408
rect 19576 14396 19582 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 19576 14368 20913 14396
rect 19576 14356 19582 14368
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 10226 14288 10232 14340
rect 10284 14288 10290 14340
rect 13354 14288 13360 14340
rect 13412 14328 13418 14340
rect 15657 14331 15715 14337
rect 13412 14300 14688 14328
rect 13412 14288 13418 14300
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 10870 14260 10876 14272
rect 9916 14232 10876 14260
rect 9916 14220 9922 14232
rect 10870 14220 10876 14232
rect 10928 14260 10934 14272
rect 11701 14263 11759 14269
rect 11701 14260 11713 14263
rect 10928 14232 11713 14260
rect 10928 14220 10934 14232
rect 11701 14229 11713 14232
rect 11747 14229 11759 14263
rect 14660 14260 14688 14300
rect 15657 14297 15669 14331
rect 15703 14328 15715 14331
rect 15930 14328 15936 14340
rect 15703 14300 15936 14328
rect 15703 14297 15715 14300
rect 15657 14291 15715 14297
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 18785 14331 18843 14337
rect 16882 14300 17540 14328
rect 15562 14260 15568 14272
rect 14660 14232 15568 14260
rect 11701 14223 11759 14229
rect 15562 14220 15568 14232
rect 15620 14260 15626 14272
rect 16390 14260 16396 14272
rect 15620 14232 16396 14260
rect 15620 14220 15626 14232
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 16960 14260 16988 14300
rect 17512 14269 17540 14300
rect 18785 14297 18797 14331
rect 18831 14328 18843 14331
rect 21082 14328 21088 14340
rect 18831 14300 21088 14328
rect 18831 14297 18843 14300
rect 18785 14291 18843 14297
rect 21082 14288 21088 14300
rect 21140 14288 21146 14340
rect 23382 14328 23388 14340
rect 22402 14300 23388 14328
rect 22940 14272 22968 14300
rect 23382 14288 23388 14300
rect 23440 14288 23446 14340
rect 16540 14232 16988 14260
rect 17497 14263 17555 14269
rect 16540 14220 16546 14232
rect 17497 14229 17509 14263
rect 17543 14260 17555 14263
rect 18506 14260 18512 14272
rect 17543 14232 18512 14260
rect 17543 14229 17555 14232
rect 17497 14223 17555 14229
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 19426 14220 19432 14272
rect 19484 14220 19490 14272
rect 19978 14220 19984 14272
rect 20036 14260 20042 14272
rect 20254 14260 20260 14272
rect 20036 14232 20260 14260
rect 20036 14220 20042 14232
rect 20254 14220 20260 14232
rect 20312 14220 20318 14272
rect 21818 14220 21824 14272
rect 21876 14260 21882 14272
rect 22649 14263 22707 14269
rect 22649 14260 22661 14263
rect 21876 14232 22661 14260
rect 21876 14220 21882 14232
rect 22649 14229 22661 14232
rect 22695 14229 22707 14263
rect 22649 14223 22707 14229
rect 22922 14220 22928 14272
rect 22980 14220 22986 14272
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 9950 14056 9956 14068
rect 8128 14028 9956 14056
rect 8128 13988 8156 14028
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10778 14056 10784 14068
rect 10192 14028 10784 14056
rect 10192 14016 10198 14028
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 12158 14016 12164 14068
rect 12216 14056 12222 14068
rect 12253 14059 12311 14065
rect 12253 14056 12265 14059
rect 12216 14028 12265 14056
rect 12216 14016 12222 14028
rect 12253 14025 12265 14028
rect 12299 14025 12311 14059
rect 12253 14019 12311 14025
rect 12713 14059 12771 14065
rect 12713 14025 12725 14059
rect 12759 14056 12771 14059
rect 13722 14056 13728 14068
rect 12759 14028 13728 14056
rect 12759 14025 12771 14028
rect 12713 14019 12771 14025
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 17586 14016 17592 14068
rect 17644 14056 17650 14068
rect 19610 14056 19616 14068
rect 17644 14028 19616 14056
rect 17644 14016 17650 14028
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 21174 14016 21180 14068
rect 21232 14056 21238 14068
rect 21450 14056 21456 14068
rect 21232 14028 21456 14056
rect 21232 14016 21238 14028
rect 21450 14016 21456 14028
rect 21508 14056 21514 14068
rect 21821 14059 21879 14065
rect 21821 14056 21833 14059
rect 21508 14028 21833 14056
rect 21508 14016 21514 14028
rect 21821 14025 21833 14028
rect 21867 14025 21879 14059
rect 21821 14019 21879 14025
rect 23017 14059 23075 14065
rect 23017 14025 23029 14059
rect 23063 14056 23075 14059
rect 23382 14056 23388 14068
rect 23063 14028 23388 14056
rect 23063 14025 23075 14028
rect 23017 14019 23075 14025
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 9766 13988 9772 14000
rect 8036 13960 8156 13988
rect 9522 13960 9772 13988
rect 1762 13880 1768 13932
rect 1820 13880 1826 13932
rect 1854 13880 1860 13932
rect 1912 13920 1918 13932
rect 5442 13920 5448 13932
rect 1912 13892 5448 13920
rect 1912 13880 1918 13892
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 8036 13929 8064 13960
rect 9766 13948 9772 13960
rect 9824 13988 9830 14000
rect 10045 13991 10103 13997
rect 10045 13988 10057 13991
rect 9824 13960 10057 13988
rect 9824 13948 9830 13960
rect 10045 13957 10057 13960
rect 10091 13957 10103 13991
rect 10045 13951 10103 13957
rect 11238 13948 11244 14000
rect 11296 13988 11302 14000
rect 13541 13991 13599 13997
rect 13541 13988 13553 13991
rect 11296 13960 13553 13988
rect 11296 13948 11302 13960
rect 13541 13957 13553 13960
rect 13587 13988 13599 13991
rect 14001 13991 14059 13997
rect 14001 13988 14013 13991
rect 13587 13960 14013 13988
rect 13587 13957 13599 13960
rect 13541 13951 13599 13957
rect 14001 13957 14013 13960
rect 14047 13957 14059 13991
rect 14001 13951 14059 13957
rect 17402 13948 17408 14000
rect 17460 13948 17466 14000
rect 19705 13991 19763 13997
rect 19705 13957 19717 13991
rect 19751 13988 19763 13991
rect 19978 13988 19984 14000
rect 19751 13960 19984 13988
rect 19751 13957 19763 13960
rect 19705 13951 19763 13957
rect 19978 13948 19984 13960
rect 20036 13948 20042 14000
rect 20714 13948 20720 14000
rect 20772 13988 20778 14000
rect 21361 13991 21419 13997
rect 20772 13960 21312 13988
rect 20772 13948 20778 13960
rect 8021 13923 8079 13929
rect 8021 13889 8033 13923
rect 8067 13889 8079 13923
rect 8021 13883 8079 13889
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 10410 13920 10416 13932
rect 9640 13892 10416 13920
rect 9640 13880 9646 13892
rect 10410 13880 10416 13892
rect 10468 13920 10474 13932
rect 12621 13923 12679 13929
rect 12621 13920 12633 13923
rect 10468 13892 12633 13920
rect 10468 13880 10474 13892
rect 12621 13889 12633 13892
rect 12667 13889 12679 13923
rect 12621 13883 12679 13889
rect 16574 13880 16580 13932
rect 16632 13920 16638 13932
rect 17126 13920 17132 13932
rect 16632 13892 17132 13920
rect 16632 13880 16638 13892
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 18506 13880 18512 13932
rect 18564 13920 18570 13932
rect 18564 13892 19288 13920
rect 18564 13880 18570 13892
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 9769 13855 9827 13861
rect 9769 13852 9781 13855
rect 9548 13824 9781 13852
rect 9548 13812 9554 13824
rect 9769 13821 9781 13824
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 12805 13855 12863 13861
rect 12805 13821 12817 13855
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 11790 13744 11796 13796
rect 11848 13784 11854 13796
rect 12820 13784 12848 13815
rect 13446 13812 13452 13864
rect 13504 13852 13510 13864
rect 13725 13855 13783 13861
rect 13725 13852 13737 13855
rect 13504 13824 13737 13852
rect 13504 13812 13510 13824
rect 13725 13821 13737 13824
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 18877 13855 18935 13861
rect 18877 13821 18889 13855
rect 18923 13852 18935 13855
rect 19150 13852 19156 13864
rect 18923 13824 19156 13852
rect 18923 13821 18935 13824
rect 18877 13815 18935 13821
rect 19150 13812 19156 13824
rect 19208 13812 19214 13864
rect 19260 13861 19288 13892
rect 20346 13880 20352 13932
rect 20404 13920 20410 13932
rect 20441 13923 20499 13929
rect 20441 13920 20453 13923
rect 20404 13892 20453 13920
rect 20404 13880 20410 13892
rect 20441 13889 20453 13892
rect 20487 13889 20499 13923
rect 20441 13883 20499 13889
rect 21174 13880 21180 13932
rect 21232 13880 21238 13932
rect 21284 13920 21312 13960
rect 21361 13957 21373 13991
rect 21407 13988 21419 13991
rect 21726 13988 21732 14000
rect 21407 13960 21732 13988
rect 21407 13957 21419 13960
rect 21361 13951 21419 13957
rect 21726 13948 21732 13960
rect 21784 13948 21790 14000
rect 22186 13948 22192 14000
rect 22244 13988 22250 14000
rect 22244 13960 23980 13988
rect 22244 13948 22250 13960
rect 23952 13929 23980 13960
rect 25130 13948 25136 14000
rect 25188 13948 25194 14000
rect 23201 13923 23259 13929
rect 23201 13920 23213 13923
rect 21284 13892 23213 13920
rect 23201 13889 23213 13892
rect 23247 13889 23259 13923
rect 23201 13883 23259 13889
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13852 19303 13855
rect 19889 13855 19947 13861
rect 19291 13824 19564 13852
rect 19291 13821 19303 13824
rect 19245 13815 19303 13821
rect 11848 13756 12848 13784
rect 19536 13784 19564 13824
rect 19889 13821 19901 13855
rect 19935 13852 19947 13855
rect 20162 13852 20168 13864
rect 19935 13824 20168 13852
rect 19935 13821 19947 13824
rect 19889 13815 19947 13821
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20530 13812 20536 13864
rect 20588 13852 20594 13864
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20588 13824 20637 13852
rect 20588 13812 20594 13824
rect 20625 13821 20637 13824
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 21358 13812 21364 13864
rect 21416 13852 21422 13864
rect 23750 13852 23756 13864
rect 21416 13824 23756 13852
rect 21416 13812 21422 13824
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 19536 13756 22048 13784
rect 11848 13744 11854 13756
rect 22020 13728 22048 13756
rect 8284 13719 8342 13725
rect 8284 13685 8296 13719
rect 8330 13716 8342 13719
rect 9858 13716 9864 13728
rect 8330 13688 9864 13716
rect 8330 13685 8342 13688
rect 8284 13679 8342 13685
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 22002 13676 22008 13728
rect 22060 13716 22066 13728
rect 22922 13716 22928 13728
rect 22060 13688 22928 13716
rect 22060 13676 22066 13688
rect 22922 13676 22928 13688
rect 22980 13676 22986 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 5868 13484 9996 13512
rect 5868 13472 5874 13484
rect 9033 13447 9091 13453
rect 9033 13413 9045 13447
rect 9079 13444 9091 13447
rect 9766 13444 9772 13456
rect 9079 13416 9772 13444
rect 9079 13413 9091 13416
rect 9033 13407 9091 13413
rect 6546 13336 6552 13388
rect 6604 13376 6610 13388
rect 6822 13376 6828 13388
rect 6604 13348 6828 13376
rect 6604 13336 6610 13348
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7558 13376 7564 13388
rect 7156 13348 7564 13376
rect 7156 13336 7162 13348
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 9048 13308 9076 13407
rect 9766 13404 9772 13416
rect 9824 13404 9830 13456
rect 9858 13336 9864 13388
rect 9916 13336 9922 13388
rect 9968 13376 9996 13484
rect 11514 13472 11520 13524
rect 11572 13512 11578 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 11572 13484 11621 13512
rect 11572 13472 11578 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 11609 13475 11667 13481
rect 11974 13472 11980 13524
rect 12032 13472 12038 13524
rect 12342 13472 12348 13524
rect 12400 13472 12406 13524
rect 13449 13515 13507 13521
rect 13449 13481 13461 13515
rect 13495 13512 13507 13515
rect 13722 13512 13728 13524
rect 13495 13484 13728 13512
rect 13495 13481 13507 13484
rect 13449 13475 13507 13481
rect 13722 13472 13728 13484
rect 13780 13512 13786 13524
rect 13780 13484 15884 13512
rect 13780 13472 13786 13484
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 9968 13348 10149 13376
rect 10137 13345 10149 13348
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 12710 13336 12716 13388
rect 12768 13376 12774 13388
rect 12897 13379 12955 13385
rect 12897 13376 12909 13379
rect 12768 13348 12909 13376
rect 12768 13336 12774 13348
rect 12897 13345 12909 13348
rect 12943 13345 12955 13379
rect 12897 13339 12955 13345
rect 14553 13379 14611 13385
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15378 13376 15384 13388
rect 14599 13348 15384 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 15856 13376 15884 13484
rect 15930 13472 15936 13524
rect 15988 13512 15994 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 15988 13484 16313 13512
rect 15988 13472 15994 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 20346 13472 20352 13524
rect 20404 13512 20410 13524
rect 20717 13515 20775 13521
rect 20717 13512 20729 13515
rect 20404 13484 20729 13512
rect 20404 13472 20410 13484
rect 20717 13481 20729 13484
rect 20763 13481 20775 13515
rect 20717 13475 20775 13481
rect 18322 13404 18328 13456
rect 18380 13444 18386 13456
rect 18874 13444 18880 13456
rect 18380 13416 18880 13444
rect 18380 13404 18386 13416
rect 18874 13404 18880 13416
rect 18932 13404 18938 13456
rect 19150 13404 19156 13456
rect 19208 13444 19214 13456
rect 19208 13416 20024 13444
rect 19208 13404 19214 13416
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 15856 13348 18245 13376
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 18417 13379 18475 13385
rect 18417 13345 18429 13379
rect 18463 13376 18475 13379
rect 18506 13376 18512 13388
rect 18463 13348 18512 13376
rect 18463 13345 18475 13348
rect 18417 13339 18475 13345
rect 8234 13294 9076 13308
rect 8220 13280 9076 13294
rect 12805 13311 12863 13317
rect 6454 13132 6460 13184
rect 6512 13172 6518 13184
rect 8220 13172 8248 13280
rect 12805 13277 12817 13311
rect 12851 13308 12863 13311
rect 18248 13308 18276 13339
rect 18506 13336 18512 13348
rect 18564 13336 18570 13388
rect 19886 13336 19892 13388
rect 19944 13336 19950 13388
rect 19996 13385 20024 13416
rect 19981 13379 20039 13385
rect 19981 13345 19993 13379
rect 20027 13345 20039 13379
rect 19981 13339 20039 13345
rect 18785 13311 18843 13317
rect 18785 13308 18797 13311
rect 12851 13280 14596 13308
rect 18248 13280 18797 13308
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 11606 13240 11612 13252
rect 11362 13212 11612 13240
rect 11606 13200 11612 13212
rect 11664 13240 11670 13252
rect 11974 13240 11980 13252
rect 11664 13212 11980 13240
rect 11664 13200 11670 13212
rect 11974 13200 11980 13212
rect 12032 13200 12038 13252
rect 12713 13243 12771 13249
rect 12713 13209 12725 13243
rect 12759 13240 12771 13243
rect 14458 13240 14464 13252
rect 12759 13212 14464 13240
rect 12759 13209 12771 13212
rect 12713 13203 12771 13209
rect 14458 13200 14464 13212
rect 14516 13200 14522 13252
rect 6512 13144 8248 13172
rect 8573 13175 8631 13181
rect 6512 13132 6518 13144
rect 8573 13141 8585 13175
rect 8619 13172 8631 13175
rect 8754 13172 8760 13184
rect 8619 13144 8760 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 8754 13132 8760 13144
rect 8812 13132 8818 13184
rect 14568 13172 14596 13280
rect 18785 13277 18797 13280
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19797 13311 19855 13317
rect 19797 13308 19809 13311
rect 19484 13280 19809 13308
rect 19484 13268 19490 13280
rect 19797 13277 19809 13280
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 22646 13268 22652 13320
rect 22704 13268 22710 13320
rect 14826 13200 14832 13252
rect 14884 13200 14890 13252
rect 16482 13240 16488 13252
rect 16054 13212 16488 13240
rect 16482 13200 16488 13212
rect 16540 13200 16546 13252
rect 18141 13243 18199 13249
rect 18141 13209 18153 13243
rect 18187 13240 18199 13243
rect 18322 13240 18328 13252
rect 18187 13212 18328 13240
rect 18187 13209 18199 13212
rect 18141 13203 18199 13209
rect 18322 13200 18328 13212
rect 18380 13200 18386 13252
rect 23845 13243 23903 13249
rect 23845 13209 23857 13243
rect 23891 13240 23903 13243
rect 25682 13240 25688 13252
rect 23891 13212 25688 13240
rect 23891 13209 23903 13212
rect 23845 13203 23903 13209
rect 25682 13200 25688 13212
rect 25740 13200 25746 13252
rect 15470 13172 15476 13184
rect 14568 13144 15476 13172
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 16853 13175 16911 13181
rect 16853 13141 16865 13175
rect 16899 13172 16911 13175
rect 17218 13172 17224 13184
rect 16899 13144 17224 13172
rect 16899 13141 16911 13144
rect 16853 13135 16911 13141
rect 17218 13132 17224 13144
rect 17276 13132 17282 13184
rect 17770 13132 17776 13184
rect 17828 13132 17834 13184
rect 19429 13175 19487 13181
rect 19429 13141 19441 13175
rect 19475 13172 19487 13175
rect 19794 13172 19800 13184
rect 19475 13144 19800 13172
rect 19475 13141 19487 13144
rect 19429 13135 19487 13141
rect 19794 13132 19800 13144
rect 19852 13132 19858 13184
rect 21358 13132 21364 13184
rect 21416 13172 21422 13184
rect 21545 13175 21603 13181
rect 21545 13172 21557 13175
rect 21416 13144 21557 13172
rect 21416 13132 21422 13144
rect 21545 13141 21557 13144
rect 21591 13172 21603 13175
rect 22002 13172 22008 13184
rect 21591 13144 22008 13172
rect 21591 13141 21603 13144
rect 21545 13135 21603 13141
rect 22002 13132 22008 13144
rect 22060 13132 22066 13184
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 8662 12928 8668 12980
rect 8720 12928 8726 12980
rect 11149 12971 11207 12977
rect 11149 12937 11161 12971
rect 11195 12968 11207 12971
rect 11790 12968 11796 12980
rect 11195 12940 11796 12968
rect 11195 12937 11207 12940
rect 11149 12931 11207 12937
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 12710 12968 12716 12980
rect 12584 12940 12716 12968
rect 12584 12928 12590 12940
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 15746 12928 15752 12980
rect 15804 12968 15810 12980
rect 15841 12971 15899 12977
rect 15841 12968 15853 12971
rect 15804 12940 15853 12968
rect 15804 12928 15810 12940
rect 15841 12937 15853 12940
rect 15887 12937 15899 12971
rect 15841 12931 15899 12937
rect 16482 12928 16488 12980
rect 16540 12928 16546 12980
rect 17218 12928 17224 12980
rect 17276 12928 17282 12980
rect 18506 12928 18512 12980
rect 18564 12968 18570 12980
rect 21453 12971 21511 12977
rect 21453 12968 21465 12971
rect 18564 12940 21465 12968
rect 18564 12928 18570 12940
rect 21453 12937 21465 12940
rect 21499 12937 21511 12971
rect 21453 12931 21511 12937
rect 9674 12900 9680 12912
rect 9416 12872 9680 12900
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 9416 12841 9444 12872
rect 9674 12860 9680 12872
rect 9732 12900 9738 12912
rect 9950 12900 9956 12912
rect 9732 12872 9956 12900
rect 9732 12860 9738 12872
rect 9950 12860 9956 12872
rect 10008 12860 10014 12912
rect 11606 12900 11612 12912
rect 10902 12872 11612 12900
rect 11606 12860 11612 12872
rect 11664 12860 11670 12912
rect 14366 12860 14372 12912
rect 14424 12900 14430 12912
rect 14461 12903 14519 12909
rect 14461 12900 14473 12903
rect 14424 12872 14473 12900
rect 14424 12860 14430 12872
rect 14461 12869 14473 12872
rect 14507 12900 14519 12903
rect 14921 12903 14979 12909
rect 14921 12900 14933 12903
rect 14507 12872 14933 12900
rect 14507 12869 14519 12872
rect 14461 12863 14519 12869
rect 14921 12869 14933 12872
rect 14967 12869 14979 12903
rect 14921 12863 14979 12869
rect 15381 12903 15439 12909
rect 15381 12869 15393 12903
rect 15427 12900 15439 12903
rect 15764 12900 15792 12928
rect 15427 12872 15792 12900
rect 15427 12869 15439 12872
rect 15381 12863 15439 12869
rect 17034 12860 17040 12912
rect 17092 12900 17098 12912
rect 17313 12903 17371 12909
rect 17313 12900 17325 12903
rect 17092 12872 17325 12900
rect 17092 12860 17098 12872
rect 17313 12869 17325 12872
rect 17359 12869 17371 12903
rect 17313 12863 17371 12869
rect 18874 12860 18880 12912
rect 18932 12900 18938 12912
rect 18969 12903 19027 12909
rect 18969 12900 18981 12903
rect 18932 12872 18981 12900
rect 18932 12860 18938 12872
rect 18969 12869 18981 12872
rect 19015 12869 19027 12903
rect 21358 12900 21364 12912
rect 21206 12872 21364 12900
rect 18969 12863 19027 12869
rect 21358 12860 21364 12872
rect 21416 12860 21422 12912
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 6604 12804 8585 12832
rect 6604 12792 6610 12804
rect 8573 12801 8585 12804
rect 8619 12801 8631 12835
rect 8573 12795 8631 12801
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 13688 12804 13737 12832
rect 13688 12792 13694 12804
rect 13725 12801 13737 12804
rect 13771 12832 13783 12835
rect 13814 12832 13820 12844
rect 13771 12804 13820 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 15930 12792 15936 12844
rect 15988 12832 15994 12844
rect 18509 12835 18567 12841
rect 15988 12804 17448 12832
rect 15988 12792 15994 12804
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 17420 12773 17448 12804
rect 18509 12801 18521 12835
rect 18555 12832 18567 12835
rect 18892 12832 18920 12860
rect 18555 12804 18920 12832
rect 18555 12801 18567 12804
rect 18509 12795 18567 12801
rect 22830 12792 22836 12844
rect 22888 12792 22894 12844
rect 23290 12792 23296 12844
rect 23348 12832 23354 12844
rect 23937 12835 23995 12841
rect 23937 12832 23949 12835
rect 23348 12804 23949 12832
rect 23348 12792 23354 12804
rect 23937 12801 23949 12804
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 9677 12767 9735 12773
rect 9677 12764 9689 12767
rect 8812 12736 9689 12764
rect 8812 12724 8818 12736
rect 9677 12733 9689 12736
rect 9723 12733 9735 12767
rect 9677 12727 9735 12733
rect 17405 12767 17463 12773
rect 17405 12733 17417 12767
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 19518 12724 19524 12776
rect 19576 12764 19582 12776
rect 19705 12767 19763 12773
rect 19705 12764 19717 12767
rect 19576 12736 19717 12764
rect 19576 12724 19582 12736
rect 19705 12733 19717 12736
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12764 20039 12767
rect 21818 12764 21824 12776
rect 20027 12736 21824 12764
rect 20027 12733 20039 12736
rect 19981 12727 20039 12733
rect 21818 12724 21824 12736
rect 21876 12724 21882 12776
rect 22002 12724 22008 12776
rect 22060 12724 22066 12776
rect 24762 12724 24768 12776
rect 24820 12724 24826 12776
rect 13909 12699 13967 12705
rect 13909 12665 13921 12699
rect 13955 12696 13967 12699
rect 14366 12696 14372 12708
rect 13955 12668 14372 12696
rect 13955 12665 13967 12668
rect 13909 12659 13967 12665
rect 14366 12656 14372 12668
rect 14424 12656 14430 12708
rect 14642 12656 14648 12708
rect 14700 12656 14706 12708
rect 15565 12699 15623 12705
rect 15565 12665 15577 12699
rect 15611 12696 15623 12699
rect 16206 12696 16212 12708
rect 15611 12668 16212 12696
rect 15611 12665 15623 12668
rect 15565 12659 15623 12665
rect 16206 12656 16212 12668
rect 16264 12656 16270 12708
rect 8205 12631 8263 12637
rect 8205 12597 8217 12631
rect 8251 12628 8263 12631
rect 10962 12628 10968 12640
rect 8251 12600 10968 12628
rect 8251 12597 8263 12600
rect 8205 12591 8263 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 16853 12631 16911 12637
rect 16853 12597 16865 12631
rect 16899 12628 16911 12631
rect 17678 12628 17684 12640
rect 16899 12600 17684 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 17678 12588 17684 12600
rect 17736 12588 17742 12640
rect 18598 12588 18604 12640
rect 18656 12588 18662 12640
rect 22649 12631 22707 12637
rect 22649 12597 22661 12631
rect 22695 12628 22707 12631
rect 24578 12628 24584 12640
rect 22695 12600 24584 12628
rect 22695 12597 22707 12600
rect 22649 12591 22707 12597
rect 24578 12588 24584 12600
rect 24636 12588 24642 12640
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 8938 12384 8944 12436
rect 8996 12424 9002 12436
rect 10134 12424 10140 12436
rect 8996 12396 10140 12424
rect 8996 12384 9002 12396
rect 10134 12384 10140 12396
rect 10192 12384 10198 12436
rect 12158 12384 12164 12436
rect 12216 12424 12222 12436
rect 12342 12424 12348 12436
rect 12216 12396 12348 12424
rect 12216 12384 12222 12396
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 13872 12396 14105 12424
rect 13872 12384 13878 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 14093 12387 14151 12393
rect 14458 12384 14464 12436
rect 14516 12384 14522 12436
rect 15654 12384 15660 12436
rect 15712 12384 15718 12436
rect 17402 12424 17408 12436
rect 16040 12396 17408 12424
rect 11790 12248 11796 12300
rect 11848 12248 11854 12300
rect 13998 12248 14004 12300
rect 14056 12288 14062 12300
rect 15105 12291 15163 12297
rect 15105 12288 15117 12291
rect 14056 12260 15117 12288
rect 14056 12248 14062 12260
rect 15105 12257 15117 12260
rect 15151 12288 15163 12291
rect 15654 12288 15660 12300
rect 15151 12260 15660 12288
rect 15151 12257 15163 12260
rect 15105 12251 15163 12257
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 11514 12220 11520 12232
rect 9732 12192 11520 12220
rect 9732 12180 9738 12192
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 16040 12229 16068 12396
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 17494 12384 17500 12436
rect 17552 12424 17558 12436
rect 18877 12427 18935 12433
rect 18877 12424 18889 12427
rect 17552 12396 18889 12424
rect 17552 12384 17558 12396
rect 18877 12393 18889 12396
rect 18923 12393 18935 12427
rect 18877 12387 18935 12393
rect 20441 12359 20499 12365
rect 20441 12325 20453 12359
rect 20487 12356 20499 12359
rect 23290 12356 23296 12368
rect 20487 12328 23296 12356
rect 20487 12325 20499 12328
rect 20441 12319 20499 12325
rect 23290 12316 23296 12328
rect 23348 12316 23354 12368
rect 16114 12248 16120 12300
rect 16172 12288 16178 12300
rect 16209 12291 16267 12297
rect 16209 12288 16221 12291
rect 16172 12260 16221 12288
rect 16172 12248 16178 12260
rect 16209 12257 16221 12260
rect 16255 12257 16267 12291
rect 16209 12251 16267 12257
rect 17126 12248 17132 12300
rect 17184 12248 17190 12300
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12288 17463 12291
rect 19978 12288 19984 12300
rect 17451 12260 19984 12288
rect 17451 12257 17463 12260
rect 17405 12251 17463 12257
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 21266 12248 21272 12300
rect 21324 12288 21330 12300
rect 21545 12291 21603 12297
rect 21545 12288 21557 12291
rect 21324 12260 21557 12288
rect 21324 12248 21330 12260
rect 21545 12257 21557 12260
rect 21591 12257 21603 12291
rect 21545 12251 21603 12257
rect 21729 12291 21787 12297
rect 21729 12257 21741 12291
rect 21775 12288 21787 12291
rect 21818 12288 21824 12300
rect 21775 12260 21824 12288
rect 21775 12257 21787 12260
rect 21729 12251 21787 12257
rect 21818 12248 21824 12260
rect 21876 12248 21882 12300
rect 21910 12248 21916 12300
rect 21968 12288 21974 12300
rect 21968 12260 23428 12288
rect 21968 12248 21974 12260
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 19334 12180 19340 12232
rect 19392 12220 19398 12232
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 19392 12192 20637 12220
rect 19392 12180 19398 12192
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 21453 12223 21511 12229
rect 21453 12189 21465 12223
rect 21499 12220 21511 12223
rect 22002 12220 22008 12232
rect 21499 12192 22008 12220
rect 21499 12189 21511 12192
rect 21453 12183 21511 12189
rect 22002 12180 22008 12192
rect 22060 12180 22066 12232
rect 23400 12229 23428 12260
rect 23385 12223 23443 12229
rect 23385 12189 23397 12223
rect 23431 12189 23443 12223
rect 23385 12183 23443 12189
rect 10226 12112 10232 12164
rect 10284 12152 10290 12164
rect 12066 12152 12072 12164
rect 10284 12124 12072 12152
rect 10284 12112 10290 12124
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 13633 12155 13691 12161
rect 13633 12152 13645 12155
rect 13018 12124 13645 12152
rect 13633 12121 13645 12124
rect 13679 12152 13691 12155
rect 14182 12152 14188 12164
rect 13679 12124 14188 12152
rect 13679 12121 13691 12124
rect 13633 12115 13691 12121
rect 14182 12112 14188 12124
rect 14240 12112 14246 12164
rect 14829 12155 14887 12161
rect 14829 12121 14841 12155
rect 14875 12152 14887 12155
rect 17310 12152 17316 12164
rect 14875 12124 17316 12152
rect 14875 12121 14887 12124
rect 14829 12115 14887 12121
rect 17310 12112 17316 12124
rect 17368 12112 17374 12164
rect 18630 12124 18736 12152
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 9582 12084 9588 12096
rect 3568 12056 9588 12084
rect 3568 12044 3574 12056
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 13228 12056 13277 12084
rect 13228 12044 13234 12056
rect 13265 12053 13277 12056
rect 13311 12053 13323 12087
rect 13265 12047 13323 12053
rect 13909 12087 13967 12093
rect 13909 12053 13921 12087
rect 13955 12084 13967 12087
rect 14918 12084 14924 12096
rect 13955 12056 14924 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 14918 12044 14924 12056
rect 14976 12084 14982 12096
rect 15286 12084 15292 12096
rect 14976 12056 15292 12084
rect 14976 12044 14982 12056
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 15378 12044 15384 12096
rect 15436 12084 15442 12096
rect 16117 12087 16175 12093
rect 16117 12084 16129 12087
rect 15436 12056 16129 12084
rect 15436 12044 15442 12056
rect 16117 12053 16129 12056
rect 16163 12084 16175 12087
rect 18322 12084 18328 12096
rect 16163 12056 18328 12084
rect 16163 12053 16175 12056
rect 16117 12047 16175 12053
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 18708 12084 18736 12124
rect 19337 12087 19395 12093
rect 19337 12084 19349 12087
rect 18708 12056 19349 12084
rect 19337 12053 19349 12056
rect 19383 12084 19395 12087
rect 19886 12084 19892 12096
rect 19383 12056 19892 12084
rect 19383 12053 19395 12056
rect 19337 12047 19395 12053
rect 19886 12044 19892 12056
rect 19944 12044 19950 12096
rect 21082 12044 21088 12096
rect 21140 12044 21146 12096
rect 23201 12087 23259 12093
rect 23201 12053 23213 12087
rect 23247 12084 23259 12087
rect 24854 12084 24860 12096
rect 23247 12056 24860 12084
rect 23247 12053 23259 12056
rect 23201 12047 23259 12053
rect 24854 12044 24860 12056
rect 24912 12044 24918 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 12400 11852 14412 11880
rect 12400 11840 12406 11852
rect 5166 11772 5172 11824
rect 5224 11812 5230 11824
rect 10686 11812 10692 11824
rect 5224 11784 10692 11812
rect 5224 11772 5230 11784
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 14384 11812 14412 11852
rect 14550 11840 14556 11892
rect 14608 11840 14614 11892
rect 16117 11883 16175 11889
rect 16117 11849 16129 11883
rect 16163 11880 16175 11883
rect 16482 11880 16488 11892
rect 16163 11852 16488 11880
rect 16163 11849 16175 11852
rect 16117 11843 16175 11849
rect 15473 11815 15531 11821
rect 15473 11812 15485 11815
rect 14384 11784 15485 11812
rect 15473 11781 15485 11784
rect 15519 11781 15531 11815
rect 15473 11775 15531 11781
rect 11514 11704 11520 11756
rect 11572 11744 11578 11756
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 11572 11716 12817 11744
rect 11572 11704 11578 11716
rect 12805 11713 12817 11716
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 14182 11704 14188 11756
rect 14240 11704 14246 11756
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 14792 11716 15393 11744
rect 14792 11704 14798 11716
rect 15381 11713 15393 11716
rect 15427 11713 15439 11747
rect 16132 11744 16160 11843
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 17494 11840 17500 11892
rect 17552 11840 17558 11892
rect 19518 11880 19524 11892
rect 18248 11852 19524 11880
rect 16945 11815 17003 11821
rect 16945 11781 16957 11815
rect 16991 11812 17003 11815
rect 17512 11812 17540 11840
rect 16991 11784 17540 11812
rect 16991 11781 17003 11784
rect 16945 11775 17003 11781
rect 18248 11753 18276 11852
rect 19518 11840 19524 11852
rect 19576 11840 19582 11892
rect 19978 11840 19984 11892
rect 20036 11840 20042 11892
rect 18506 11772 18512 11824
rect 18564 11772 18570 11824
rect 20714 11772 20720 11824
rect 20772 11812 20778 11824
rect 20901 11815 20959 11821
rect 20901 11812 20913 11815
rect 20772 11784 20913 11812
rect 20772 11772 20778 11784
rect 20901 11781 20913 11784
rect 20947 11812 20959 11815
rect 21361 11815 21419 11821
rect 21361 11812 21373 11815
rect 20947 11784 21373 11812
rect 20947 11781 20959 11784
rect 20901 11775 20959 11781
rect 21361 11781 21373 11784
rect 21407 11781 21419 11815
rect 21361 11775 21419 11781
rect 25130 11772 25136 11824
rect 25188 11772 25194 11824
rect 15381 11707 15439 11713
rect 15488 11716 16160 11744
rect 18233 11747 18291 11753
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11676 13139 11679
rect 13170 11676 13176 11688
rect 13127 11648 13176 11676
rect 13127 11645 13139 11648
rect 13081 11639 13139 11645
rect 13170 11636 13176 11648
rect 13228 11676 13234 11688
rect 14200 11676 14228 11704
rect 15488 11676 15516 11716
rect 18233 11713 18245 11747
rect 18279 11713 18291 11747
rect 19886 11744 19892 11756
rect 19642 11716 19892 11744
rect 18233 11707 18291 11713
rect 19886 11704 19892 11716
rect 19944 11744 19950 11756
rect 19944 11716 20576 11744
rect 19944 11704 19950 11716
rect 13228 11648 14136 11676
rect 14200 11648 15516 11676
rect 15565 11679 15623 11685
rect 13228 11636 13234 11648
rect 14108 11608 14136 11648
rect 15565 11645 15577 11679
rect 15611 11645 15623 11679
rect 15565 11639 15623 11645
rect 15580 11608 15608 11639
rect 17402 11636 17408 11688
rect 17460 11676 17466 11688
rect 20438 11676 20444 11688
rect 17460 11648 20444 11676
rect 17460 11636 17466 11648
rect 20438 11636 20444 11648
rect 20496 11636 20502 11688
rect 14108 11580 15608 11608
rect 15013 11543 15071 11549
rect 15013 11509 15025 11543
rect 15059 11540 15071 11543
rect 15746 11540 15752 11552
rect 15059 11512 15752 11540
rect 15059 11509 15071 11512
rect 15013 11503 15071 11509
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 17037 11543 17095 11549
rect 17037 11540 17049 11543
rect 16816 11512 17049 11540
rect 16816 11500 16822 11512
rect 17037 11509 17049 11512
rect 17083 11509 17095 11543
rect 17037 11503 17095 11509
rect 20349 11543 20407 11549
rect 20349 11509 20361 11543
rect 20395 11540 20407 11543
rect 20548 11540 20576 11716
rect 22554 11704 22560 11756
rect 22612 11744 22618 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 22612 11716 23949 11744
rect 22612 11704 22618 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 21085 11611 21143 11617
rect 21085 11577 21097 11611
rect 21131 11608 21143 11611
rect 22094 11608 22100 11620
rect 21131 11580 22100 11608
rect 21131 11577 21143 11580
rect 21085 11571 21143 11577
rect 22094 11568 22100 11580
rect 22152 11568 22158 11620
rect 21358 11540 21364 11552
rect 20395 11512 21364 11540
rect 20395 11509 20407 11512
rect 20349 11503 20407 11509
rect 21358 11500 21364 11512
rect 21416 11540 21422 11552
rect 24486 11540 24492 11552
rect 21416 11512 24492 11540
rect 21416 11500 21422 11512
rect 24486 11500 24492 11512
rect 24544 11500 24550 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 15470 11296 15476 11348
rect 15528 11296 15534 11348
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 16850 11336 16856 11348
rect 16724 11308 16856 11336
rect 16724 11296 16730 11308
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 14734 11160 14740 11212
rect 14792 11160 14798 11212
rect 15654 11160 15660 11212
rect 15712 11200 15718 11212
rect 16025 11203 16083 11209
rect 16025 11200 16037 11203
rect 15712 11172 16037 11200
rect 15712 11160 15718 11172
rect 16025 11169 16037 11172
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 15930 11092 15936 11144
rect 15988 11132 15994 11144
rect 17586 11132 17592 11144
rect 15988 11104 17592 11132
rect 15988 11092 15994 11104
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 15841 11067 15899 11073
rect 15841 11033 15853 11067
rect 15887 11064 15899 11067
rect 20622 11064 20628 11076
rect 15887 11036 20628 11064
rect 15887 11033 15899 11036
rect 15841 11027 15899 11033
rect 20622 11024 20628 11036
rect 20680 11024 20686 11076
rect 20806 11024 20812 11076
rect 20864 11024 20870 11076
rect 20993 11067 21051 11073
rect 20993 11033 21005 11067
rect 21039 11064 21051 11067
rect 23842 11064 23848 11076
rect 21039 11036 23848 11064
rect 21039 11033 21051 11036
rect 20993 11027 21051 11033
rect 23842 11024 23848 11036
rect 23900 11024 23906 11076
rect 19610 10956 19616 11008
rect 19668 10956 19674 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 19521 10795 19579 10801
rect 19521 10761 19533 10795
rect 19567 10792 19579 10795
rect 19610 10792 19616 10804
rect 19567 10764 19616 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 19610 10752 19616 10764
rect 19668 10752 19674 10804
rect 20349 10795 20407 10801
rect 20349 10761 20361 10795
rect 20395 10761 20407 10795
rect 20349 10755 20407 10761
rect 10962 10684 10968 10736
rect 11020 10724 11026 10736
rect 11020 10696 14872 10724
rect 11020 10684 11026 10696
rect 12066 10616 12072 10668
rect 12124 10616 12130 10668
rect 14844 10665 14872 10696
rect 17678 10684 17684 10736
rect 17736 10724 17742 10736
rect 20364 10724 20392 10755
rect 17736 10696 18736 10724
rect 20364 10696 23428 10724
rect 17736 10684 17742 10696
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10625 14887 10659
rect 14829 10619 14887 10625
rect 15746 10616 15752 10668
rect 15804 10656 15810 10668
rect 18417 10659 18475 10665
rect 18417 10656 18429 10659
rect 15804 10628 18429 10656
rect 15804 10616 15810 10628
rect 18417 10625 18429 10628
rect 18463 10625 18475 10659
rect 18708 10656 18736 10696
rect 23400 10665 23428 10696
rect 20533 10659 20591 10665
rect 20533 10656 20545 10659
rect 18708 10628 20545 10656
rect 18417 10619 18475 10625
rect 20533 10625 20545 10628
rect 20579 10625 20591 10659
rect 20533 10619 20591 10625
rect 23385 10659 23443 10665
rect 23385 10625 23397 10659
rect 23431 10625 23443 10659
rect 23385 10619 23443 10625
rect 23937 10659 23995 10665
rect 23937 10625 23949 10659
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 17770 10548 17776 10600
rect 17828 10588 17834 10600
rect 19613 10591 19671 10597
rect 19613 10588 19625 10591
rect 17828 10560 19625 10588
rect 17828 10548 17834 10560
rect 19613 10557 19625 10560
rect 19659 10557 19671 10591
rect 19613 10551 19671 10557
rect 19797 10591 19855 10597
rect 19797 10557 19809 10591
rect 19843 10588 19855 10591
rect 19978 10588 19984 10600
rect 19843 10560 19984 10588
rect 19843 10557 19855 10560
rect 19797 10551 19855 10557
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 21542 10548 21548 10600
rect 21600 10588 21606 10600
rect 23952 10588 23980 10619
rect 21600 10560 23980 10588
rect 21600 10548 21606 10560
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 12253 10523 12311 10529
rect 12253 10489 12265 10523
rect 12299 10520 12311 10523
rect 12526 10520 12532 10532
rect 12299 10492 12532 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 14645 10523 14703 10529
rect 14645 10489 14657 10523
rect 14691 10520 14703 10523
rect 20806 10520 20812 10532
rect 14691 10492 20812 10520
rect 14691 10489 14703 10492
rect 14645 10483 14703 10489
rect 20806 10480 20812 10492
rect 20864 10480 20870 10532
rect 5258 10412 5264 10464
rect 5316 10452 5322 10464
rect 9858 10452 9864 10464
rect 5316 10424 9864 10452
rect 5316 10412 5322 10424
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 18230 10412 18236 10464
rect 18288 10412 18294 10464
rect 19153 10455 19211 10461
rect 19153 10421 19165 10455
rect 19199 10452 19211 10455
rect 21726 10452 21732 10464
rect 19199 10424 21732 10452
rect 19199 10421 19211 10424
rect 19153 10415 19211 10421
rect 21726 10412 21732 10424
rect 21784 10412 21790 10464
rect 23201 10455 23259 10461
rect 23201 10421 23213 10455
rect 23247 10452 23259 10455
rect 23934 10452 23940 10464
rect 23247 10424 23940 10452
rect 23247 10421 23259 10424
rect 23201 10415 23259 10421
rect 23934 10412 23940 10424
rect 23992 10412 23998 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 21269 10183 21327 10189
rect 21269 10149 21281 10183
rect 21315 10180 21327 10183
rect 22554 10180 22560 10192
rect 21315 10152 22560 10180
rect 21315 10149 21327 10152
rect 21269 10143 21327 10149
rect 22554 10140 22560 10152
rect 22612 10140 22618 10192
rect 18230 10072 18236 10124
rect 18288 10112 18294 10124
rect 18288 10084 22232 10112
rect 18288 10072 18294 10084
rect 13630 10004 13636 10056
rect 13688 10044 13694 10056
rect 14645 10047 14703 10053
rect 14645 10044 14657 10047
rect 13688 10016 14657 10044
rect 13688 10004 13694 10016
rect 14645 10013 14657 10016
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 14829 10047 14887 10053
rect 14829 10013 14841 10047
rect 14875 10044 14887 10047
rect 19426 10044 19432 10056
rect 14875 10016 19432 10044
rect 14875 10013 14887 10016
rect 14829 10007 14887 10013
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 19794 10004 19800 10056
rect 19852 10044 19858 10056
rect 22204 10053 22232 10084
rect 21453 10047 21511 10053
rect 21453 10044 21465 10047
rect 19852 10016 21465 10044
rect 19852 10004 19858 10016
rect 21453 10013 21465 10016
rect 21499 10013 21511 10047
rect 21453 10007 21511 10013
rect 22189 10047 22247 10053
rect 22189 10013 22201 10047
rect 22235 10013 22247 10047
rect 22189 10007 22247 10013
rect 22649 10047 22707 10053
rect 22649 10013 22661 10047
rect 22695 10013 22707 10047
rect 22649 10007 22707 10013
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10044 23903 10047
rect 24946 10044 24952 10056
rect 23891 10016 24952 10044
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 16761 9979 16819 9985
rect 16761 9945 16773 9979
rect 16807 9976 16819 9979
rect 18414 9976 18420 9988
rect 16807 9948 18420 9976
rect 16807 9945 16819 9948
rect 16761 9939 16819 9945
rect 18414 9936 18420 9948
rect 18472 9936 18478 9988
rect 22664 9976 22692 10007
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 22020 9948 22692 9976
rect 16850 9868 16856 9920
rect 16908 9868 16914 9920
rect 22020 9917 22048 9948
rect 23290 9936 23296 9988
rect 23348 9976 23354 9988
rect 24673 9979 24731 9985
rect 24673 9976 24685 9979
rect 23348 9948 24685 9976
rect 23348 9936 23354 9948
rect 24673 9945 24685 9948
rect 24719 9945 24731 9979
rect 24673 9939 24731 9945
rect 22005 9911 22063 9917
rect 22005 9877 22017 9911
rect 22051 9877 22063 9911
rect 22005 9871 22063 9877
rect 24026 9868 24032 9920
rect 24084 9908 24090 9920
rect 24765 9911 24823 9917
rect 24765 9908 24777 9911
rect 24084 9880 24777 9908
rect 24084 9868 24090 9880
rect 24765 9877 24777 9880
rect 24811 9877 24823 9911
rect 24765 9871 24823 9877
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 9490 9596 9496 9648
rect 9548 9636 9554 9648
rect 13906 9636 13912 9648
rect 9548 9608 13912 9636
rect 9548 9596 9554 9608
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 15562 9596 15568 9648
rect 15620 9636 15626 9648
rect 16945 9639 17003 9645
rect 16945 9636 16957 9639
rect 15620 9608 16957 9636
rect 15620 9596 15626 9608
rect 16945 9605 16957 9608
rect 16991 9605 17003 9639
rect 16945 9599 17003 9605
rect 18690 9596 18696 9648
rect 18748 9636 18754 9648
rect 19061 9639 19119 9645
rect 19061 9636 19073 9639
rect 18748 9608 19073 9636
rect 18748 9596 18754 9608
rect 19061 9605 19073 9608
rect 19107 9605 19119 9639
rect 19061 9599 19119 9605
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 5859 9540 6929 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 21082 9528 21088 9580
rect 21140 9568 21146 9580
rect 22925 9571 22983 9577
rect 22925 9568 22937 9571
rect 21140 9540 22937 9568
rect 21140 9528 21146 9540
rect 22925 9537 22937 9540
rect 22971 9537 22983 9571
rect 22925 9531 22983 9537
rect 23842 9528 23848 9580
rect 23900 9568 23906 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 23900 9540 23949 9568
rect 23900 9528 23906 9540
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 5592 9472 7021 9500
rect 5592 9460 5598 9472
rect 7009 9469 7021 9472
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 7098 9460 7104 9512
rect 7156 9460 7162 9512
rect 24670 9460 24676 9512
rect 24728 9460 24734 9512
rect 6546 9392 6552 9444
rect 6604 9392 6610 9444
rect 17129 9435 17187 9441
rect 17129 9401 17141 9435
rect 17175 9432 17187 9435
rect 17678 9432 17684 9444
rect 17175 9404 17684 9432
rect 17175 9401 17187 9404
rect 17129 9395 17187 9401
rect 17678 9392 17684 9404
rect 17736 9392 17742 9444
rect 19245 9435 19303 9441
rect 19245 9401 19257 9435
rect 19291 9432 19303 9435
rect 23842 9432 23848 9444
rect 19291 9404 23848 9432
rect 19291 9401 19303 9404
rect 19245 9395 19303 9401
rect 23842 9392 23848 9404
rect 23900 9392 23906 9444
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 11698 9364 11704 9376
rect 7156 9336 11704 9364
rect 7156 9324 7162 9336
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 22738 9324 22744 9376
rect 22796 9324 22802 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 3050 9120 3056 9172
rect 3108 9160 3114 9172
rect 5902 9160 5908 9172
rect 3108 9132 5908 9160
rect 3108 9120 3114 9132
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 22830 9052 22836 9104
rect 22888 9092 22894 9104
rect 24673 9095 24731 9101
rect 24673 9092 24685 9095
rect 22888 9064 24685 9092
rect 22888 9052 22894 9064
rect 24673 9061 24685 9064
rect 24719 9061 24731 9095
rect 24673 9055 24731 9061
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 15010 8956 15016 8968
rect 7800 8928 15016 8956
rect 7800 8916 7806 8928
rect 15010 8916 15016 8928
rect 15068 8916 15074 8968
rect 21726 8916 21732 8968
rect 21784 8916 21790 8968
rect 23382 8916 23388 8968
rect 23440 8956 23446 8968
rect 23937 8959 23995 8965
rect 23937 8956 23949 8959
rect 23440 8928 23949 8956
rect 23440 8916 23446 8928
rect 23937 8925 23949 8928
rect 23983 8925 23995 8959
rect 23937 8919 23995 8925
rect 24578 8916 24584 8968
rect 24636 8956 24642 8968
rect 24857 8959 24915 8965
rect 24857 8956 24869 8959
rect 24636 8928 24869 8956
rect 24636 8916 24642 8928
rect 24857 8925 24869 8928
rect 24903 8925 24915 8959
rect 24857 8919 24915 8925
rect 21545 8823 21603 8829
rect 21545 8789 21557 8823
rect 21591 8820 21603 8823
rect 23290 8820 23296 8832
rect 21591 8792 23296 8820
rect 21591 8789 21603 8792
rect 21545 8783 21603 8789
rect 23290 8780 23296 8792
rect 23348 8780 23354 8832
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 23753 8823 23811 8829
rect 23753 8820 23765 8823
rect 23532 8792 23765 8820
rect 23532 8780 23538 8792
rect 23753 8789 23765 8792
rect 23799 8789 23811 8823
rect 23753 8783 23811 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 18874 8508 18880 8560
rect 18932 8548 18938 8560
rect 19153 8551 19211 8557
rect 19153 8548 19165 8551
rect 18932 8520 19165 8548
rect 18932 8508 18938 8520
rect 19153 8517 19165 8520
rect 19199 8517 19211 8551
rect 19153 8511 19211 8517
rect 20717 8551 20775 8557
rect 20717 8517 20729 8551
rect 20763 8548 20775 8551
rect 20898 8548 20904 8560
rect 20763 8520 20904 8548
rect 20763 8517 20775 8520
rect 20717 8511 20775 8517
rect 20898 8508 20904 8520
rect 20956 8508 20962 8560
rect 25130 8508 25136 8560
rect 25188 8508 25194 8560
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8480 22339 8483
rect 22327 8452 23520 8480
rect 22327 8449 22339 8452
rect 22281 8443 22339 8449
rect 20901 8415 20959 8421
rect 20901 8381 20913 8415
rect 20947 8412 20959 8415
rect 21266 8412 21272 8424
rect 20947 8384 21272 8412
rect 20947 8381 20959 8384
rect 20901 8375 20959 8381
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 22370 8372 22376 8424
rect 22428 8412 22434 8424
rect 22557 8415 22615 8421
rect 22557 8412 22569 8415
rect 22428 8384 22569 8412
rect 22428 8372 22434 8384
rect 22557 8381 22569 8384
rect 22603 8381 22615 8415
rect 23492 8412 23520 8452
rect 23934 8440 23940 8492
rect 23992 8440 23998 8492
rect 24946 8412 24952 8424
rect 23492 8384 24952 8412
rect 22557 8375 22615 8381
rect 24946 8372 24952 8384
rect 25004 8372 25010 8424
rect 11606 8304 11612 8356
rect 11664 8344 11670 8356
rect 18414 8344 18420 8356
rect 11664 8316 18420 8344
rect 11664 8304 11670 8316
rect 18414 8304 18420 8316
rect 18472 8304 18478 8356
rect 19337 8347 19395 8353
rect 19337 8313 19349 8347
rect 19383 8344 19395 8347
rect 22002 8344 22008 8356
rect 19383 8316 22008 8344
rect 19383 8313 19395 8316
rect 19337 8307 19395 8313
rect 22002 8304 22008 8316
rect 22060 8304 22066 8356
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 6454 8032 6460 8084
rect 6512 8032 6518 8084
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 12710 8072 12716 8084
rect 11940 8044 12716 8072
rect 11940 8032 11946 8044
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 6822 7936 6828 7948
rect 4111 7908 6828 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 23382 7896 23388 7948
rect 23440 7896 23446 7948
rect 6454 7868 6460 7880
rect 5474 7840 6460 7868
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 20438 7828 20444 7880
rect 20496 7828 20502 7880
rect 20622 7828 20628 7880
rect 20680 7868 20686 7880
rect 21269 7871 21327 7877
rect 21269 7868 21281 7871
rect 20680 7840 21281 7868
rect 20680 7828 20686 7840
rect 21269 7837 21281 7840
rect 21315 7837 21327 7871
rect 21269 7831 21327 7837
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7868 22891 7871
rect 23474 7868 23480 7880
rect 22879 7840 23480 7868
rect 22879 7837 22891 7840
rect 22833 7831 22891 7837
rect 23474 7828 23480 7840
rect 23532 7828 23538 7880
rect 24854 7828 24860 7880
rect 24912 7828 24918 7880
rect 2774 7760 2780 7812
rect 2832 7800 2838 7812
rect 4341 7803 4399 7809
rect 4341 7800 4353 7803
rect 2832 7772 4353 7800
rect 2832 7760 2838 7772
rect 4341 7769 4353 7772
rect 4387 7769 4399 7803
rect 4341 7763 4399 7769
rect 6089 7803 6147 7809
rect 6089 7769 6101 7803
rect 6135 7800 6147 7803
rect 9122 7800 9128 7812
rect 6135 7772 9128 7800
rect 6135 7769 6147 7772
rect 6089 7763 6147 7769
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 20257 7735 20315 7741
rect 20257 7701 20269 7735
rect 20303 7732 20315 7735
rect 20806 7732 20812 7744
rect 20303 7704 20812 7732
rect 20303 7701 20315 7704
rect 20257 7695 20315 7701
rect 20806 7692 20812 7704
rect 20864 7692 20870 7744
rect 21082 7692 21088 7744
rect 21140 7692 21146 7744
rect 24118 7692 24124 7744
rect 24176 7732 24182 7744
rect 24673 7735 24731 7741
rect 24673 7732 24685 7735
rect 24176 7704 24685 7732
rect 24176 7692 24182 7704
rect 24673 7701 24685 7704
rect 24719 7701 24731 7735
rect 24673 7695 24731 7701
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 17310 7420 17316 7472
rect 17368 7460 17374 7472
rect 18785 7463 18843 7469
rect 18785 7460 18797 7463
rect 17368 7432 18797 7460
rect 17368 7420 17374 7432
rect 18785 7429 18797 7432
rect 18831 7429 18843 7463
rect 18785 7423 18843 7429
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20898 7392 20904 7404
rect 20303 7364 20904 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 22002 7352 22008 7404
rect 22060 7392 22066 7404
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 22060 7364 22109 7392
rect 22060 7352 22066 7364
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 23934 7352 23940 7404
rect 23992 7352 23998 7404
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 22186 7324 22192 7336
rect 21315 7296 22192 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 22186 7284 22192 7296
rect 22244 7284 22250 7336
rect 22278 7284 22284 7336
rect 22336 7324 22342 7336
rect 22557 7327 22615 7333
rect 22557 7324 22569 7327
rect 22336 7296 22569 7324
rect 22336 7284 22342 7296
rect 22557 7293 22569 7296
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 18969 7259 19027 7265
rect 18969 7225 18981 7259
rect 19015 7256 19027 7259
rect 20622 7256 20628 7268
rect 19015 7228 20628 7256
rect 19015 7225 19027 7228
rect 18969 7219 19027 7225
rect 20622 7216 20628 7228
rect 20680 7216 20686 7268
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 16482 6740 16488 6792
rect 16540 6780 16546 6792
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 16540 6752 19717 6780
rect 16540 6740 16546 6752
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 20806 6740 20812 6792
rect 20864 6740 20870 6792
rect 22830 6740 22836 6792
rect 22888 6740 22894 6792
rect 3050 6672 3056 6724
rect 3108 6712 3114 6724
rect 5994 6712 6000 6724
rect 3108 6684 6000 6712
rect 3108 6672 3114 6684
rect 5994 6672 6000 6684
rect 6052 6672 6058 6724
rect 22002 6672 22008 6724
rect 22060 6672 22066 6724
rect 23845 6715 23903 6721
rect 23845 6681 23857 6715
rect 23891 6712 23903 6715
rect 24946 6712 24952 6724
rect 23891 6684 24952 6712
rect 23891 6681 23903 6684
rect 23845 6675 23903 6681
rect 24946 6672 24952 6684
rect 25004 6672 25010 6724
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 19521 6647 19579 6653
rect 19521 6644 19533 6647
rect 18564 6616 19533 6644
rect 18564 6604 18570 6616
rect 19521 6613 19533 6616
rect 19567 6613 19579 6647
rect 19521 6607 19579 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 11238 6332 11244 6384
rect 11296 6372 11302 6384
rect 16390 6372 16396 6384
rect 11296 6344 16396 6372
rect 11296 6332 11302 6344
rect 16390 6332 16396 6344
rect 16448 6332 16454 6384
rect 21269 6375 21327 6381
rect 21269 6341 21281 6375
rect 21315 6372 21327 6375
rect 22646 6372 22652 6384
rect 21315 6344 22652 6372
rect 21315 6341 21327 6344
rect 21269 6335 21327 6341
rect 22646 6332 22652 6344
rect 22704 6332 22710 6384
rect 25130 6332 25136 6384
rect 25188 6332 25194 6384
rect 18414 6264 18420 6316
rect 18472 6264 18478 6316
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6304 20315 6307
rect 21082 6304 21088 6316
rect 20303 6276 21088 6304
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 22094 6264 22100 6316
rect 22152 6264 22158 6316
rect 24026 6264 24032 6316
rect 24084 6264 24090 6316
rect 19245 6239 19303 6245
rect 19245 6205 19257 6239
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 19260 6168 19288 6199
rect 21910 6196 21916 6248
rect 21968 6236 21974 6248
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 21968 6208 22477 6236
rect 21968 6196 21974 6208
rect 22465 6205 22477 6208
rect 22511 6205 22523 6239
rect 22465 6199 22523 6205
rect 22830 6168 22836 6180
rect 19260 6140 22836 6168
rect 22830 6128 22836 6140
rect 22888 6128 22894 6180
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 20898 5856 20904 5908
rect 20956 5896 20962 5908
rect 24765 5899 24823 5905
rect 24765 5896 24777 5899
rect 20956 5868 24777 5896
rect 20956 5856 20962 5868
rect 24765 5865 24777 5868
rect 24811 5865 24823 5899
rect 24765 5859 24823 5865
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 20993 5763 21051 5769
rect 20993 5760 21005 5763
rect 20772 5732 21005 5760
rect 20772 5720 20778 5732
rect 20993 5729 21005 5732
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 21542 5720 21548 5772
rect 21600 5760 21606 5772
rect 22833 5763 22891 5769
rect 22833 5760 22845 5763
rect 21600 5732 22845 5760
rect 21600 5720 21606 5732
rect 22833 5729 22845 5732
rect 22879 5729 22891 5763
rect 22833 5723 22891 5729
rect 2590 5652 2596 5704
rect 2648 5692 2654 5704
rect 8754 5692 8760 5704
rect 2648 5664 8760 5692
rect 2648 5652 2654 5664
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 20530 5652 20536 5704
rect 20588 5652 20594 5704
rect 20622 5652 20628 5704
rect 20680 5692 20686 5704
rect 22373 5695 22431 5701
rect 22373 5692 22385 5695
rect 20680 5664 22385 5692
rect 20680 5652 20686 5664
rect 22373 5661 22385 5664
rect 22419 5661 22431 5695
rect 22373 5655 22431 5661
rect 22554 5652 22560 5704
rect 22612 5692 22618 5704
rect 24673 5695 24731 5701
rect 24673 5692 24685 5695
rect 22612 5664 24685 5692
rect 22612 5652 22618 5664
rect 24673 5661 24685 5664
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 15102 5624 15108 5636
rect 10100 5596 15108 5624
rect 10100 5584 10106 5596
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 11422 5556 11428 5568
rect 9364 5528 11428 5556
rect 9364 5516 9370 5528
rect 11422 5516 11428 5528
rect 11480 5516 11486 5568
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 18785 5287 18843 5293
rect 18785 5253 18797 5287
rect 18831 5284 18843 5287
rect 19610 5284 19616 5296
rect 18831 5256 19616 5284
rect 18831 5253 18843 5256
rect 18785 5247 18843 5253
rect 19610 5244 19616 5256
rect 19668 5244 19674 5296
rect 17770 5176 17776 5228
rect 17828 5176 17834 5228
rect 19518 5176 19524 5228
rect 19576 5176 19582 5228
rect 21818 5176 21824 5228
rect 21876 5216 21882 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21876 5188 22017 5216
rect 21876 5176 21882 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 24118 5176 24124 5228
rect 24176 5176 24182 5228
rect 19334 5108 19340 5160
rect 19392 5148 19398 5160
rect 19889 5151 19947 5157
rect 19889 5148 19901 5151
rect 19392 5120 19901 5148
rect 19392 5108 19398 5120
rect 19889 5117 19901 5120
rect 19935 5117 19947 5151
rect 19889 5111 19947 5117
rect 22462 5108 22468 5160
rect 22520 5108 22526 5160
rect 24762 5108 24768 5160
rect 24820 5108 24826 5160
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 17770 4700 17776 4752
rect 17828 4740 17834 4752
rect 17828 4712 23520 4740
rect 17828 4700 17834 4712
rect 19886 4632 19892 4684
rect 19944 4632 19950 4684
rect 21729 4675 21787 4681
rect 21729 4672 21741 4675
rect 19996 4644 21741 4672
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4604 17739 4607
rect 18506 4604 18512 4616
rect 17727 4576 18512 4604
rect 17727 4573 17739 4576
rect 17681 4567 17739 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 18598 4564 18604 4616
rect 18656 4604 18662 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 18656 4576 19441 4604
rect 18656 4564 18662 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 19702 4564 19708 4616
rect 19760 4604 19766 4616
rect 19996 4604 20024 4644
rect 21729 4641 21741 4644
rect 21775 4641 21787 4675
rect 21729 4635 21787 4641
rect 22738 4632 22744 4684
rect 22796 4672 22802 4684
rect 23492 4681 23520 4712
rect 24854 4700 24860 4752
rect 24912 4700 24918 4752
rect 23201 4675 23259 4681
rect 23201 4672 23213 4675
rect 22796 4644 23213 4672
rect 22796 4632 22802 4644
rect 23201 4641 23213 4644
rect 23247 4641 23259 4675
rect 23201 4635 23259 4641
rect 23477 4675 23535 4681
rect 23477 4641 23489 4675
rect 23523 4641 23535 4675
rect 23477 4635 23535 4641
rect 19760 4576 20024 4604
rect 19760 4564 19766 4576
rect 21266 4564 21272 4616
rect 21324 4564 21330 4616
rect 23290 4564 23296 4616
rect 23348 4604 23354 4616
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 23348 4576 24685 4604
rect 23348 4564 23354 4576
rect 24673 4573 24685 4576
rect 24719 4573 24731 4607
rect 24673 4567 24731 4573
rect 18693 4539 18751 4545
rect 18693 4505 18705 4539
rect 18739 4536 18751 4539
rect 20622 4536 20628 4548
rect 18739 4508 20628 4536
rect 18739 4505 18751 4508
rect 18693 4499 18751 4505
rect 20622 4496 20628 4508
rect 20680 4496 20686 4548
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 8202 4156 8208 4208
rect 8260 4196 8266 4208
rect 10318 4196 10324 4208
rect 8260 4168 10324 4196
rect 8260 4156 8266 4168
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 12618 4156 12624 4208
rect 12676 4196 12682 4208
rect 14182 4196 14188 4208
rect 12676 4168 14188 4196
rect 12676 4156 12682 4168
rect 14182 4156 14188 4168
rect 14240 4156 14246 4208
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 1504 4100 1777 4128
rect 1504 3924 1532 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 13446 4088 13452 4140
rect 13504 4128 13510 4140
rect 13541 4131 13599 4137
rect 13541 4128 13553 4131
rect 13504 4100 13553 4128
rect 13504 4088 13510 4100
rect 13541 4097 13553 4100
rect 13587 4097 13599 4131
rect 13541 4091 13599 4097
rect 16114 4088 16120 4140
rect 16172 4088 16178 4140
rect 16666 4088 16672 4140
rect 16724 4128 16730 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16724 4100 16865 4128
rect 16724 4088 16730 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 18690 4088 18696 4140
rect 18748 4088 18754 4140
rect 22094 4088 22100 4140
rect 22152 4088 22158 4140
rect 23842 4088 23848 4140
rect 23900 4088 23906 4140
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 6178 4060 6184 4072
rect 3200 4032 6184 4060
rect 3200 4020 3206 4032
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 11606 4060 11612 4072
rect 11379 4032 11612 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11606 4020 11612 4032
rect 11664 4060 11670 4072
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 11664 4032 11713 4060
rect 11664 4020 11670 4032
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11701 4023 11759 4029
rect 11977 4063 12035 4069
rect 11977 4029 11989 4063
rect 12023 4029 12035 4063
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 11977 4023 12035 4029
rect 13464 4032 14013 4060
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 2774 3992 2780 4004
rect 1627 3964 2780 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 9953 3995 10011 4001
rect 9953 3992 9965 3995
rect 9088 3964 9965 3992
rect 9088 3952 9094 3964
rect 9953 3961 9965 3964
rect 9999 3961 10011 3995
rect 9953 3955 10011 3961
rect 2041 3927 2099 3933
rect 2041 3924 2053 3927
rect 1504 3896 2053 3924
rect 2041 3893 2053 3896
rect 2087 3924 2099 3927
rect 2866 3924 2872 3936
rect 2087 3896 2872 3924
rect 2087 3893 2099 3896
rect 2041 3887 2099 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6144 3896 6377 3924
rect 6144 3884 6150 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 9456 3896 9505 3924
rect 9456 3884 9462 3896
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 9493 3887 9551 3893
rect 9766 3884 9772 3936
rect 9824 3884 9830 3936
rect 10502 3884 10508 3936
rect 10560 3924 10566 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10560 3896 11069 3924
rect 10560 3884 10566 3896
rect 11057 3893 11069 3896
rect 11103 3893 11115 3927
rect 11992 3924 12020 4023
rect 13464 4004 13492 4032
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16448 4032 17325 4060
rect 16448 4020 16454 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 17552 4032 19165 4060
rect 17552 4020 17558 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 20070 4020 20076 4072
rect 20128 4060 20134 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 20128 4032 22477 4060
rect 20128 4020 20134 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 13446 3952 13452 4004
rect 13504 3952 13510 4004
rect 16298 3952 16304 4004
rect 16356 3952 16362 4004
rect 21174 3952 21180 4004
rect 21232 3992 21238 4004
rect 24320 3992 24348 4023
rect 21232 3964 24348 3992
rect 21232 3952 21238 3964
rect 15930 3924 15936 3936
rect 11992 3896 15936 3924
rect 11057 3887 11115 3893
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 19610 3884 19616 3936
rect 19668 3924 19674 3936
rect 22370 3924 22376 3936
rect 19668 3896 22376 3924
rect 19668 3884 19674 3896
rect 22370 3884 22376 3896
rect 22428 3884 22434 3936
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 5258 3680 5264 3732
rect 5316 3680 5322 3732
rect 6730 3680 6736 3732
rect 6788 3680 6794 3732
rect 8202 3680 8208 3732
rect 8260 3680 8266 3732
rect 9309 3723 9367 3729
rect 9309 3689 9321 3723
rect 9355 3720 9367 3723
rect 9490 3720 9496 3732
rect 9355 3692 9496 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 10042 3680 10048 3732
rect 10100 3680 10106 3732
rect 22830 3680 22836 3732
rect 22888 3720 22894 3732
rect 24946 3720 24952 3732
rect 22888 3692 24952 3720
rect 22888 3680 22894 3692
rect 24946 3680 24952 3692
rect 25004 3680 25010 3732
rect 1765 3655 1823 3661
rect 1765 3621 1777 3655
rect 1811 3652 1823 3655
rect 5534 3652 5540 3664
rect 1811 3624 5540 3652
rect 1811 3621 1823 3624
rect 1765 3615 1823 3621
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 5905 3655 5963 3661
rect 5905 3621 5917 3655
rect 5951 3652 5963 3655
rect 16114 3652 16120 3664
rect 5951 3624 16120 3652
rect 5951 3621 5963 3624
rect 5905 3615 5963 3621
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 16574 3612 16580 3664
rect 16632 3652 16638 3664
rect 16632 3624 17724 3652
rect 16632 3612 16638 3624
rect 7561 3587 7619 3593
rect 7561 3553 7573 3587
rect 7607 3584 7619 3587
rect 8294 3584 8300 3596
rect 7607 3556 8300 3584
rect 7607 3553 7619 3556
rect 7561 3547 7619 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 11238 3544 11244 3596
rect 11296 3544 11302 3596
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 12805 3587 12863 3593
rect 12805 3584 12817 3587
rect 12768 3556 12817 3584
rect 12768 3544 12774 3556
rect 12805 3553 12817 3556
rect 12851 3553 12863 3587
rect 12805 3547 12863 3553
rect 14918 3544 14924 3596
rect 14976 3584 14982 3596
rect 15473 3587 15531 3593
rect 15473 3584 15485 3587
rect 14976 3556 15485 3584
rect 14976 3544 14982 3556
rect 15473 3553 15485 3556
rect 15519 3553 15531 3587
rect 15473 3547 15531 3553
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 16080 3556 17325 3584
rect 16080 3544 16086 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 1949 3519 2007 3525
rect 1949 3516 1961 3519
rect 1728 3488 1961 3516
rect 1728 3476 1734 3488
rect 1949 3485 1961 3488
rect 1995 3516 2007 3519
rect 2409 3519 2467 3525
rect 2409 3516 2421 3519
rect 1995 3488 2421 3516
rect 1995 3485 2007 3488
rect 1949 3479 2007 3485
rect 2409 3485 2421 3488
rect 2455 3485 2467 3519
rect 5077 3519 5135 3525
rect 5077 3516 5089 3519
rect 2409 3479 2467 3485
rect 5000 3488 5089 3516
rect 3145 3451 3203 3457
rect 3145 3417 3157 3451
rect 3191 3448 3203 3451
rect 3326 3448 3332 3460
rect 3191 3420 3332 3448
rect 3191 3417 3203 3420
rect 3145 3411 3203 3417
rect 3326 3408 3332 3420
rect 3384 3408 3390 3460
rect 5000 3392 5028 3488
rect 5077 3485 5089 3488
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 6086 3476 6092 3528
rect 6144 3476 6150 3528
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6512 3488 6561 3516
rect 6512 3476 6518 3488
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 6549 3479 6607 3485
rect 7852 3488 8033 3516
rect 7852 3392 7880 3488
rect 8021 3485 8033 3488
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3516 9183 3519
rect 9398 3516 9404 3528
rect 9171 3488 9404 3516
rect 9171 3485 9183 3488
rect 9125 3479 9183 3485
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9824 3488 9873 3516
rect 9824 3476 9830 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 10870 3516 10876 3528
rect 10551 3488 10876 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 10870 3476 10876 3488
rect 10928 3516 10934 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 10928 3488 10977 3516
rect 10928 3476 10934 3488
rect 10965 3485 10977 3488
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 12434 3476 12440 3528
rect 12492 3476 12498 3528
rect 15102 3476 15108 3528
rect 15160 3476 15166 3528
rect 16206 3476 16212 3528
rect 16264 3516 16270 3528
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16264 3488 16865 3516
rect 16264 3476 16270 3488
rect 16853 3485 16865 3488
rect 16899 3485 16911 3519
rect 17696 3516 17724 3624
rect 17862 3544 17868 3596
rect 17920 3584 17926 3596
rect 19889 3587 19947 3593
rect 19889 3584 19901 3587
rect 17920 3556 19901 3584
rect 17920 3544 17926 3556
rect 19889 3553 19901 3556
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 17696 3488 19441 3516
rect 16853 3479 16911 3485
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 20990 3476 20996 3528
rect 21048 3516 21054 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 21048 3488 21281 3516
rect 21048 3476 21054 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 18966 3408 18972 3460
rect 19024 3448 19030 3460
rect 21744 3448 21772 3547
rect 19024 3420 21772 3448
rect 19024 3408 19030 3420
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 2096 3352 2237 3380
rect 2096 3340 2102 3352
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 2225 3343 2283 3349
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 2869 3383 2927 3389
rect 2869 3380 2881 3383
rect 2832 3352 2881 3380
rect 2832 3340 2838 3352
rect 2869 3349 2881 3352
rect 2915 3349 2927 3383
rect 2869 3343 2927 3349
rect 3237 3383 3295 3389
rect 3237 3349 3249 3383
rect 3283 3380 3295 3383
rect 3418 3380 3424 3392
rect 3283 3352 3424 3380
rect 3283 3349 3295 3352
rect 3237 3343 3295 3349
rect 3418 3340 3424 3352
rect 3476 3340 3482 3392
rect 3605 3383 3663 3389
rect 3605 3349 3617 3383
rect 3651 3380 3663 3383
rect 3878 3380 3884 3392
rect 3651 3352 3884 3380
rect 3651 3349 3663 3352
rect 3605 3343 3663 3349
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 4801 3383 4859 3389
rect 4801 3349 4813 3383
rect 4847 3380 4859 3383
rect 4982 3380 4988 3392
rect 4847 3352 4988 3380
rect 4847 3349 4859 3352
rect 4801 3343 4859 3349
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7193 3383 7251 3389
rect 7193 3380 7205 3383
rect 6880 3352 7205 3380
rect 6880 3340 6886 3352
rect 7193 3349 7205 3352
rect 7239 3349 7251 3383
rect 7193 3343 7251 3349
rect 7745 3383 7803 3389
rect 7745 3349 7757 3383
rect 7791 3380 7803 3383
rect 7834 3380 7840 3392
rect 7791 3352 7840 3380
rect 7791 3349 7803 3352
rect 7745 3343 7803 3349
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 8662 3340 8668 3392
rect 8720 3340 8726 3392
rect 10689 3383 10747 3389
rect 10689 3349 10701 3383
rect 10735 3380 10747 3383
rect 11238 3380 11244 3392
rect 10735 3352 11244 3380
rect 10735 3349 10747 3352
rect 10689 3343 10747 3349
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 22002 3340 22008 3392
rect 22060 3380 22066 3392
rect 22830 3380 22836 3392
rect 22060 3352 22836 3380
rect 22060 3340 22066 3352
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 23566 3340 23572 3392
rect 23624 3380 23630 3392
rect 24118 3380 24124 3392
rect 23624 3352 24124 3380
rect 23624 3340 23630 3352
rect 24118 3340 24124 3352
rect 24176 3380 24182 3392
rect 25409 3383 25467 3389
rect 25409 3380 25421 3383
rect 24176 3352 25421 3380
rect 24176 3340 24182 3352
rect 25409 3349 25421 3352
rect 25455 3349 25467 3383
rect 25409 3343 25467 3349
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 2682 3136 2688 3188
rect 2740 3136 2746 3188
rect 5166 3136 5172 3188
rect 5224 3136 5230 3188
rect 5902 3136 5908 3188
rect 5960 3136 5966 3188
rect 7006 3136 7012 3188
rect 7064 3136 7070 3188
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7248 3148 7757 3176
rect 7248 3136 7254 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 8478 3136 8484 3188
rect 8536 3136 8542 3188
rect 11882 3136 11888 3188
rect 11940 3136 11946 3188
rect 24670 3136 24676 3188
rect 24728 3176 24734 3188
rect 24857 3179 24915 3185
rect 24857 3176 24869 3179
rect 24728 3148 24869 3176
rect 24728 3136 24734 3148
rect 24857 3145 24869 3148
rect 24903 3145 24915 3179
rect 24857 3139 24915 3145
rect 14826 3108 14832 3120
rect 10612 3080 14832 3108
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2038 3040 2044 3052
rect 1903 3012 2044 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2038 3000 2044 3012
rect 2096 3000 2102 3052
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2774 3040 2780 3052
rect 2547 3012 2780 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 3510 3000 3516 3052
rect 3568 3000 3574 3052
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3040 4767 3043
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4755 3012 4997 3040
rect 4755 3009 4767 3012
rect 4709 3003 4767 3009
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 5350 3040 5356 3052
rect 5031 3012 5356 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5718 3000 5724 3052
rect 5776 3000 5782 3052
rect 6822 3000 6828 3052
rect 6880 3000 6886 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 8202 3040 8208 3052
rect 7607 3012 8208 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 8662 3040 8668 3052
rect 8343 3012 8668 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 9306 3000 9312 3052
rect 9364 3000 9370 3052
rect 10612 3049 10640 3080
rect 14826 3068 14832 3080
rect 14884 3068 14890 3120
rect 18598 3068 18604 3120
rect 18656 3108 18662 3120
rect 19886 3108 19892 3120
rect 18656 3080 19892 3108
rect 18656 3068 18662 3080
rect 19886 3068 19892 3080
rect 19944 3068 19950 3120
rect 23566 3068 23572 3120
rect 23624 3068 23630 3120
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11296 3012 11713 3040
rect 11296 3000 11302 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 12618 3000 12624 3052
rect 12676 3000 12682 3052
rect 14274 3000 14280 3052
rect 14332 3000 14338 3052
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16816 3012 16865 3040
rect 16816 3000 16822 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 16942 3000 16948 3052
rect 17000 3040 17006 3052
rect 18693 3043 18751 3049
rect 18693 3040 18705 3043
rect 17000 3012 18705 3040
rect 17000 3000 17006 3012
rect 18693 3009 18705 3012
rect 18739 3009 18751 3043
rect 18693 3003 18751 3009
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2972 3295 2975
rect 3326 2972 3332 2984
rect 3283 2944 3332 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 9030 2932 9036 2984
rect 9088 2932 9094 2984
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2972 10379 2975
rect 10502 2972 10508 2984
rect 10367 2944 10508 2972
rect 10367 2941 10379 2944
rect 10321 2935 10379 2941
rect 10502 2932 10508 2944
rect 10560 2932 10566 2984
rect 13354 2932 13360 2984
rect 13412 2932 13418 2984
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14240 2944 14749 2972
rect 14240 2932 14246 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15712 2944 17325 2972
rect 15712 2932 15718 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 2041 2907 2099 2913
rect 2041 2873 2053 2907
rect 2087 2904 2099 2907
rect 4890 2904 4896 2916
rect 2087 2876 4896 2904
rect 2087 2873 2099 2876
rect 2041 2867 2099 2873
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
rect 17126 2864 17132 2916
rect 17184 2904 17190 2916
rect 19168 2904 19196 2935
rect 17184 2876 19196 2904
rect 17184 2864 17190 2876
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 23382 2904 23388 2916
rect 20680 2876 23388 2904
rect 20680 2864 20686 2876
rect 23382 2864 23388 2876
rect 23440 2864 23446 2916
rect 1486 2796 1492 2848
rect 1544 2796 1550 2848
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 4341 2839 4399 2845
rect 4341 2836 4353 2839
rect 4304 2808 4353 2836
rect 4304 2796 4310 2808
rect 4341 2805 4353 2808
rect 4387 2805 4399 2839
rect 4341 2799 4399 2805
rect 6454 2796 6460 2848
rect 6512 2796 6518 2848
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 19886 2836 19892 2848
rect 16816 2808 19892 2836
rect 16816 2796 16822 2808
rect 19886 2796 19892 2808
rect 19944 2796 19950 2848
rect 20806 2796 20812 2848
rect 20864 2836 20870 2848
rect 22462 2836 22468 2848
rect 20864 2808 22468 2836
rect 20864 2796 20870 2808
rect 22462 2796 22468 2808
rect 22520 2796 22526 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 1854 2592 1860 2644
rect 1912 2592 1918 2644
rect 2590 2592 2596 2644
rect 2648 2592 2654 2644
rect 4154 2592 4160 2644
rect 4212 2592 4218 2644
rect 7098 2592 7104 2644
rect 7156 2592 7162 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 11790 2632 11796 2644
rect 9815 2604 11796 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 11790 2592 11796 2604
rect 11848 2592 11854 2644
rect 3329 2567 3387 2573
rect 3329 2533 3341 2567
rect 3375 2564 3387 2567
rect 4798 2564 4804 2576
rect 3375 2536 4804 2564
rect 3375 2533 3387 2536
rect 3329 2527 3387 2533
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 8938 2564 8944 2576
rect 6886 2536 8944 2564
rect 4985 2499 5043 2505
rect 4985 2465 4997 2499
rect 5031 2496 5043 2499
rect 6886 2496 6914 2536
rect 8938 2524 8944 2536
rect 8996 2524 9002 2576
rect 12802 2564 12808 2576
rect 10612 2536 12808 2564
rect 5031 2468 6914 2496
rect 5031 2465 5043 2468
rect 4985 2459 5043 2465
rect 7742 2456 7748 2508
rect 7800 2496 7806 2508
rect 10612 2505 10640 2536
rect 12802 2524 12808 2536
rect 12860 2524 12866 2576
rect 7929 2499 7987 2505
rect 7929 2496 7941 2499
rect 7800 2468 7941 2496
rect 7800 2456 7806 2468
rect 7929 2465 7941 2468
rect 7975 2465 7987 2499
rect 7929 2459 7987 2465
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2465 10655 2499
rect 11974 2496 11980 2508
rect 10597 2459 10655 2465
rect 11900 2468 11980 2496
rect 1486 2388 1492 2440
rect 1544 2428 1550 2440
rect 1673 2431 1731 2437
rect 1673 2428 1685 2431
rect 1544 2400 1685 2428
rect 1544 2388 1550 2400
rect 1673 2397 1685 2400
rect 1719 2428 1731 2431
rect 2314 2428 2320 2440
rect 1719 2400 2320 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2428 3203 2431
rect 3878 2428 3884 2440
rect 3191 2400 3884 2428
rect 3191 2397 3203 2400
rect 3145 2391 3203 2397
rect 2424 2360 2452 2391
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4246 2428 4252 2440
rect 4019 2400 4252 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 4614 2388 4620 2440
rect 4672 2428 4678 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4672 2400 4721 2428
rect 4672 2388 4678 2400
rect 4709 2397 4721 2400
rect 4755 2428 4767 2431
rect 5813 2431 5871 2437
rect 5813 2428 5825 2431
rect 4755 2400 5825 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5813 2397 5825 2400
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6503 2400 6929 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 6917 2397 6929 2400
rect 6963 2428 6975 2431
rect 7190 2428 7196 2440
rect 6963 2400 7196 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7616 2400 7665 2428
rect 7616 2388 7622 2400
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9585 2431 9643 2437
rect 9585 2428 9597 2431
rect 9171 2400 9597 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9585 2397 9597 2400
rect 9631 2428 9643 2431
rect 10134 2428 10140 2440
rect 9631 2400 10140 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 11900 2437 11928 2468
rect 11974 2456 11980 2468
rect 12032 2496 12038 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 12032 2468 14105 2496
rect 12032 2456 12038 2468
rect 14093 2465 14105 2468
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 14608 2468 15209 2496
rect 14608 2456 14614 2468
rect 15197 2465 15209 2468
rect 15243 2465 15255 2499
rect 15197 2459 15255 2465
rect 15286 2456 15292 2508
rect 15344 2496 15350 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 15344 2468 17325 2496
rect 15344 2456 15350 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 17678 2456 17684 2508
rect 17736 2496 17742 2508
rect 17736 2468 19564 2496
rect 17736 2456 17742 2468
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 3510 2360 3516 2372
rect 2424 2332 3516 2360
rect 3510 2320 3516 2332
rect 3568 2320 3574 2372
rect 5718 2320 5724 2372
rect 5776 2360 5782 2372
rect 6089 2363 6147 2369
rect 6089 2360 6101 2363
rect 5776 2332 6101 2360
rect 5776 2320 5782 2332
rect 6089 2329 6101 2332
rect 6135 2329 6147 2363
rect 6089 2323 6147 2329
rect 6641 2363 6699 2369
rect 6641 2329 6653 2363
rect 6687 2360 6699 2363
rect 7576 2360 7604 2388
rect 6687 2332 7604 2360
rect 9309 2363 9367 2369
rect 6687 2329 6699 2332
rect 6641 2323 6699 2329
rect 9309 2329 9321 2363
rect 9355 2360 9367 2363
rect 10336 2360 10364 2391
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 14642 2388 14648 2440
rect 14700 2388 14706 2440
rect 16850 2388 16856 2440
rect 16908 2388 16914 2440
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 19536 2428 19564 2468
rect 19886 2456 19892 2508
rect 19944 2456 19950 2508
rect 22465 2499 22523 2505
rect 22465 2465 22477 2499
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 19536 2400 22017 2428
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 12342 2360 12348 2372
rect 9355 2332 12348 2360
rect 9355 2329 9367 2332
rect 9309 2323 9367 2329
rect 12342 2320 12348 2332
rect 12400 2320 12406 2372
rect 13541 2363 13599 2369
rect 13541 2329 13553 2363
rect 13587 2360 13599 2363
rect 13814 2360 13820 2372
rect 13587 2332 13820 2360
rect 13587 2329 13599 2332
rect 13541 2323 13599 2329
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 18322 2320 18328 2372
rect 18380 2360 18386 2372
rect 22480 2360 22508 2459
rect 25314 2388 25320 2440
rect 25372 2388 25378 2440
rect 18380 2332 22508 2360
rect 18380 2320 18386 2332
rect 11701 2295 11759 2301
rect 11701 2261 11713 2295
rect 11747 2292 11759 2295
rect 15378 2292 15384 2304
rect 11747 2264 15384 2292
rect 11747 2261 11759 2264
rect 11701 2255 11759 2261
rect 15378 2252 15384 2264
rect 15436 2252 15442 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 3142 2048 3148 2100
rect 3200 2088 3206 2100
rect 9030 2088 9036 2100
rect 3200 2060 9036 2088
rect 3200 2048 3206 2060
rect 9030 2048 9036 2060
rect 9088 2048 9094 2100
rect 8294 1980 8300 2032
rect 8352 2020 8358 2032
rect 15930 2020 15936 2032
rect 8352 1992 15936 2020
rect 8352 1980 8358 1992
rect 15930 1980 15936 1992
rect 15988 1980 15994 2032
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 9956 54272 10008 54324
rect 14740 54272 14792 54324
rect 16212 54272 16264 54324
rect 7840 54204 7892 54256
rect 11428 54204 11480 54256
rect 4528 54136 4580 54188
rect 4620 54179 4672 54188
rect 4620 54145 4629 54179
rect 4629 54145 4663 54179
rect 4663 54145 4672 54179
rect 4620 54136 4672 54145
rect 5908 54068 5960 54120
rect 9956 54179 10008 54188
rect 9956 54145 9965 54179
rect 9965 54145 9999 54179
rect 9999 54145 10008 54179
rect 9956 54136 10008 54145
rect 12900 54204 12952 54256
rect 12348 54179 12400 54188
rect 12348 54145 12357 54179
rect 12357 54145 12391 54179
rect 12391 54145 12400 54179
rect 12348 54136 12400 54145
rect 15200 54136 15252 54188
rect 24492 54315 24544 54324
rect 24492 54281 24501 54315
rect 24501 54281 24535 54315
rect 24535 54281 24544 54315
rect 24492 54272 24544 54281
rect 17684 54204 17736 54256
rect 18880 54204 18932 54256
rect 16948 54136 17000 54188
rect 11244 54068 11296 54120
rect 12532 54068 12584 54120
rect 18420 54068 18472 54120
rect 19524 54136 19576 54188
rect 20720 54136 20772 54188
rect 21364 54136 21416 54188
rect 22468 54136 22520 54188
rect 24952 54179 25004 54188
rect 24952 54145 24961 54179
rect 24961 54145 24995 54179
rect 24995 54145 25004 54179
rect 24952 54136 25004 54145
rect 19708 54068 19760 54120
rect 15384 54000 15436 54052
rect 25136 54043 25188 54052
rect 25136 54009 25145 54043
rect 25145 54009 25179 54043
rect 25179 54009 25188 54043
rect 25136 54000 25188 54009
rect 11704 53975 11756 53984
rect 11704 53941 11713 53975
rect 11713 53941 11747 53975
rect 11747 53941 11756 53975
rect 11704 53932 11756 53941
rect 14096 53932 14148 53984
rect 15292 53932 15344 53984
rect 17040 53975 17092 53984
rect 17040 53941 17049 53975
rect 17049 53941 17083 53975
rect 17083 53941 17092 53975
rect 17040 53932 17092 53941
rect 18512 53975 18564 53984
rect 18512 53941 18521 53975
rect 18521 53941 18555 53975
rect 18555 53941 18564 53975
rect 18512 53932 18564 53941
rect 19340 53932 19392 53984
rect 20904 53932 20956 53984
rect 21548 53932 21600 53984
rect 22192 53975 22244 53984
rect 22192 53941 22201 53975
rect 22201 53941 22235 53975
rect 22235 53941 22244 53975
rect 22192 53932 22244 53941
rect 22744 53932 22796 53984
rect 24124 53932 24176 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 16580 53728 16632 53780
rect 18880 53771 18932 53780
rect 18880 53737 18889 53771
rect 18889 53737 18923 53771
rect 18923 53737 18932 53771
rect 18880 53728 18932 53737
rect 5540 53660 5592 53712
rect 21640 53660 21692 53712
rect 22376 53660 22428 53712
rect 7380 53592 7432 53644
rect 8852 53592 8904 53644
rect 11060 53635 11112 53644
rect 11060 53601 11069 53635
rect 11069 53601 11103 53635
rect 11103 53601 11112 53635
rect 11060 53592 11112 53601
rect 12164 53592 12216 53644
rect 6828 53524 6880 53576
rect 9128 53524 9180 53576
rect 10416 53567 10468 53576
rect 10416 53533 10425 53567
rect 10425 53533 10459 53567
rect 10459 53533 10468 53567
rect 10416 53524 10468 53533
rect 12624 53524 12676 53576
rect 14004 53524 14056 53576
rect 15476 53524 15528 53576
rect 16580 53524 16632 53576
rect 17316 53524 17368 53576
rect 18328 53524 18380 53576
rect 19156 53524 19208 53576
rect 19892 53524 19944 53576
rect 20996 53524 21048 53576
rect 21732 53524 21784 53576
rect 22100 53524 22152 53576
rect 22836 53524 22888 53576
rect 23388 53524 23440 53576
rect 24768 53524 24820 53576
rect 7380 53456 7432 53508
rect 16396 53456 16448 53508
rect 20444 53499 20496 53508
rect 20444 53465 20453 53499
rect 20453 53465 20487 53499
rect 20487 53465 20496 53499
rect 20444 53456 20496 53465
rect 24216 53456 24268 53508
rect 14464 53431 14516 53440
rect 14464 53397 14473 53431
rect 14473 53397 14507 53431
rect 14507 53397 14516 53431
rect 14464 53388 14516 53397
rect 16856 53431 16908 53440
rect 16856 53397 16865 53431
rect 16865 53397 16899 53431
rect 16899 53397 16908 53431
rect 16856 53388 16908 53397
rect 17408 53431 17460 53440
rect 17408 53397 17417 53431
rect 17417 53397 17451 53431
rect 17451 53397 17460 53431
rect 17408 53388 17460 53397
rect 18328 53431 18380 53440
rect 18328 53397 18337 53431
rect 18337 53397 18371 53431
rect 18371 53397 18380 53431
rect 18328 53388 18380 53397
rect 19616 53431 19668 53440
rect 19616 53397 19625 53431
rect 19625 53397 19659 53431
rect 19659 53397 19668 53431
rect 19616 53388 19668 53397
rect 21364 53388 21416 53440
rect 22468 53431 22520 53440
rect 22468 53397 22477 53431
rect 22477 53397 22511 53431
rect 22511 53397 22520 53431
rect 22468 53388 22520 53397
rect 25872 53388 25924 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 2780 53184 2832 53236
rect 17316 53227 17368 53236
rect 17316 53193 17325 53227
rect 17325 53193 17359 53227
rect 17359 53193 17368 53227
rect 17316 53184 17368 53193
rect 19156 53184 19208 53236
rect 19708 53227 19760 53236
rect 19708 53193 19717 53227
rect 19717 53193 19751 53227
rect 19751 53193 19760 53227
rect 19708 53184 19760 53193
rect 20996 53227 21048 53236
rect 20996 53193 21005 53227
rect 21005 53193 21039 53227
rect 21039 53193 21048 53227
rect 20996 53184 21048 53193
rect 21732 53184 21784 53236
rect 22100 53184 22152 53236
rect 22560 53227 22612 53236
rect 22560 53193 22569 53227
rect 22569 53193 22603 53227
rect 22603 53193 22612 53227
rect 22560 53184 22612 53193
rect 23296 53184 23348 53236
rect 4436 53116 4488 53168
rect 6276 53116 6328 53168
rect 9220 53116 9272 53168
rect 13636 53116 13688 53168
rect 20720 53116 20772 53168
rect 6368 53048 6420 53100
rect 5632 52980 5684 53032
rect 9680 53048 9732 53100
rect 11888 53091 11940 53100
rect 11888 53057 11897 53091
rect 11897 53057 11931 53091
rect 11931 53057 11940 53091
rect 11888 53048 11940 53057
rect 14372 53048 14424 53100
rect 15844 53048 15896 53100
rect 18788 53048 18840 53100
rect 20260 53048 20312 53100
rect 23572 53048 23624 53100
rect 25044 53091 25096 53100
rect 25044 53057 25053 53091
rect 25053 53057 25087 53091
rect 25087 53057 25096 53091
rect 25044 53048 25096 53057
rect 10232 52980 10284 53032
rect 10324 53023 10376 53032
rect 10324 52989 10333 53023
rect 10333 52989 10367 53023
rect 10367 52989 10376 53023
rect 10324 52980 10376 52989
rect 11796 52980 11848 53032
rect 3976 52912 4028 52964
rect 14004 52955 14056 52964
rect 14004 52921 14013 52955
rect 14013 52921 14047 52955
rect 14047 52921 14056 52955
rect 14004 52912 14056 52921
rect 1860 52844 1912 52896
rect 3516 52844 3568 52896
rect 14464 52887 14516 52896
rect 14464 52853 14473 52887
rect 14473 52853 14507 52887
rect 14507 52853 14516 52887
rect 14464 52844 14516 52853
rect 15936 52887 15988 52896
rect 15936 52853 15945 52887
rect 15945 52853 15979 52887
rect 15979 52853 15988 52887
rect 15936 52844 15988 52853
rect 18604 52844 18656 52896
rect 20168 52844 20220 52896
rect 22192 52844 22244 52896
rect 23940 52887 23992 52896
rect 23940 52853 23949 52887
rect 23949 52853 23983 52887
rect 23983 52853 23992 52887
rect 23940 52844 23992 52853
rect 25228 52887 25280 52896
rect 25228 52853 25237 52887
rect 25237 52853 25271 52887
rect 25271 52853 25280 52887
rect 25228 52844 25280 52853
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 2228 52640 2280 52692
rect 3424 52640 3476 52692
rect 12624 52683 12676 52692
rect 12624 52649 12633 52683
rect 12633 52649 12667 52683
rect 12667 52649 12676 52683
rect 12624 52640 12676 52649
rect 13636 52640 13688 52692
rect 24768 52640 24820 52692
rect 1308 52572 1360 52624
rect 3792 52572 3844 52624
rect 3700 52504 3752 52556
rect 25596 52572 25648 52624
rect 5172 52436 5224 52488
rect 5724 52436 5776 52488
rect 6644 52436 6696 52488
rect 7288 52479 7340 52488
rect 7288 52445 7297 52479
rect 7297 52445 7331 52479
rect 7331 52445 7340 52479
rect 7288 52436 7340 52445
rect 7748 52547 7800 52556
rect 7748 52513 7757 52547
rect 7757 52513 7791 52547
rect 7791 52513 7800 52547
rect 7748 52504 7800 52513
rect 10692 52504 10744 52556
rect 8944 52436 8996 52488
rect 10784 52479 10836 52488
rect 10784 52445 10793 52479
rect 10793 52445 10827 52479
rect 10827 52445 10836 52479
rect 10784 52436 10836 52445
rect 12808 52479 12860 52488
rect 12808 52445 12817 52479
rect 12817 52445 12851 52479
rect 12851 52445 12860 52479
rect 12808 52436 12860 52445
rect 13544 52436 13596 52488
rect 24768 52479 24820 52488
rect 24768 52445 24777 52479
rect 24777 52445 24811 52479
rect 24811 52445 24820 52479
rect 24768 52436 24820 52445
rect 13360 52368 13412 52420
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 5632 52096 5684 52148
rect 11888 52096 11940 52148
rect 12348 52139 12400 52148
rect 12348 52105 12357 52139
rect 12357 52105 12391 52139
rect 12391 52105 12400 52139
rect 12348 52096 12400 52105
rect 13360 52096 13412 52148
rect 24952 52096 25004 52148
rect 4896 52028 4948 52080
rect 9036 52028 9088 52080
rect 4712 52003 4764 52012
rect 4712 51969 4721 52003
rect 4721 51969 4755 52003
rect 4755 51969 4764 52003
rect 4712 51960 4764 51969
rect 10140 52028 10192 52080
rect 9772 52003 9824 52012
rect 9772 51969 9781 52003
rect 9781 51969 9815 52003
rect 9815 51969 9824 52003
rect 9772 51960 9824 51969
rect 10876 51960 10928 52012
rect 11980 51960 12032 52012
rect 3332 51935 3384 51944
rect 3332 51901 3341 51935
rect 3341 51901 3375 51935
rect 3375 51901 3384 51935
rect 3332 51892 3384 51901
rect 4804 51892 4856 51944
rect 8484 51935 8536 51944
rect 8484 51901 8493 51935
rect 8493 51901 8527 51935
rect 8527 51901 8536 51935
rect 8484 51892 8536 51901
rect 9864 51892 9916 51944
rect 25504 51799 25556 51808
rect 25504 51765 25513 51799
rect 25513 51765 25547 51799
rect 25547 51765 25556 51799
rect 25504 51756 25556 51765
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 3792 51595 3844 51604
rect 3792 51561 3801 51595
rect 3801 51561 3835 51595
rect 3835 51561 3844 51595
rect 3792 51552 3844 51561
rect 9956 51552 10008 51604
rect 2872 51459 2924 51468
rect 2872 51425 2881 51459
rect 2881 51425 2915 51459
rect 2915 51425 2924 51459
rect 2872 51416 2924 51425
rect 5540 51416 5592 51468
rect 7012 51416 7064 51468
rect 6736 51348 6788 51400
rect 7104 51391 7156 51400
rect 7104 51357 7113 51391
rect 7113 51357 7147 51391
rect 7147 51357 7156 51391
rect 7104 51348 7156 51357
rect 9220 51348 9272 51400
rect 25504 51348 25556 51400
rect 5540 51280 5592 51332
rect 25688 51212 25740 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 5540 51008 5592 51060
rect 4344 50940 4396 50992
rect 4528 50940 4580 50992
rect 4160 50915 4212 50924
rect 4160 50881 4169 50915
rect 4169 50881 4203 50915
rect 4203 50881 4212 50915
rect 4160 50872 4212 50881
rect 7656 50872 7708 50924
rect 10784 50940 10836 50992
rect 7840 50872 7892 50924
rect 25044 50915 25096 50924
rect 25044 50881 25053 50915
rect 25053 50881 25087 50915
rect 25087 50881 25096 50915
rect 25044 50872 25096 50881
rect 2780 50847 2832 50856
rect 2780 50813 2789 50847
rect 2789 50813 2823 50847
rect 2823 50813 2832 50847
rect 2780 50804 2832 50813
rect 4252 50804 4304 50856
rect 7472 50847 7524 50856
rect 7472 50813 7481 50847
rect 7481 50813 7515 50847
rect 7515 50813 7524 50847
rect 7472 50804 7524 50813
rect 15844 50804 15896 50856
rect 16856 50804 16908 50856
rect 25412 50668 25464 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 6828 50507 6880 50516
rect 6828 50473 6837 50507
rect 6837 50473 6871 50507
rect 6871 50473 6880 50507
rect 6828 50464 6880 50473
rect 9128 50464 9180 50516
rect 1308 50328 1360 50380
rect 3424 50260 3476 50312
rect 5816 50260 5868 50312
rect 8392 50260 8444 50312
rect 7564 50192 7616 50244
rect 5080 50124 5132 50176
rect 25320 50124 25372 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 3516 49852 3568 49904
rect 3332 49784 3384 49836
rect 10232 49920 10284 49972
rect 20996 49920 21048 49972
rect 7748 49784 7800 49836
rect 9680 49852 9732 49904
rect 9496 49784 9548 49836
rect 25320 49827 25372 49836
rect 25320 49793 25329 49827
rect 25329 49793 25363 49827
rect 25363 49793 25372 49827
rect 25320 49784 25372 49793
rect 8852 49716 8904 49768
rect 11704 49716 11756 49768
rect 12716 49716 12768 49768
rect 3976 49580 4028 49632
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 11980 49376 12032 49428
rect 1492 49240 1544 49292
rect 10600 49172 10652 49224
rect 10692 49172 10744 49224
rect 25320 49215 25372 49224
rect 25320 49181 25329 49215
rect 25329 49181 25363 49215
rect 25363 49181 25372 49215
rect 25320 49172 25372 49181
rect 25136 49079 25188 49088
rect 25136 49045 25145 49079
rect 25145 49045 25179 49079
rect 25179 49045 25188 49079
rect 25136 49036 25188 49045
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 12808 48832 12860 48884
rect 12532 48696 12584 48748
rect 25780 48492 25832 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 17316 48220 17368 48272
rect 17684 48220 17736 48272
rect 18512 48220 18564 48272
rect 25320 48127 25372 48136
rect 25320 48093 25329 48127
rect 25329 48093 25363 48127
rect 25363 48093 25372 48127
rect 25320 48084 25372 48093
rect 1308 48016 1360 48068
rect 8300 48016 8352 48068
rect 24860 47948 24912 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 9036 47744 9088 47796
rect 15936 47744 15988 47796
rect 17316 47787 17368 47796
rect 17316 47753 17325 47787
rect 17325 47753 17359 47787
rect 17359 47753 17368 47787
rect 17316 47744 17368 47753
rect 17408 47744 17460 47796
rect 18328 47676 18380 47728
rect 18788 47676 18840 47728
rect 11796 47608 11848 47660
rect 25780 47608 25832 47660
rect 16304 47472 16356 47524
rect 18696 47583 18748 47592
rect 18696 47549 18705 47583
rect 18705 47549 18739 47583
rect 18739 47549 18748 47583
rect 18696 47540 18748 47549
rect 23848 47540 23900 47592
rect 16580 47404 16632 47456
rect 17500 47404 17552 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 18696 47200 18748 47252
rect 19340 47243 19392 47252
rect 19340 47209 19349 47243
rect 19349 47209 19383 47243
rect 19383 47209 19392 47243
rect 19340 47200 19392 47209
rect 20444 47200 20496 47252
rect 18512 47132 18564 47184
rect 10232 47107 10284 47116
rect 10232 47073 10241 47107
rect 10241 47073 10275 47107
rect 10275 47073 10284 47107
rect 10232 47064 10284 47073
rect 16672 47064 16724 47116
rect 17224 47064 17276 47116
rect 18604 47107 18656 47116
rect 18604 47073 18613 47107
rect 18613 47073 18647 47107
rect 18647 47073 18656 47107
rect 18604 47064 18656 47073
rect 19340 47064 19392 47116
rect 25596 47132 25648 47184
rect 22468 47107 22520 47116
rect 22468 47073 22477 47107
rect 22477 47073 22511 47107
rect 22511 47073 22520 47107
rect 22468 47064 22520 47073
rect 22560 47107 22612 47116
rect 22560 47073 22569 47107
rect 22569 47073 22603 47107
rect 22603 47073 22612 47107
rect 22560 47064 22612 47073
rect 10784 46928 10836 46980
rect 12164 46860 12216 46912
rect 16396 46928 16448 46980
rect 18604 46928 18656 46980
rect 24768 46928 24820 46980
rect 13912 46860 13964 46912
rect 17592 46860 17644 46912
rect 22008 46903 22060 46912
rect 22008 46869 22017 46903
rect 22017 46869 22051 46903
rect 22051 46869 22060 46903
rect 22008 46860 22060 46869
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 7472 46656 7524 46708
rect 10876 46699 10928 46708
rect 10876 46665 10885 46699
rect 10885 46665 10919 46699
rect 10919 46665 10928 46699
rect 10876 46656 10928 46665
rect 14188 46656 14240 46708
rect 18696 46656 18748 46708
rect 18972 46656 19024 46708
rect 21916 46656 21968 46708
rect 22100 46656 22152 46708
rect 23940 46656 23992 46708
rect 13912 46588 13964 46640
rect 17592 46588 17644 46640
rect 9312 46520 9364 46572
rect 11060 46563 11112 46572
rect 11060 46529 11069 46563
rect 11069 46529 11103 46563
rect 11103 46529 11112 46563
rect 11060 46520 11112 46529
rect 11888 46316 11940 46368
rect 13360 46316 13412 46368
rect 16672 46452 16724 46504
rect 16856 46495 16908 46504
rect 16856 46461 16865 46495
rect 16865 46461 16899 46495
rect 16899 46461 16908 46495
rect 16856 46452 16908 46461
rect 18788 46452 18840 46504
rect 13728 46316 13780 46368
rect 16304 46359 16356 46368
rect 16304 46325 16313 46359
rect 16313 46325 16347 46359
rect 16347 46325 16356 46359
rect 16304 46316 16356 46325
rect 19340 46495 19392 46504
rect 19340 46461 19349 46495
rect 19349 46461 19383 46495
rect 19383 46461 19392 46495
rect 19340 46452 19392 46461
rect 20536 46452 20588 46504
rect 22652 46384 22704 46436
rect 24492 46495 24544 46504
rect 24492 46461 24501 46495
rect 24501 46461 24535 46495
rect 24535 46461 24544 46495
rect 24492 46452 24544 46461
rect 24676 46452 24728 46504
rect 19524 46316 19576 46368
rect 23296 46316 23348 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 5724 46112 5776 46164
rect 9220 46112 9272 46164
rect 10692 46155 10744 46164
rect 10692 46121 10701 46155
rect 10701 46121 10735 46155
rect 10735 46121 10744 46155
rect 10692 46112 10744 46121
rect 24492 46112 24544 46164
rect 24768 46112 24820 46164
rect 7656 46044 7708 46096
rect 9220 45976 9272 46028
rect 11888 46019 11940 46028
rect 11888 45985 11897 46019
rect 11897 45985 11931 46019
rect 11931 45985 11940 46019
rect 11888 45976 11940 45985
rect 12164 46019 12216 46028
rect 12164 45985 12173 46019
rect 12173 45985 12207 46019
rect 12207 45985 12216 46019
rect 12164 45976 12216 45985
rect 20168 46019 20220 46028
rect 20168 45985 20177 46019
rect 20177 45985 20211 46019
rect 20211 45985 20220 46019
rect 20168 45976 20220 45985
rect 20444 45976 20496 46028
rect 21364 46019 21416 46028
rect 21364 45985 21373 46019
rect 21373 45985 21407 46019
rect 21407 45985 21416 46019
rect 21364 45976 21416 45985
rect 21548 46019 21600 46028
rect 21548 45985 21557 46019
rect 21557 45985 21591 46019
rect 21591 45985 21600 46019
rect 21548 45976 21600 45985
rect 1308 45908 1360 45960
rect 8668 45908 8720 45960
rect 10968 45908 11020 45960
rect 20904 45908 20956 45960
rect 7380 45840 7432 45892
rect 11704 45840 11756 45892
rect 13912 45840 13964 45892
rect 11152 45815 11204 45824
rect 11152 45781 11161 45815
rect 11161 45781 11195 45815
rect 11195 45781 11204 45815
rect 11152 45772 11204 45781
rect 13636 45815 13688 45824
rect 13636 45781 13645 45815
rect 13645 45781 13679 45815
rect 13679 45781 13688 45815
rect 13636 45772 13688 45781
rect 15016 45772 15068 45824
rect 16396 45815 16448 45824
rect 16396 45781 16405 45815
rect 16405 45781 16439 45815
rect 16439 45781 16448 45815
rect 16396 45772 16448 45781
rect 17592 45772 17644 45824
rect 19064 45772 19116 45824
rect 19616 45840 19668 45892
rect 19892 45772 19944 45824
rect 20720 45772 20772 45824
rect 23480 45951 23532 45960
rect 23480 45917 23489 45951
rect 23489 45917 23523 45951
rect 23523 45917 23532 45951
rect 23480 45908 23532 45917
rect 24952 45772 25004 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 1308 45568 1360 45620
rect 19340 45568 19392 45620
rect 8760 45500 8812 45552
rect 9496 45543 9548 45552
rect 9496 45509 9505 45543
rect 9505 45509 9539 45543
rect 9539 45509 9548 45543
rect 9496 45500 9548 45509
rect 10876 45500 10928 45552
rect 15936 45500 15988 45552
rect 20536 45500 20588 45552
rect 21548 45500 21600 45552
rect 24032 45432 24084 45484
rect 24400 45432 24452 45484
rect 8760 45228 8812 45280
rect 10784 45296 10836 45348
rect 12256 45296 12308 45348
rect 10232 45228 10284 45280
rect 10876 45228 10928 45280
rect 12440 45228 12492 45280
rect 16304 45364 16356 45416
rect 18328 45364 18380 45416
rect 20076 45364 20128 45416
rect 14832 45228 14884 45280
rect 16120 45271 16172 45280
rect 16120 45237 16129 45271
rect 16129 45237 16163 45271
rect 16163 45237 16172 45271
rect 16120 45228 16172 45237
rect 20536 45271 20588 45280
rect 20536 45237 20545 45271
rect 20545 45237 20579 45271
rect 20579 45237 20588 45271
rect 20536 45228 20588 45237
rect 20812 45271 20864 45280
rect 20812 45237 20821 45271
rect 20821 45237 20855 45271
rect 20855 45237 20864 45271
rect 20812 45228 20864 45237
rect 22744 45364 22796 45416
rect 24492 45407 24544 45416
rect 24492 45373 24501 45407
rect 24501 45373 24535 45407
rect 24535 45373 24544 45407
rect 24492 45364 24544 45373
rect 22284 45228 22336 45280
rect 24032 45271 24084 45280
rect 24032 45237 24041 45271
rect 24041 45237 24075 45271
rect 24075 45237 24084 45271
rect 24032 45228 24084 45237
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 6368 45024 6420 45076
rect 11244 45024 11296 45076
rect 12532 45024 12584 45076
rect 15936 45024 15988 45076
rect 16764 45024 16816 45076
rect 17592 45024 17644 45076
rect 22100 45024 22152 45076
rect 22560 45024 22612 45076
rect 7288 44956 7340 45008
rect 10416 44888 10468 44940
rect 12624 44888 12676 44940
rect 13728 44888 13780 44940
rect 12440 44820 12492 44872
rect 13452 44820 13504 44872
rect 14832 44820 14884 44872
rect 16856 44888 16908 44940
rect 20536 44888 20588 44940
rect 19524 44863 19576 44872
rect 19524 44829 19533 44863
rect 19533 44829 19567 44863
rect 19567 44829 19576 44863
rect 19524 44820 19576 44829
rect 8576 44752 8628 44804
rect 11520 44795 11572 44804
rect 11520 44761 11529 44795
rect 11529 44761 11563 44795
rect 11563 44761 11572 44795
rect 11520 44752 11572 44761
rect 15660 44752 15712 44804
rect 15936 44752 15988 44804
rect 19800 44795 19852 44804
rect 19800 44761 19809 44795
rect 19809 44761 19843 44795
rect 19843 44761 19852 44795
rect 19800 44752 19852 44761
rect 21456 44888 21508 44940
rect 22284 44863 22336 44872
rect 22284 44829 22293 44863
rect 22293 44829 22327 44863
rect 22327 44829 22336 44863
rect 22284 44820 22336 44829
rect 24032 44820 24084 44872
rect 24584 44820 24636 44872
rect 25504 44820 25556 44872
rect 25780 44820 25832 44872
rect 22560 44795 22612 44804
rect 22560 44761 22569 44795
rect 22569 44761 22603 44795
rect 22603 44761 22612 44795
rect 22560 44752 22612 44761
rect 6460 44727 6512 44736
rect 6460 44693 6469 44727
rect 6469 44693 6503 44727
rect 6503 44693 6512 44727
rect 6460 44684 6512 44693
rect 7380 44684 7432 44736
rect 9680 44727 9732 44736
rect 9680 44693 9689 44727
rect 9689 44693 9723 44727
rect 9723 44693 9732 44727
rect 9680 44684 9732 44693
rect 15200 44684 15252 44736
rect 16672 44684 16724 44736
rect 16948 44684 17000 44736
rect 20628 44684 20680 44736
rect 22744 44684 22796 44736
rect 24492 44684 24544 44736
rect 25504 44727 25556 44736
rect 25504 44693 25513 44727
rect 25513 44693 25547 44727
rect 25547 44693 25556 44727
rect 25504 44684 25556 44693
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 5816 44523 5868 44532
rect 5816 44489 5825 44523
rect 5825 44489 5859 44523
rect 5859 44489 5868 44523
rect 5816 44480 5868 44489
rect 6736 44523 6788 44532
rect 6736 44489 6745 44523
rect 6745 44489 6779 44523
rect 6779 44489 6788 44523
rect 6736 44480 6788 44489
rect 7472 44523 7524 44532
rect 7472 44489 7481 44523
rect 7481 44489 7515 44523
rect 7515 44489 7524 44523
rect 7472 44480 7524 44489
rect 7840 44480 7892 44532
rect 9772 44480 9824 44532
rect 11152 44480 11204 44532
rect 15108 44480 15160 44532
rect 7104 44412 7156 44464
rect 10324 44412 10376 44464
rect 11612 44412 11664 44464
rect 12348 44412 12400 44464
rect 5356 44344 5408 44396
rect 6460 44344 6512 44396
rect 7380 44387 7432 44396
rect 7380 44353 7389 44387
rect 7389 44353 7423 44387
rect 7423 44353 7432 44387
rect 7380 44344 7432 44353
rect 7472 44344 7524 44396
rect 9404 44387 9456 44396
rect 9404 44353 9413 44387
rect 9413 44353 9447 44387
rect 9447 44353 9456 44387
rect 9404 44344 9456 44353
rect 11520 44344 11572 44396
rect 13360 44412 13412 44464
rect 15016 44412 15068 44464
rect 17592 44412 17644 44464
rect 19800 44480 19852 44532
rect 20444 44480 20496 44532
rect 21456 44480 21508 44532
rect 22560 44480 22612 44532
rect 20260 44412 20312 44464
rect 20536 44412 20588 44464
rect 22100 44412 22152 44464
rect 22652 44412 22704 44464
rect 24584 44412 24636 44464
rect 25320 44344 25372 44396
rect 10600 44276 10652 44328
rect 11152 44276 11204 44328
rect 12256 44208 12308 44260
rect 14188 44276 14240 44328
rect 16856 44319 16908 44328
rect 16856 44285 16865 44319
rect 16865 44285 16899 44319
rect 16899 44285 16908 44319
rect 16856 44276 16908 44285
rect 18972 44276 19024 44328
rect 19524 44319 19576 44328
rect 19524 44285 19533 44319
rect 19533 44285 19567 44319
rect 19567 44285 19576 44319
rect 19524 44276 19576 44285
rect 21180 44276 21232 44328
rect 22284 44319 22336 44328
rect 22284 44285 22293 44319
rect 22293 44285 22327 44319
rect 22327 44285 22336 44319
rect 22284 44276 22336 44285
rect 22652 44276 22704 44328
rect 23940 44276 23992 44328
rect 11520 44183 11572 44192
rect 11520 44149 11529 44183
rect 11529 44149 11563 44183
rect 11563 44149 11572 44183
rect 11520 44140 11572 44149
rect 13636 44140 13688 44192
rect 15016 44140 15068 44192
rect 18328 44140 18380 44192
rect 18788 44140 18840 44192
rect 22284 44140 22336 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 4712 43936 4764 43988
rect 8392 43979 8444 43988
rect 8392 43945 8401 43979
rect 8401 43945 8435 43979
rect 8435 43945 8444 43979
rect 8392 43936 8444 43945
rect 11612 43979 11664 43988
rect 11612 43945 11621 43979
rect 11621 43945 11655 43979
rect 11655 43945 11664 43979
rect 11612 43936 11664 43945
rect 16028 43800 16080 43852
rect 22192 43800 22244 43852
rect 23388 43800 23440 43852
rect 9036 43732 9088 43784
rect 9128 43775 9180 43784
rect 9128 43741 9137 43775
rect 9137 43741 9171 43775
rect 9171 43741 9180 43775
rect 9128 43732 9180 43741
rect 10784 43664 10836 43716
rect 11888 43664 11940 43716
rect 17408 43664 17460 43716
rect 18604 43664 18656 43716
rect 10324 43596 10376 43648
rect 10692 43596 10744 43648
rect 11244 43596 11296 43648
rect 17592 43596 17644 43648
rect 19524 43596 19576 43648
rect 20812 43596 20864 43648
rect 21732 43664 21784 43716
rect 21916 43596 21968 43648
rect 24584 43596 24636 43648
rect 25320 43639 25372 43648
rect 25320 43605 25329 43639
rect 25329 43605 25363 43639
rect 25363 43605 25372 43639
rect 25320 43596 25372 43605
rect 25504 43596 25556 43648
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 7748 43435 7800 43444
rect 7748 43401 7757 43435
rect 7757 43401 7791 43435
rect 7791 43401 7800 43435
rect 7748 43392 7800 43401
rect 8944 43392 8996 43444
rect 9496 43435 9548 43444
rect 9496 43401 9505 43435
rect 9505 43401 9539 43435
rect 9539 43401 9548 43435
rect 9496 43392 9548 43401
rect 10140 43392 10192 43444
rect 4620 43324 4672 43376
rect 12624 43367 12676 43376
rect 12624 43333 12633 43367
rect 12633 43333 12667 43367
rect 12667 43333 12676 43367
rect 12624 43324 12676 43333
rect 14464 43392 14516 43444
rect 16764 43435 16816 43444
rect 16764 43401 16773 43435
rect 16773 43401 16807 43435
rect 16807 43401 16816 43435
rect 16764 43392 16816 43401
rect 17500 43435 17552 43444
rect 17500 43401 17509 43435
rect 17509 43401 17543 43435
rect 17543 43401 17552 43435
rect 17500 43392 17552 43401
rect 20076 43435 20128 43444
rect 20076 43401 20085 43435
rect 20085 43401 20119 43435
rect 20119 43401 20128 43435
rect 20076 43392 20128 43401
rect 22376 43392 22428 43444
rect 15476 43324 15528 43376
rect 17592 43324 17644 43376
rect 20536 43324 20588 43376
rect 23572 43324 23624 43376
rect 24584 43324 24636 43376
rect 1308 43256 1360 43308
rect 6920 43256 6972 43308
rect 8484 43299 8536 43308
rect 8484 43265 8493 43299
rect 8493 43265 8527 43299
rect 8527 43265 8536 43299
rect 8484 43256 8536 43265
rect 8760 43256 8812 43308
rect 8944 43256 8996 43308
rect 9220 43188 9272 43240
rect 9588 43231 9640 43240
rect 9588 43197 9597 43231
rect 9597 43197 9631 43231
rect 9631 43197 9640 43231
rect 9588 43188 9640 43197
rect 10416 43256 10468 43308
rect 12348 43299 12400 43308
rect 12348 43265 12357 43299
rect 12357 43265 12391 43299
rect 12391 43265 12400 43299
rect 12348 43256 12400 43265
rect 13728 43256 13780 43308
rect 15384 43256 15436 43308
rect 21640 43256 21692 43308
rect 3976 43120 4028 43172
rect 11152 43120 11204 43172
rect 14740 43120 14792 43172
rect 15660 43188 15712 43240
rect 17224 43188 17276 43240
rect 18328 43231 18380 43240
rect 18328 43197 18337 43231
rect 18337 43197 18371 43231
rect 18371 43197 18380 43231
rect 18328 43188 18380 43197
rect 10784 43052 10836 43104
rect 12164 43052 12216 43104
rect 14648 43095 14700 43104
rect 14648 43061 14657 43095
rect 14657 43061 14691 43095
rect 14691 43061 14700 43095
rect 14648 43052 14700 43061
rect 15384 43052 15436 43104
rect 17040 43095 17092 43104
rect 17040 43061 17049 43095
rect 17049 43061 17083 43095
rect 17083 43061 17092 43095
rect 17040 43052 17092 43061
rect 20628 43188 20680 43240
rect 22652 43231 22704 43240
rect 22652 43197 22661 43231
rect 22661 43197 22695 43231
rect 22695 43197 22704 43231
rect 22652 43188 22704 43197
rect 23480 43188 23532 43240
rect 19708 43120 19760 43172
rect 19248 43052 19300 43104
rect 20536 43052 20588 43104
rect 20904 43052 20956 43104
rect 21640 43095 21692 43104
rect 21640 43061 21649 43095
rect 21649 43061 21683 43095
rect 21683 43061 21692 43095
rect 21640 43052 21692 43061
rect 24952 43052 25004 43104
rect 25504 43052 25556 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 8484 42848 8536 42900
rect 8944 42848 8996 42900
rect 12440 42780 12492 42832
rect 14556 42780 14608 42832
rect 4896 42712 4948 42764
rect 9128 42712 9180 42764
rect 12348 42712 12400 42764
rect 14832 42755 14884 42764
rect 14832 42721 14841 42755
rect 14841 42721 14875 42755
rect 14875 42721 14884 42755
rect 14832 42712 14884 42721
rect 15108 42712 15160 42764
rect 20352 42848 20404 42900
rect 21548 42848 21600 42900
rect 12164 42644 12216 42696
rect 12624 42644 12676 42696
rect 22008 42712 22060 42764
rect 22560 42712 22612 42764
rect 22192 42644 22244 42696
rect 8852 42576 8904 42628
rect 5264 42551 5316 42560
rect 5264 42517 5273 42551
rect 5273 42517 5307 42551
rect 5307 42517 5316 42551
rect 5264 42508 5316 42517
rect 8300 42508 8352 42560
rect 8760 42508 8812 42560
rect 8944 42551 8996 42560
rect 8944 42517 8953 42551
rect 8953 42517 8987 42551
rect 8987 42517 8996 42551
rect 8944 42508 8996 42517
rect 10416 42508 10468 42560
rect 10876 42508 10928 42560
rect 12440 42508 12492 42560
rect 12624 42508 12676 42560
rect 13728 42508 13780 42560
rect 15016 42508 15068 42560
rect 19800 42576 19852 42628
rect 20536 42576 20588 42628
rect 25136 42712 25188 42764
rect 23664 42644 23716 42696
rect 23756 42644 23808 42696
rect 24860 42644 24912 42696
rect 16764 42508 16816 42560
rect 19156 42508 19208 42560
rect 21272 42551 21324 42560
rect 21272 42517 21281 42551
rect 21281 42517 21315 42551
rect 21315 42517 21324 42551
rect 21272 42508 21324 42517
rect 21824 42551 21876 42560
rect 21824 42517 21833 42551
rect 21833 42517 21867 42551
rect 21867 42517 21876 42551
rect 21824 42508 21876 42517
rect 22192 42551 22244 42560
rect 22192 42517 22201 42551
rect 22201 42517 22235 42551
rect 22235 42517 22244 42551
rect 22192 42508 22244 42517
rect 24584 42576 24636 42628
rect 24860 42508 24912 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 4344 42347 4396 42356
rect 4344 42313 4353 42347
rect 4353 42313 4387 42347
rect 4387 42313 4396 42347
rect 4344 42304 4396 42313
rect 5080 42347 5132 42356
rect 5080 42313 5089 42347
rect 5089 42313 5123 42347
rect 5123 42313 5132 42347
rect 5080 42304 5132 42313
rect 4160 42236 4212 42288
rect 4252 42211 4304 42220
rect 4252 42177 4261 42211
rect 4261 42177 4295 42211
rect 4295 42177 4304 42211
rect 4252 42168 4304 42177
rect 8484 42304 8536 42356
rect 10232 42304 10284 42356
rect 11796 42347 11848 42356
rect 11796 42313 11805 42347
rect 11805 42313 11839 42347
rect 11839 42313 11848 42347
rect 11796 42304 11848 42313
rect 13452 42304 13504 42356
rect 15200 42304 15252 42356
rect 19616 42304 19668 42356
rect 6736 42168 6788 42220
rect 8852 42168 8904 42220
rect 6276 41964 6328 42016
rect 7748 42143 7800 42152
rect 7748 42109 7757 42143
rect 7757 42109 7791 42143
rect 7791 42109 7800 42143
rect 7748 42100 7800 42109
rect 10140 42143 10192 42152
rect 10140 42109 10149 42143
rect 10149 42109 10183 42143
rect 10183 42109 10192 42143
rect 10140 42100 10192 42109
rect 15108 42236 15160 42288
rect 20720 42347 20772 42356
rect 20720 42313 20729 42347
rect 20729 42313 20763 42347
rect 20763 42313 20772 42347
rect 20720 42304 20772 42313
rect 20904 42304 20956 42356
rect 23388 42304 23440 42356
rect 11152 42168 11204 42220
rect 15752 42211 15804 42220
rect 15752 42177 15761 42211
rect 15761 42177 15795 42211
rect 15795 42177 15804 42211
rect 15752 42168 15804 42177
rect 12440 42143 12492 42152
rect 12440 42109 12449 42143
rect 12449 42109 12483 42143
rect 12483 42109 12492 42143
rect 12440 42100 12492 42109
rect 12532 42100 12584 42152
rect 7196 42007 7248 42016
rect 7196 41973 7205 42007
rect 7205 41973 7239 42007
rect 7239 41973 7248 42007
rect 7196 41964 7248 41973
rect 7564 41964 7616 42016
rect 14188 42032 14240 42084
rect 9220 42007 9272 42016
rect 9220 41973 9229 42007
rect 9229 41973 9263 42007
rect 9263 41973 9272 42007
rect 9220 41964 9272 41973
rect 9312 41964 9364 42016
rect 10784 42007 10836 42016
rect 10784 41973 10793 42007
rect 10793 41973 10827 42007
rect 10827 41973 10836 42007
rect 10784 41964 10836 41973
rect 13452 41964 13504 42016
rect 13636 41964 13688 42016
rect 23756 42236 23808 42288
rect 24492 42236 24544 42288
rect 16396 42007 16448 42016
rect 16396 41973 16405 42007
rect 16405 41973 16439 42007
rect 16439 41973 16448 42007
rect 20628 42211 20680 42220
rect 20628 42177 20637 42211
rect 20637 42177 20671 42211
rect 20671 42177 20680 42211
rect 20628 42168 20680 42177
rect 19248 42100 19300 42152
rect 19984 42100 20036 42152
rect 21272 42100 21324 42152
rect 22284 42100 22336 42152
rect 22836 42143 22888 42152
rect 22836 42109 22845 42143
rect 22845 42109 22879 42143
rect 22879 42109 22888 42143
rect 23480 42143 23532 42152
rect 22836 42100 22888 42109
rect 23480 42109 23489 42143
rect 23489 42109 23523 42143
rect 23523 42109 23532 42143
rect 23480 42100 23532 42109
rect 25504 42100 25556 42152
rect 16396 41964 16448 41973
rect 18328 41964 18380 42016
rect 20260 42007 20312 42016
rect 20260 41973 20269 42007
rect 20269 41973 20303 42007
rect 20303 41973 20312 42007
rect 20260 41964 20312 41973
rect 24860 41964 24912 42016
rect 25044 41964 25096 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 5172 41803 5224 41812
rect 5172 41769 5181 41803
rect 5181 41769 5215 41803
rect 5215 41769 5224 41803
rect 5172 41760 5224 41769
rect 7748 41760 7800 41812
rect 6184 41624 6236 41676
rect 6736 41624 6788 41676
rect 8300 41760 8352 41812
rect 8852 41760 8904 41812
rect 11060 41760 11112 41812
rect 14464 41760 14516 41812
rect 16396 41760 16448 41812
rect 17316 41803 17368 41812
rect 17316 41769 17325 41803
rect 17325 41769 17359 41803
rect 17359 41769 17368 41803
rect 17316 41760 17368 41769
rect 9220 41692 9272 41744
rect 10876 41692 10928 41744
rect 15752 41692 15804 41744
rect 19340 41692 19392 41744
rect 21180 41803 21232 41812
rect 21180 41769 21189 41803
rect 21189 41769 21223 41803
rect 21223 41769 21232 41803
rect 21180 41760 21232 41769
rect 23204 41760 23256 41812
rect 25320 41760 25372 41812
rect 22560 41692 22612 41744
rect 25044 41692 25096 41744
rect 10232 41624 10284 41676
rect 10692 41624 10744 41676
rect 12348 41624 12400 41676
rect 12808 41624 12860 41676
rect 13636 41624 13688 41676
rect 15200 41624 15252 41676
rect 16120 41624 16172 41676
rect 18512 41624 18564 41676
rect 18972 41624 19024 41676
rect 19248 41624 19300 41676
rect 10324 41556 10376 41608
rect 11888 41556 11940 41608
rect 16672 41599 16724 41608
rect 16672 41565 16681 41599
rect 16681 41565 16715 41599
rect 16715 41565 16724 41599
rect 16672 41556 16724 41565
rect 17500 41556 17552 41608
rect 20904 41624 20956 41676
rect 22468 41624 22520 41676
rect 23296 41667 23348 41676
rect 23296 41633 23305 41667
rect 23305 41633 23339 41667
rect 23339 41633 23348 41667
rect 23296 41624 23348 41633
rect 23480 41624 23532 41676
rect 23572 41624 23624 41676
rect 25688 41624 25740 41676
rect 5724 41420 5776 41472
rect 10416 41488 10468 41540
rect 10784 41488 10836 41540
rect 18328 41488 18380 41540
rect 25320 41599 25372 41608
rect 25320 41565 25329 41599
rect 25329 41565 25363 41599
rect 25363 41565 25372 41599
rect 25320 41556 25372 41565
rect 19984 41488 20036 41540
rect 21088 41488 21140 41540
rect 22284 41488 22336 41540
rect 7012 41420 7064 41472
rect 11060 41463 11112 41472
rect 11060 41429 11069 41463
rect 11069 41429 11103 41463
rect 11103 41429 11112 41463
rect 11060 41420 11112 41429
rect 14188 41420 14240 41472
rect 16488 41420 16540 41472
rect 17316 41420 17368 41472
rect 18420 41420 18472 41472
rect 18880 41420 18932 41472
rect 22008 41463 22060 41472
rect 22008 41429 22017 41463
rect 22017 41429 22051 41463
rect 22051 41429 22060 41463
rect 22008 41420 22060 41429
rect 24584 41420 24636 41472
rect 25136 41463 25188 41472
rect 25136 41429 25145 41463
rect 25145 41429 25179 41463
rect 25179 41429 25188 41463
rect 25136 41420 25188 41429
rect 25320 41420 25372 41472
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 3332 41259 3384 41268
rect 3332 41225 3341 41259
rect 3341 41225 3375 41259
rect 3375 41225 3384 41259
rect 3332 41216 3384 41225
rect 11704 41259 11756 41268
rect 11704 41225 11713 41259
rect 11713 41225 11747 41259
rect 11747 41225 11756 41259
rect 11704 41216 11756 41225
rect 14924 41216 14976 41268
rect 1308 41080 1360 41132
rect 4620 41080 4672 41132
rect 9128 41148 9180 41200
rect 10876 41012 10928 41064
rect 1584 40919 1636 40928
rect 1584 40885 1593 40919
rect 1593 40885 1627 40919
rect 1627 40885 1636 40919
rect 1584 40876 1636 40885
rect 9956 40876 10008 40928
rect 10692 40919 10744 40928
rect 10692 40885 10701 40919
rect 10701 40885 10735 40919
rect 10735 40885 10744 40919
rect 10692 40876 10744 40885
rect 12072 41123 12124 41132
rect 12072 41089 12081 41123
rect 12081 41089 12115 41123
rect 12115 41089 12124 41123
rect 12072 41080 12124 41089
rect 13636 41123 13688 41132
rect 13636 41089 13645 41123
rect 13645 41089 13679 41123
rect 13679 41089 13688 41123
rect 13636 41080 13688 41089
rect 15016 41080 15068 41132
rect 19248 41216 19300 41268
rect 20168 41216 20220 41268
rect 21088 41216 21140 41268
rect 21548 41216 21600 41268
rect 22008 41259 22060 41268
rect 22008 41225 22017 41259
rect 22017 41225 22051 41259
rect 22051 41225 22060 41259
rect 22008 41216 22060 41225
rect 23480 41216 23532 41268
rect 18420 41148 18472 41200
rect 19892 41191 19944 41200
rect 19892 41157 19901 41191
rect 19901 41157 19935 41191
rect 19935 41157 19944 41191
rect 19892 41148 19944 41157
rect 12256 41055 12308 41064
rect 12256 41021 12265 41055
rect 12265 41021 12299 41055
rect 12299 41021 12308 41055
rect 12256 41012 12308 41021
rect 14004 41012 14056 41064
rect 15200 41012 15252 41064
rect 11336 40876 11388 40928
rect 12256 40876 12308 40928
rect 12624 40876 12676 40928
rect 15568 40876 15620 40928
rect 18604 41080 18656 41132
rect 21088 41123 21140 41132
rect 21088 41089 21097 41123
rect 21097 41089 21131 41123
rect 21131 41089 21140 41123
rect 21088 41080 21140 41089
rect 16764 41012 16816 41064
rect 19708 41012 19760 41064
rect 19984 41055 20036 41064
rect 19984 41021 19993 41055
rect 19993 41021 20027 41055
rect 20027 41021 20036 41055
rect 19984 41012 20036 41021
rect 20720 41012 20772 41064
rect 20996 41012 21048 41064
rect 22376 41148 22428 41200
rect 24492 41148 24544 41200
rect 25320 41123 25372 41132
rect 25320 41089 25329 41123
rect 25329 41089 25363 41123
rect 25363 41089 25372 41123
rect 25320 41080 25372 41089
rect 22836 41012 22888 41064
rect 23664 41012 23716 41064
rect 18420 40876 18472 40928
rect 18696 40876 18748 40928
rect 18880 40876 18932 40928
rect 19432 40919 19484 40928
rect 19432 40885 19441 40919
rect 19441 40885 19475 40919
rect 19475 40885 19484 40919
rect 19432 40876 19484 40885
rect 20904 40876 20956 40928
rect 21088 40876 21140 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 8300 40715 8352 40724
rect 8300 40681 8309 40715
rect 8309 40681 8343 40715
rect 8343 40681 8352 40715
rect 8300 40672 8352 40681
rect 9496 40672 9548 40724
rect 10232 40604 10284 40656
rect 11336 40604 11388 40656
rect 6552 40536 6604 40588
rect 6184 40511 6236 40520
rect 6184 40477 6193 40511
rect 6193 40477 6227 40511
rect 6227 40477 6236 40511
rect 6184 40468 6236 40477
rect 9404 40536 9456 40588
rect 9588 40536 9640 40588
rect 9680 40536 9732 40588
rect 14832 40672 14884 40724
rect 18604 40672 18656 40724
rect 22192 40672 22244 40724
rect 13360 40604 13412 40656
rect 13636 40536 13688 40588
rect 12716 40468 12768 40520
rect 15844 40604 15896 40656
rect 16948 40604 17000 40656
rect 15476 40536 15528 40588
rect 15752 40579 15804 40588
rect 15752 40545 15761 40579
rect 15761 40545 15795 40579
rect 15795 40545 15804 40579
rect 15752 40536 15804 40545
rect 17040 40536 17092 40588
rect 19800 40604 19852 40656
rect 20536 40604 20588 40656
rect 22008 40604 22060 40656
rect 24860 40672 24912 40724
rect 22468 40647 22520 40656
rect 22468 40613 22477 40647
rect 22477 40613 22511 40647
rect 22511 40613 22520 40647
rect 22468 40604 22520 40613
rect 22744 40604 22796 40656
rect 18880 40536 18932 40588
rect 21364 40579 21416 40588
rect 21364 40545 21373 40579
rect 21373 40545 21407 40579
rect 21407 40545 21416 40579
rect 21364 40536 21416 40545
rect 21456 40536 21508 40588
rect 23112 40604 23164 40656
rect 23848 40604 23900 40656
rect 8300 40400 8352 40452
rect 9220 40400 9272 40452
rect 9588 40443 9640 40452
rect 9588 40409 9597 40443
rect 9597 40409 9631 40443
rect 9631 40409 9640 40443
rect 9588 40400 9640 40409
rect 7104 40332 7156 40384
rect 7748 40332 7800 40384
rect 9404 40332 9456 40384
rect 11428 40375 11480 40384
rect 11428 40341 11437 40375
rect 11437 40341 11471 40375
rect 11471 40341 11480 40375
rect 11428 40332 11480 40341
rect 12440 40400 12492 40452
rect 14832 40332 14884 40384
rect 15200 40375 15252 40384
rect 15200 40341 15209 40375
rect 15209 40341 15243 40375
rect 15243 40341 15252 40375
rect 15200 40332 15252 40341
rect 17684 40400 17736 40452
rect 20168 40400 20220 40452
rect 17040 40375 17092 40384
rect 17040 40341 17049 40375
rect 17049 40341 17083 40375
rect 17083 40341 17092 40375
rect 17040 40332 17092 40341
rect 17316 40332 17368 40384
rect 18880 40332 18932 40384
rect 20996 40332 21048 40384
rect 21456 40400 21508 40452
rect 25412 40536 25464 40588
rect 22560 40468 22612 40520
rect 22928 40511 22980 40520
rect 22928 40477 22937 40511
rect 22937 40477 22971 40511
rect 22971 40477 22980 40511
rect 22928 40468 22980 40477
rect 23296 40468 23348 40520
rect 24032 40468 24084 40520
rect 24492 40468 24544 40520
rect 24768 40468 24820 40520
rect 21640 40400 21692 40452
rect 22192 40400 22244 40452
rect 23572 40400 23624 40452
rect 23296 40332 23348 40384
rect 24032 40375 24084 40384
rect 24032 40341 24041 40375
rect 24041 40341 24075 40375
rect 24075 40341 24084 40375
rect 24032 40332 24084 40341
rect 24216 40375 24268 40384
rect 24216 40341 24225 40375
rect 24225 40341 24259 40375
rect 24259 40341 24268 40375
rect 24216 40332 24268 40341
rect 24584 40332 24636 40384
rect 25320 40332 25372 40384
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 8668 40128 8720 40180
rect 9588 40128 9640 40180
rect 8760 40060 8812 40112
rect 9220 40060 9272 40112
rect 10968 40060 11020 40112
rect 8484 40035 8536 40044
rect 8484 40001 8493 40035
rect 8493 40001 8527 40035
rect 8527 40001 8536 40035
rect 8484 39992 8536 40001
rect 15016 40171 15068 40180
rect 15016 40137 15025 40171
rect 15025 40137 15059 40171
rect 15059 40137 15068 40171
rect 15016 40128 15068 40137
rect 15108 40128 15160 40180
rect 20628 40128 20680 40180
rect 21456 40128 21508 40180
rect 22100 40128 22152 40180
rect 15844 40060 15896 40112
rect 16948 40060 17000 40112
rect 12716 39992 12768 40044
rect 12808 39992 12860 40044
rect 14280 39992 14332 40044
rect 17132 39992 17184 40044
rect 20996 40060 21048 40112
rect 22008 40060 22060 40112
rect 22836 40060 22888 40112
rect 24032 40060 24084 40112
rect 7748 39967 7800 39976
rect 7748 39933 7757 39967
rect 7757 39933 7791 39967
rect 7791 39933 7800 39967
rect 7748 39924 7800 39933
rect 7840 39967 7892 39976
rect 7840 39933 7849 39967
rect 7849 39933 7883 39967
rect 7883 39933 7892 39967
rect 7840 39924 7892 39933
rect 9956 39924 10008 39976
rect 10968 39967 11020 39976
rect 10968 39933 10977 39967
rect 10977 39933 11011 39967
rect 11011 39933 11020 39967
rect 10968 39924 11020 39933
rect 15568 39924 15620 39976
rect 16028 39967 16080 39976
rect 16028 39933 16037 39967
rect 16037 39933 16071 39967
rect 16071 39933 16080 39967
rect 16028 39924 16080 39933
rect 18512 39924 18564 39976
rect 18788 39967 18840 39976
rect 18788 39933 18797 39967
rect 18797 39933 18831 39967
rect 18831 39933 18840 39967
rect 18788 39924 18840 39933
rect 19524 39924 19576 39976
rect 19800 39924 19852 39976
rect 20352 39967 20404 39976
rect 20352 39933 20361 39967
rect 20361 39933 20395 39967
rect 20395 39933 20404 39967
rect 20352 39924 20404 39933
rect 22560 39924 22612 39976
rect 24492 39924 24544 39976
rect 10784 39788 10836 39840
rect 14556 39788 14608 39840
rect 14740 39788 14792 39840
rect 19248 39788 19300 39840
rect 23756 39788 23808 39840
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 6552 39584 6604 39636
rect 7748 39584 7800 39636
rect 10876 39584 10928 39636
rect 12900 39584 12952 39636
rect 13084 39627 13136 39636
rect 13084 39593 13093 39627
rect 13093 39593 13127 39627
rect 13127 39593 13136 39627
rect 13084 39584 13136 39593
rect 14280 39584 14332 39636
rect 17040 39584 17092 39636
rect 22284 39584 22336 39636
rect 6736 39516 6788 39568
rect 8576 39516 8628 39568
rect 12716 39516 12768 39568
rect 16028 39516 16080 39568
rect 25136 39584 25188 39636
rect 6184 39448 6236 39500
rect 10232 39491 10284 39500
rect 10232 39457 10241 39491
rect 10241 39457 10275 39491
rect 10275 39457 10284 39491
rect 10232 39448 10284 39457
rect 8576 39380 8628 39432
rect 12624 39448 12676 39500
rect 12808 39448 12860 39500
rect 15660 39448 15712 39500
rect 17868 39448 17920 39500
rect 18604 39448 18656 39500
rect 18788 39448 18840 39500
rect 19432 39448 19484 39500
rect 20076 39491 20128 39500
rect 20076 39457 20085 39491
rect 20085 39457 20119 39491
rect 20119 39457 20128 39491
rect 20076 39448 20128 39457
rect 21364 39448 21416 39500
rect 22376 39448 22428 39500
rect 22560 39448 22612 39500
rect 12256 39380 12308 39432
rect 13084 39380 13136 39432
rect 5816 39244 5868 39296
rect 11520 39312 11572 39364
rect 15016 39312 15068 39364
rect 18604 39312 18656 39364
rect 7380 39244 7432 39296
rect 8300 39244 8352 39296
rect 12256 39244 12308 39296
rect 12716 39287 12768 39296
rect 12716 39253 12725 39287
rect 12725 39253 12759 39287
rect 12759 39253 12768 39287
rect 12716 39244 12768 39253
rect 13820 39287 13872 39296
rect 13820 39253 13829 39287
rect 13829 39253 13863 39287
rect 13863 39253 13872 39287
rect 13820 39244 13872 39253
rect 14740 39287 14792 39296
rect 14740 39253 14749 39287
rect 14749 39253 14783 39287
rect 14783 39253 14792 39287
rect 14740 39244 14792 39253
rect 15384 39244 15436 39296
rect 16028 39287 16080 39296
rect 16028 39253 16037 39287
rect 16037 39253 16071 39287
rect 16071 39253 16080 39287
rect 16028 39244 16080 39253
rect 18420 39244 18472 39296
rect 19524 39244 19576 39296
rect 20352 39380 20404 39432
rect 23480 39448 23532 39500
rect 23572 39380 23624 39432
rect 25044 39491 25096 39500
rect 25044 39457 25053 39491
rect 25053 39457 25087 39491
rect 25087 39457 25096 39491
rect 25044 39448 25096 39457
rect 25504 39448 25556 39500
rect 20444 39355 20496 39364
rect 20444 39321 20453 39355
rect 20453 39321 20487 39355
rect 20487 39321 20496 39355
rect 20444 39312 20496 39321
rect 22192 39312 22244 39364
rect 20996 39244 21048 39296
rect 24584 39287 24636 39296
rect 24584 39253 24593 39287
rect 24593 39253 24627 39287
rect 24627 39253 24636 39287
rect 24584 39244 24636 39253
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 7380 39083 7432 39092
rect 7380 39049 7389 39083
rect 7389 39049 7423 39083
rect 7423 39049 7432 39083
rect 7380 39040 7432 39049
rect 9220 39040 9272 39092
rect 9496 39083 9548 39092
rect 9496 39049 9505 39083
rect 9505 39049 9539 39083
rect 9539 39049 9548 39083
rect 9496 39040 9548 39049
rect 10968 39040 11020 39092
rect 12256 39040 12308 39092
rect 8668 38972 8720 39024
rect 11980 38972 12032 39024
rect 10784 38904 10836 38956
rect 12624 38972 12676 39024
rect 14740 39040 14792 39092
rect 15936 39040 15988 39092
rect 16028 39040 16080 39092
rect 20720 39083 20772 39092
rect 20720 39049 20729 39083
rect 20729 39049 20763 39083
rect 20763 39049 20772 39083
rect 20720 39040 20772 39049
rect 17776 38972 17828 39024
rect 20904 38972 20956 39024
rect 8852 38836 8904 38888
rect 9588 38879 9640 38888
rect 9588 38845 9597 38879
rect 9597 38845 9631 38879
rect 9631 38845 9640 38879
rect 9588 38836 9640 38845
rect 14280 38904 14332 38956
rect 19156 38904 19208 38956
rect 8484 38768 8536 38820
rect 14556 38836 14608 38888
rect 11152 38768 11204 38820
rect 9128 38743 9180 38752
rect 9128 38709 9137 38743
rect 9137 38709 9171 38743
rect 9171 38709 9180 38743
rect 9128 38700 9180 38709
rect 11704 38700 11756 38752
rect 15660 38836 15712 38888
rect 16120 38836 16172 38888
rect 16856 38879 16908 38888
rect 16856 38845 16865 38879
rect 16865 38845 16899 38879
rect 16899 38845 16908 38879
rect 16856 38836 16908 38845
rect 18420 38879 18472 38888
rect 18420 38845 18429 38879
rect 18429 38845 18463 38879
rect 18463 38845 18472 38879
rect 18420 38836 18472 38845
rect 19156 38768 19208 38820
rect 13912 38700 13964 38752
rect 15476 38700 15528 38752
rect 16028 38743 16080 38752
rect 16028 38709 16037 38743
rect 16037 38709 16071 38743
rect 16071 38709 16080 38743
rect 16028 38700 16080 38709
rect 16212 38700 16264 38752
rect 18236 38700 18288 38752
rect 18696 38700 18748 38752
rect 19892 38904 19944 38956
rect 23756 38972 23808 39024
rect 25780 38972 25832 39024
rect 24032 38904 24084 38956
rect 24216 38904 24268 38956
rect 24860 38904 24912 38956
rect 25320 38947 25372 38956
rect 25320 38913 25329 38947
rect 25329 38913 25363 38947
rect 25363 38913 25372 38947
rect 25320 38904 25372 38913
rect 20444 38836 20496 38888
rect 20904 38879 20956 38888
rect 20904 38845 20913 38879
rect 20913 38845 20947 38879
rect 20947 38845 20956 38879
rect 20904 38836 20956 38845
rect 22100 38879 22152 38888
rect 22100 38845 22109 38879
rect 22109 38845 22143 38879
rect 22143 38845 22152 38879
rect 22100 38836 22152 38845
rect 23388 38836 23440 38888
rect 21732 38768 21784 38820
rect 23572 38768 23624 38820
rect 25872 38768 25924 38820
rect 21272 38700 21324 38752
rect 23664 38700 23716 38752
rect 25136 38743 25188 38752
rect 25136 38709 25145 38743
rect 25145 38709 25179 38743
rect 25179 38709 25188 38743
rect 25136 38700 25188 38709
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 7564 38496 7616 38548
rect 11060 38496 11112 38548
rect 14188 38496 14240 38548
rect 14832 38496 14884 38548
rect 7656 38428 7708 38480
rect 6460 38360 6512 38412
rect 6920 38360 6972 38412
rect 7840 38360 7892 38412
rect 9128 38360 9180 38412
rect 1308 38292 1360 38344
rect 7380 38292 7432 38344
rect 8300 38292 8352 38344
rect 9220 38292 9272 38344
rect 10140 38428 10192 38480
rect 10876 38360 10928 38412
rect 11428 38360 11480 38412
rect 12716 38360 12768 38412
rect 16580 38496 16632 38548
rect 17776 38496 17828 38548
rect 18604 38428 18656 38480
rect 18236 38360 18288 38412
rect 19156 38496 19208 38548
rect 19340 38496 19392 38548
rect 20168 38496 20220 38548
rect 21456 38496 21508 38548
rect 21640 38496 21692 38548
rect 25596 38496 25648 38548
rect 18880 38428 18932 38480
rect 22376 38428 22428 38480
rect 22836 38428 22888 38480
rect 23388 38428 23440 38480
rect 14280 38292 14332 38344
rect 15200 38292 15252 38344
rect 15936 38335 15988 38344
rect 15936 38301 15945 38335
rect 15945 38301 15979 38335
rect 15979 38301 15988 38335
rect 15936 38292 15988 38301
rect 17776 38292 17828 38344
rect 19432 38360 19484 38412
rect 20260 38360 20312 38412
rect 21180 38403 21232 38412
rect 21180 38369 21189 38403
rect 21189 38369 21223 38403
rect 21223 38369 21232 38403
rect 21180 38360 21232 38369
rect 21916 38360 21968 38412
rect 22560 38403 22612 38412
rect 22560 38369 22569 38403
rect 22569 38369 22603 38403
rect 22603 38369 22612 38403
rect 22560 38360 22612 38369
rect 23664 38360 23716 38412
rect 23848 38360 23900 38412
rect 4068 38156 4120 38208
rect 8576 38224 8628 38276
rect 16304 38224 16356 38276
rect 18420 38224 18472 38276
rect 21640 38292 21692 38344
rect 19892 38267 19944 38276
rect 19892 38233 19901 38267
rect 19901 38233 19935 38267
rect 19935 38233 19944 38267
rect 19892 38224 19944 38233
rect 20444 38224 20496 38276
rect 23940 38292 23992 38344
rect 24952 38292 25004 38344
rect 8208 38156 8260 38208
rect 8392 38156 8444 38208
rect 10784 38199 10836 38208
rect 10784 38165 10793 38199
rect 10793 38165 10827 38199
rect 10827 38165 10836 38199
rect 10784 38156 10836 38165
rect 10876 38199 10928 38208
rect 10876 38165 10885 38199
rect 10885 38165 10919 38199
rect 10919 38165 10928 38199
rect 10876 38156 10928 38165
rect 12256 38199 12308 38208
rect 12256 38165 12265 38199
rect 12265 38165 12299 38199
rect 12299 38165 12308 38199
rect 12256 38156 12308 38165
rect 17224 38156 17276 38208
rect 17868 38156 17920 38208
rect 18512 38199 18564 38208
rect 18512 38165 18521 38199
rect 18521 38165 18555 38199
rect 18555 38165 18564 38199
rect 18512 38156 18564 38165
rect 19340 38156 19392 38208
rect 20628 38199 20680 38208
rect 20628 38165 20637 38199
rect 20637 38165 20671 38199
rect 20671 38165 20680 38199
rect 20628 38156 20680 38165
rect 20996 38199 21048 38208
rect 20996 38165 21005 38199
rect 21005 38165 21039 38199
rect 21039 38165 21048 38199
rect 20996 38156 21048 38165
rect 22284 38156 22336 38208
rect 23480 38224 23532 38276
rect 24308 38224 24360 38276
rect 23572 38199 23624 38208
rect 23572 38165 23581 38199
rect 23581 38165 23615 38199
rect 23615 38165 23624 38199
rect 23572 38156 23624 38165
rect 23664 38199 23716 38208
rect 23664 38165 23673 38199
rect 23673 38165 23707 38199
rect 23707 38165 23716 38199
rect 23664 38156 23716 38165
rect 23756 38156 23808 38208
rect 24676 38156 24728 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 5356 37952 5408 38004
rect 7840 37952 7892 38004
rect 8944 37952 8996 38004
rect 6920 37884 6972 37936
rect 7380 37884 7432 37936
rect 10784 37952 10836 38004
rect 12440 37952 12492 38004
rect 15476 37952 15528 38004
rect 16396 37995 16448 38004
rect 16396 37961 16405 37995
rect 16405 37961 16439 37995
rect 16439 37961 16448 37995
rect 16396 37952 16448 37961
rect 16856 37952 16908 38004
rect 18420 37952 18472 38004
rect 4988 37816 5040 37868
rect 18604 37884 18656 37936
rect 18880 37884 18932 37936
rect 19708 37952 19760 38004
rect 20352 37952 20404 38004
rect 24676 37952 24728 38004
rect 5816 37791 5868 37800
rect 5816 37757 5825 37791
rect 5825 37757 5859 37791
rect 5859 37757 5868 37791
rect 5816 37748 5868 37757
rect 6552 37791 6604 37800
rect 6552 37757 6561 37791
rect 6561 37757 6595 37791
rect 6595 37757 6604 37791
rect 6552 37748 6604 37757
rect 8484 37748 8536 37800
rect 6644 37612 6696 37664
rect 9956 37748 10008 37800
rect 13452 37748 13504 37800
rect 13544 37791 13596 37800
rect 13544 37757 13553 37791
rect 13553 37757 13587 37791
rect 13587 37757 13596 37791
rect 13544 37748 13596 37757
rect 15844 37816 15896 37868
rect 16120 37816 16172 37868
rect 18696 37859 18748 37868
rect 18696 37825 18705 37859
rect 18705 37825 18739 37859
rect 18739 37825 18748 37859
rect 18696 37816 18748 37825
rect 15200 37748 15252 37800
rect 15660 37791 15712 37800
rect 15660 37757 15669 37791
rect 15669 37757 15703 37791
rect 15703 37757 15712 37791
rect 15660 37748 15712 37757
rect 16028 37748 16080 37800
rect 12072 37680 12124 37732
rect 12164 37680 12216 37732
rect 16764 37680 16816 37732
rect 16948 37680 17000 37732
rect 17592 37748 17644 37800
rect 18328 37680 18380 37732
rect 18880 37680 18932 37732
rect 20168 37816 20220 37868
rect 20260 37816 20312 37868
rect 19708 37748 19760 37800
rect 20444 37748 20496 37800
rect 23480 37884 23532 37936
rect 23848 37927 23900 37936
rect 23848 37893 23857 37927
rect 23857 37893 23891 37927
rect 23891 37893 23900 37927
rect 23848 37884 23900 37893
rect 24308 37884 24360 37936
rect 22376 37859 22428 37868
rect 22376 37825 22385 37859
rect 22385 37825 22419 37859
rect 22419 37825 22428 37859
rect 22376 37816 22428 37825
rect 22744 37816 22796 37868
rect 23296 37816 23348 37868
rect 21364 37748 21416 37800
rect 21548 37680 21600 37732
rect 22836 37748 22888 37800
rect 22652 37680 22704 37732
rect 24492 37748 24544 37800
rect 10140 37612 10192 37664
rect 12808 37612 12860 37664
rect 15476 37612 15528 37664
rect 20352 37612 20404 37664
rect 22836 37612 22888 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 8576 37451 8628 37460
rect 8576 37417 8585 37451
rect 8585 37417 8619 37451
rect 8619 37417 8628 37451
rect 8576 37408 8628 37417
rect 10416 37451 10468 37460
rect 10416 37417 10425 37451
rect 10425 37417 10459 37451
rect 10459 37417 10468 37451
rect 10416 37408 10468 37417
rect 8484 37340 8536 37392
rect 12164 37340 12216 37392
rect 8300 37272 8352 37324
rect 9496 37272 9548 37324
rect 11244 37272 11296 37324
rect 11980 37272 12032 37324
rect 14004 37408 14056 37460
rect 14372 37451 14424 37460
rect 14372 37417 14381 37451
rect 14381 37417 14415 37451
rect 14415 37417 14424 37451
rect 14372 37408 14424 37417
rect 15568 37408 15620 37460
rect 14464 37340 14516 37392
rect 16304 37408 16356 37460
rect 18512 37408 18564 37460
rect 20720 37408 20772 37460
rect 23572 37408 23624 37460
rect 6552 37204 6604 37256
rect 10416 37204 10468 37256
rect 11704 37247 11756 37256
rect 11704 37213 11713 37247
rect 11713 37213 11747 37247
rect 11747 37213 11756 37247
rect 11704 37204 11756 37213
rect 13544 37204 13596 37256
rect 15016 37272 15068 37324
rect 15108 37272 15160 37324
rect 15200 37272 15252 37324
rect 15568 37272 15620 37324
rect 16396 37272 16448 37324
rect 17040 37340 17092 37392
rect 17776 37340 17828 37392
rect 18880 37340 18932 37392
rect 16764 37272 16816 37324
rect 24032 37340 24084 37392
rect 24216 37340 24268 37392
rect 14740 37204 14792 37256
rect 17776 37247 17828 37256
rect 17776 37213 17785 37247
rect 17785 37213 17819 37247
rect 17819 37213 17828 37247
rect 17776 37204 17828 37213
rect 20444 37272 20496 37324
rect 22100 37204 22152 37256
rect 7380 37136 7432 37188
rect 12808 37136 12860 37188
rect 14188 37179 14240 37188
rect 14188 37145 14197 37179
rect 14197 37145 14231 37179
rect 14231 37145 14240 37179
rect 14188 37136 14240 37145
rect 20076 37136 20128 37188
rect 20168 37179 20220 37188
rect 20168 37145 20177 37179
rect 20177 37145 20211 37179
rect 20211 37145 20220 37179
rect 20168 37136 20220 37145
rect 20720 37136 20772 37188
rect 24676 37136 24728 37188
rect 10508 37068 10560 37120
rect 12716 37068 12768 37120
rect 14740 37068 14792 37120
rect 14924 37111 14976 37120
rect 14924 37077 14933 37111
rect 14933 37077 14967 37111
rect 14967 37077 14976 37111
rect 14924 37068 14976 37077
rect 15108 37068 15160 37120
rect 15844 37068 15896 37120
rect 16304 37068 16356 37120
rect 18512 37111 18564 37120
rect 18512 37077 18521 37111
rect 18521 37077 18555 37111
rect 18555 37077 18564 37111
rect 18512 37068 18564 37077
rect 25320 37247 25372 37256
rect 25320 37213 25329 37247
rect 25329 37213 25363 37247
rect 25363 37213 25372 37247
rect 25320 37204 25372 37213
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 5540 36864 5592 36916
rect 6552 36864 6604 36916
rect 7472 36907 7524 36916
rect 7472 36873 7481 36907
rect 7481 36873 7515 36907
rect 7515 36873 7524 36907
rect 7472 36864 7524 36873
rect 8392 36864 8444 36916
rect 9036 36907 9088 36916
rect 9036 36873 9045 36907
rect 9045 36873 9079 36907
rect 9079 36873 9088 36907
rect 9036 36864 9088 36873
rect 9404 36864 9456 36916
rect 6920 36796 6972 36848
rect 7380 36796 7432 36848
rect 8668 36839 8720 36848
rect 8668 36805 8677 36839
rect 8677 36805 8711 36839
rect 8711 36805 8720 36839
rect 8668 36796 8720 36805
rect 10416 36796 10468 36848
rect 16028 36864 16080 36916
rect 17040 36907 17092 36916
rect 17040 36873 17049 36907
rect 17049 36873 17083 36907
rect 17083 36873 17092 36907
rect 17040 36864 17092 36873
rect 18512 36864 18564 36916
rect 19616 36864 19668 36916
rect 23848 36864 23900 36916
rect 14648 36796 14700 36848
rect 15200 36796 15252 36848
rect 15844 36796 15896 36848
rect 17776 36796 17828 36848
rect 19892 36796 19944 36848
rect 22652 36796 22704 36848
rect 23388 36796 23440 36848
rect 9128 36728 9180 36780
rect 9312 36728 9364 36780
rect 10600 36728 10652 36780
rect 12716 36728 12768 36780
rect 13452 36728 13504 36780
rect 14188 36728 14240 36780
rect 16764 36771 16816 36780
rect 16764 36737 16773 36771
rect 16773 36737 16807 36771
rect 16807 36737 16816 36771
rect 16764 36728 16816 36737
rect 5448 36660 5500 36712
rect 5816 36660 5868 36712
rect 6000 36660 6052 36712
rect 9588 36703 9640 36712
rect 9588 36669 9597 36703
rect 9597 36669 9631 36703
rect 9631 36669 9640 36703
rect 9588 36660 9640 36669
rect 10968 36703 11020 36712
rect 10968 36669 10977 36703
rect 10977 36669 11011 36703
rect 11011 36669 11020 36703
rect 10968 36660 11020 36669
rect 12808 36703 12860 36712
rect 12808 36669 12817 36703
rect 12817 36669 12851 36703
rect 12851 36669 12860 36703
rect 12808 36660 12860 36669
rect 13912 36703 13964 36712
rect 13912 36669 13921 36703
rect 13921 36669 13955 36703
rect 13955 36669 13964 36703
rect 13912 36660 13964 36669
rect 14372 36660 14424 36712
rect 15108 36703 15160 36712
rect 15108 36669 15117 36703
rect 15117 36669 15151 36703
rect 15151 36669 15160 36703
rect 15108 36660 15160 36669
rect 15844 36660 15896 36712
rect 19984 36728 20036 36780
rect 22100 36728 22152 36780
rect 22836 36771 22888 36780
rect 22836 36737 22845 36771
rect 22845 36737 22879 36771
rect 22879 36737 22888 36771
rect 22836 36728 22888 36737
rect 24216 36728 24268 36780
rect 24676 36728 24728 36780
rect 25320 36771 25372 36780
rect 25320 36737 25329 36771
rect 25329 36737 25363 36771
rect 25363 36737 25372 36771
rect 25320 36728 25372 36737
rect 18880 36660 18932 36712
rect 21916 36660 21968 36712
rect 24768 36660 24820 36712
rect 7656 36592 7708 36644
rect 11980 36592 12032 36644
rect 18972 36592 19024 36644
rect 10784 36524 10836 36576
rect 14464 36524 14516 36576
rect 14556 36567 14608 36576
rect 14556 36533 14565 36567
rect 14565 36533 14599 36567
rect 14599 36533 14608 36567
rect 14556 36524 14608 36533
rect 15844 36567 15896 36576
rect 15844 36533 15853 36567
rect 15853 36533 15887 36567
rect 15887 36533 15896 36567
rect 15844 36524 15896 36533
rect 17224 36524 17276 36576
rect 20076 36524 20128 36576
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 7012 36320 7064 36372
rect 7840 36320 7892 36372
rect 11888 36320 11940 36372
rect 12440 36320 12492 36372
rect 12532 36320 12584 36372
rect 15384 36320 15436 36372
rect 15844 36320 15896 36372
rect 23664 36320 23716 36372
rect 11520 36252 11572 36304
rect 15752 36252 15804 36304
rect 7472 36184 7524 36236
rect 1768 36159 1820 36168
rect 1768 36125 1777 36159
rect 1777 36125 1811 36159
rect 1811 36125 1820 36159
rect 1768 36116 1820 36125
rect 7656 36116 7708 36168
rect 12716 36184 12768 36236
rect 13820 36227 13872 36236
rect 13820 36193 13829 36227
rect 13829 36193 13863 36227
rect 13863 36193 13872 36227
rect 13820 36184 13872 36193
rect 14832 36227 14884 36236
rect 14832 36193 14841 36227
rect 14841 36193 14875 36227
rect 14875 36193 14884 36227
rect 14832 36184 14884 36193
rect 17500 36184 17552 36236
rect 19432 36295 19484 36304
rect 19432 36261 19441 36295
rect 19441 36261 19475 36295
rect 19475 36261 19484 36295
rect 19432 36252 19484 36261
rect 20996 36252 21048 36304
rect 21824 36252 21876 36304
rect 10140 36116 10192 36168
rect 12440 36116 12492 36168
rect 12716 36048 12768 36100
rect 21272 36227 21324 36236
rect 21272 36193 21281 36227
rect 21281 36193 21315 36227
rect 21315 36193 21324 36227
rect 21272 36184 21324 36193
rect 3424 35980 3476 36032
rect 7748 35980 7800 36032
rect 10324 35980 10376 36032
rect 12440 36023 12492 36032
rect 12440 35989 12449 36023
rect 12449 35989 12483 36023
rect 12483 35989 12492 36023
rect 12440 35980 12492 35989
rect 12624 35980 12676 36032
rect 14648 36023 14700 36032
rect 14648 35989 14657 36023
rect 14657 35989 14691 36023
rect 14691 35989 14700 36023
rect 14648 35980 14700 35989
rect 15752 36023 15804 36032
rect 15752 35989 15761 36023
rect 15761 35989 15795 36023
rect 15795 35989 15804 36023
rect 15752 35980 15804 35989
rect 15844 35980 15896 36032
rect 21180 36116 21232 36168
rect 23756 36227 23808 36236
rect 23756 36193 23765 36227
rect 23765 36193 23799 36227
rect 23799 36193 23808 36227
rect 23756 36184 23808 36193
rect 24492 36184 24544 36236
rect 25320 36159 25372 36168
rect 25320 36125 25329 36159
rect 25329 36125 25363 36159
rect 25363 36125 25372 36159
rect 25320 36116 25372 36125
rect 22100 36048 22152 36100
rect 25136 36048 25188 36100
rect 20352 35980 20404 36032
rect 20444 35980 20496 36032
rect 21088 35980 21140 36032
rect 23296 36023 23348 36032
rect 23296 35989 23305 36023
rect 23305 35989 23339 36023
rect 23339 35989 23348 36023
rect 23296 35980 23348 35989
rect 23664 36023 23716 36032
rect 23664 35989 23673 36023
rect 23673 35989 23707 36023
rect 23707 35989 23716 36023
rect 23664 35980 23716 35989
rect 23756 35980 23808 36032
rect 24400 35980 24452 36032
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 5540 35776 5592 35828
rect 6000 35819 6052 35828
rect 6000 35785 6009 35819
rect 6009 35785 6043 35819
rect 6043 35785 6052 35819
rect 6000 35776 6052 35785
rect 6920 35776 6972 35828
rect 8668 35708 8720 35760
rect 5816 35572 5868 35624
rect 9588 35572 9640 35624
rect 8852 35436 8904 35488
rect 9772 35436 9824 35488
rect 13544 35776 13596 35828
rect 14004 35776 14056 35828
rect 14372 35776 14424 35828
rect 14648 35776 14700 35828
rect 17776 35776 17828 35828
rect 24400 35776 24452 35828
rect 14096 35708 14148 35760
rect 17132 35708 17184 35760
rect 17868 35751 17920 35760
rect 17868 35717 17877 35751
rect 17877 35717 17911 35751
rect 17911 35717 17920 35751
rect 17868 35708 17920 35717
rect 18420 35708 18472 35760
rect 20536 35708 20588 35760
rect 23940 35708 23992 35760
rect 19248 35640 19300 35692
rect 21088 35640 21140 35692
rect 22192 35640 22244 35692
rect 22836 35640 22888 35692
rect 10968 35572 11020 35624
rect 13820 35572 13872 35624
rect 13636 35504 13688 35556
rect 10232 35479 10284 35488
rect 10232 35445 10241 35479
rect 10241 35445 10275 35479
rect 10275 35445 10284 35479
rect 10232 35436 10284 35445
rect 15936 35436 15988 35488
rect 18604 35572 18656 35624
rect 22744 35572 22796 35624
rect 23388 35615 23440 35624
rect 23388 35581 23397 35615
rect 23397 35581 23431 35615
rect 23431 35581 23440 35615
rect 23388 35572 23440 35581
rect 23940 35572 23992 35624
rect 25412 35572 25464 35624
rect 21548 35504 21600 35556
rect 17960 35436 18012 35488
rect 19800 35479 19852 35488
rect 19800 35445 19809 35479
rect 19809 35445 19843 35479
rect 19843 35445 19852 35479
rect 19800 35436 19852 35445
rect 20996 35436 21048 35488
rect 22376 35436 22428 35488
rect 22836 35436 22888 35488
rect 23480 35436 23532 35488
rect 25320 35436 25372 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 7656 35232 7708 35284
rect 8668 35232 8720 35284
rect 8760 35232 8812 35284
rect 10600 35232 10652 35284
rect 15660 35232 15712 35284
rect 8576 35164 8628 35216
rect 5540 35096 5592 35148
rect 6092 35139 6144 35148
rect 6092 35105 6101 35139
rect 6101 35105 6135 35139
rect 6135 35105 6144 35139
rect 6092 35096 6144 35105
rect 9772 35096 9824 35148
rect 12348 35164 12400 35216
rect 13452 35164 13504 35216
rect 11060 35096 11112 35148
rect 15752 35096 15804 35148
rect 14556 35028 14608 35080
rect 17868 35232 17920 35284
rect 18328 35232 18380 35284
rect 18420 35232 18472 35284
rect 20904 35232 20956 35284
rect 21088 35232 21140 35284
rect 22376 35232 22428 35284
rect 17960 35096 18012 35148
rect 18328 35096 18380 35148
rect 20168 35096 20220 35148
rect 23020 35096 23072 35148
rect 23940 35096 23992 35148
rect 24216 35096 24268 35148
rect 22192 35028 22244 35080
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 6920 34960 6972 35012
rect 8668 34960 8720 35012
rect 10140 34892 10192 34944
rect 15568 34892 15620 34944
rect 19616 34960 19668 35012
rect 20996 34960 21048 35012
rect 21180 34935 21232 34944
rect 21180 34901 21189 34935
rect 21189 34901 21223 34935
rect 21223 34901 21232 34935
rect 21180 34892 21232 34901
rect 22560 35003 22612 35012
rect 22560 34969 22569 35003
rect 22569 34969 22603 35003
rect 22603 34969 22612 35003
rect 22560 34960 22612 34969
rect 23020 34960 23072 35012
rect 23388 34892 23440 34944
rect 24952 34892 25004 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 8760 34688 8812 34740
rect 6000 34620 6052 34672
rect 6920 34620 6972 34672
rect 7288 34620 7340 34672
rect 9772 34688 9824 34740
rect 6092 34552 6144 34604
rect 8852 34595 8904 34604
rect 8852 34561 8868 34595
rect 8868 34561 8902 34595
rect 8902 34561 8904 34595
rect 8852 34552 8904 34561
rect 12808 34688 12860 34740
rect 13728 34688 13780 34740
rect 14004 34688 14056 34740
rect 14188 34688 14240 34740
rect 19800 34688 19852 34740
rect 20720 34688 20772 34740
rect 21640 34688 21692 34740
rect 22100 34688 22152 34740
rect 22468 34731 22520 34740
rect 22468 34697 22477 34731
rect 22477 34697 22511 34731
rect 22511 34697 22520 34731
rect 22468 34688 22520 34697
rect 22744 34688 22796 34740
rect 24676 34688 24728 34740
rect 6920 34484 6972 34536
rect 10416 34484 10468 34536
rect 10968 34484 11020 34536
rect 16212 34620 16264 34672
rect 20260 34620 20312 34672
rect 15568 34552 15620 34604
rect 18512 34552 18564 34604
rect 20628 34552 20680 34604
rect 21640 34552 21692 34604
rect 24032 34552 24084 34604
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 5264 34416 5316 34468
rect 5632 34416 5684 34468
rect 10232 34416 10284 34468
rect 13820 34484 13872 34536
rect 14832 34484 14884 34536
rect 15844 34416 15896 34468
rect 19800 34416 19852 34468
rect 22100 34416 22152 34468
rect 23572 34484 23624 34536
rect 23664 34527 23716 34536
rect 23664 34493 23673 34527
rect 23673 34493 23707 34527
rect 23707 34493 23716 34527
rect 23664 34484 23716 34493
rect 23848 34416 23900 34468
rect 9864 34348 9916 34400
rect 10968 34348 11020 34400
rect 11980 34391 12032 34400
rect 11980 34357 12010 34391
rect 12010 34357 12032 34391
rect 11980 34348 12032 34357
rect 20720 34391 20772 34400
rect 20720 34357 20729 34391
rect 20729 34357 20763 34391
rect 20763 34357 20772 34391
rect 20720 34348 20772 34357
rect 22008 34391 22060 34400
rect 22008 34357 22017 34391
rect 22017 34357 22051 34391
rect 22051 34357 22060 34391
rect 22008 34348 22060 34357
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 7288 34144 7340 34196
rect 9128 34187 9180 34196
rect 9128 34153 9137 34187
rect 9137 34153 9171 34187
rect 9171 34153 9180 34187
rect 9128 34144 9180 34153
rect 10692 34144 10744 34196
rect 13820 34144 13872 34196
rect 18420 34144 18472 34196
rect 19432 34144 19484 34196
rect 25320 34187 25372 34196
rect 25320 34153 25329 34187
rect 25329 34153 25363 34187
rect 25363 34153 25372 34187
rect 25320 34144 25372 34153
rect 25412 34187 25464 34196
rect 25412 34153 25421 34187
rect 25421 34153 25455 34187
rect 25455 34153 25464 34187
rect 25412 34144 25464 34153
rect 5540 34051 5592 34060
rect 5540 34017 5549 34051
rect 5549 34017 5583 34051
rect 5583 34017 5592 34051
rect 5540 34008 5592 34017
rect 5816 34008 5868 34060
rect 9220 34008 9272 34060
rect 10416 33983 10468 33992
rect 10416 33949 10425 33983
rect 10425 33949 10459 33983
rect 10459 33949 10468 33983
rect 10416 33940 10468 33949
rect 12072 33940 12124 33992
rect 13360 34008 13412 34060
rect 20260 34076 20312 34128
rect 20536 34076 20588 34128
rect 15936 34051 15988 34060
rect 15936 34017 15945 34051
rect 15945 34017 15979 34051
rect 15979 34017 15988 34051
rect 15936 34008 15988 34017
rect 17776 34008 17828 34060
rect 21180 34008 21232 34060
rect 22284 34008 22336 34060
rect 23388 34008 23440 34060
rect 13636 33940 13688 33992
rect 14096 33983 14148 33992
rect 7288 33872 7340 33924
rect 7656 33872 7708 33924
rect 9680 33872 9732 33924
rect 7380 33804 7432 33856
rect 8484 33804 8536 33856
rect 12532 33872 12584 33924
rect 14096 33949 14105 33983
rect 14105 33949 14139 33983
rect 14139 33949 14148 33983
rect 14096 33940 14148 33949
rect 17868 33940 17920 33992
rect 19432 33940 19484 33992
rect 19708 33940 19760 33992
rect 21732 33940 21784 33992
rect 12072 33804 12124 33856
rect 12808 33804 12860 33856
rect 13176 33804 13228 33856
rect 14740 33872 14792 33924
rect 13636 33804 13688 33856
rect 13912 33804 13964 33856
rect 14004 33804 14056 33856
rect 19248 33804 19300 33856
rect 20076 33872 20128 33924
rect 20904 33872 20956 33924
rect 24584 33940 24636 33992
rect 25136 33872 25188 33924
rect 20628 33847 20680 33856
rect 20628 33813 20637 33847
rect 20637 33813 20671 33847
rect 20671 33813 20680 33847
rect 20628 33804 20680 33813
rect 21456 33847 21508 33856
rect 21456 33813 21465 33847
rect 21465 33813 21499 33847
rect 21499 33813 21508 33847
rect 21456 33804 21508 33813
rect 22468 33804 22520 33856
rect 24584 33847 24636 33856
rect 24584 33813 24593 33847
rect 24593 33813 24627 33847
rect 24627 33813 24636 33847
rect 24584 33804 24636 33813
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 7288 33600 7340 33652
rect 10324 33600 10376 33652
rect 10784 33600 10836 33652
rect 12716 33600 12768 33652
rect 13820 33600 13872 33652
rect 11796 33532 11848 33584
rect 14004 33532 14056 33584
rect 1308 33464 1360 33516
rect 11612 33464 11664 33516
rect 12440 33464 12492 33516
rect 12624 33464 12676 33516
rect 12716 33464 12768 33516
rect 13176 33464 13228 33516
rect 14556 33600 14608 33652
rect 15936 33600 15988 33652
rect 17868 33600 17920 33652
rect 5356 33439 5408 33448
rect 5356 33405 5365 33439
rect 5365 33405 5399 33439
rect 5399 33405 5408 33439
rect 5356 33396 5408 33405
rect 9772 33439 9824 33448
rect 9772 33405 9781 33439
rect 9781 33405 9815 33439
rect 9815 33405 9824 33439
rect 9772 33396 9824 33405
rect 8300 33328 8352 33380
rect 11428 33396 11480 33448
rect 15936 33464 15988 33516
rect 18328 33532 18380 33584
rect 19616 33600 19668 33652
rect 20628 33643 20680 33652
rect 20628 33609 20637 33643
rect 20637 33609 20671 33643
rect 20671 33609 20680 33643
rect 20628 33600 20680 33609
rect 21456 33600 21508 33652
rect 23664 33532 23716 33584
rect 21272 33464 21324 33516
rect 22192 33464 22244 33516
rect 13544 33439 13596 33448
rect 13544 33405 13553 33439
rect 13553 33405 13587 33439
rect 13587 33405 13596 33439
rect 13544 33396 13596 33405
rect 16304 33396 16356 33448
rect 12624 33328 12676 33380
rect 19432 33328 19484 33380
rect 19892 33328 19944 33380
rect 3516 33260 3568 33312
rect 7196 33260 7248 33312
rect 10600 33260 10652 33312
rect 13452 33260 13504 33312
rect 15844 33303 15896 33312
rect 15844 33269 15853 33303
rect 15853 33269 15887 33303
rect 15887 33269 15896 33303
rect 15844 33260 15896 33269
rect 20996 33396 21048 33448
rect 23756 33439 23808 33448
rect 23756 33405 23765 33439
rect 23765 33405 23799 33439
rect 23799 33405 23808 33439
rect 23756 33396 23808 33405
rect 24216 33396 24268 33448
rect 25412 33532 25464 33584
rect 23480 33328 23532 33380
rect 21180 33260 21232 33312
rect 21272 33303 21324 33312
rect 21272 33269 21281 33303
rect 21281 33269 21315 33303
rect 21315 33269 21324 33303
rect 21272 33260 21324 33269
rect 21364 33260 21416 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 7748 33056 7800 33108
rect 9312 33056 9364 33108
rect 10600 33099 10652 33108
rect 10600 33065 10609 33099
rect 10609 33065 10643 33099
rect 10643 33065 10652 33099
rect 10600 33056 10652 33065
rect 10876 33056 10928 33108
rect 9680 32988 9732 33040
rect 15108 33056 15160 33108
rect 17408 33099 17460 33108
rect 13636 32988 13688 33040
rect 5540 32920 5592 32972
rect 7472 32920 7524 32972
rect 7288 32852 7340 32904
rect 8300 32920 8352 32972
rect 9864 32920 9916 32972
rect 11152 32920 11204 32972
rect 11520 32920 11572 32972
rect 14464 32920 14516 32972
rect 14832 32963 14884 32972
rect 14832 32929 14841 32963
rect 14841 32929 14875 32963
rect 14875 32929 14884 32963
rect 14832 32920 14884 32929
rect 9772 32895 9824 32904
rect 9772 32861 9781 32895
rect 9781 32861 9815 32895
rect 9815 32861 9824 32895
rect 9772 32852 9824 32861
rect 15476 32920 15528 32972
rect 17408 33065 17417 33099
rect 17417 33065 17451 33099
rect 17451 33065 17460 33099
rect 17408 33056 17460 33065
rect 20904 33056 20956 33108
rect 21180 33056 21232 33108
rect 21824 33056 21876 33108
rect 23940 33056 23992 33108
rect 17868 32988 17920 33040
rect 16948 32920 17000 32972
rect 22560 32988 22612 33040
rect 21456 32963 21508 32972
rect 21456 32929 21465 32963
rect 21465 32929 21499 32963
rect 21499 32929 21508 32963
rect 21456 32920 21508 32929
rect 21548 32963 21600 32972
rect 21548 32929 21557 32963
rect 21557 32929 21591 32963
rect 21591 32929 21600 32963
rect 21548 32920 21600 32929
rect 20996 32852 21048 32904
rect 22376 32895 22428 32904
rect 22376 32861 22385 32895
rect 22385 32861 22419 32895
rect 22419 32861 22428 32895
rect 22376 32852 22428 32861
rect 22744 32895 22796 32904
rect 22744 32861 22753 32895
rect 22753 32861 22787 32895
rect 22787 32861 22796 32895
rect 22744 32852 22796 32861
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 7748 32784 7800 32836
rect 11704 32784 11756 32836
rect 7840 32759 7892 32768
rect 7840 32725 7849 32759
rect 7849 32725 7883 32759
rect 7883 32725 7892 32759
rect 7840 32716 7892 32725
rect 9496 32716 9548 32768
rect 10600 32716 10652 32768
rect 11888 32716 11940 32768
rect 14004 32716 14056 32768
rect 14464 32716 14516 32768
rect 14648 32759 14700 32768
rect 14648 32725 14657 32759
rect 14657 32725 14691 32759
rect 14691 32725 14700 32759
rect 14648 32716 14700 32725
rect 16120 32759 16172 32768
rect 16120 32725 16129 32759
rect 16129 32725 16163 32759
rect 16163 32725 16172 32759
rect 16120 32716 16172 32725
rect 16212 32716 16264 32768
rect 20904 32716 20956 32768
rect 21088 32716 21140 32768
rect 21272 32716 21324 32768
rect 24124 32716 24176 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 4620 32555 4672 32564
rect 4620 32521 4629 32555
rect 4629 32521 4663 32555
rect 4663 32521 4672 32555
rect 4620 32512 4672 32521
rect 4988 32555 5040 32564
rect 4988 32521 4997 32555
rect 4997 32521 5031 32555
rect 5031 32521 5040 32555
rect 4988 32512 5040 32521
rect 5356 32555 5408 32564
rect 5356 32521 5365 32555
rect 5365 32521 5399 32555
rect 5399 32521 5408 32555
rect 5356 32512 5408 32521
rect 7840 32512 7892 32564
rect 4896 32444 4948 32496
rect 5540 32444 5592 32496
rect 7288 32444 7340 32496
rect 8484 32512 8536 32564
rect 9680 32512 9732 32564
rect 14648 32512 14700 32564
rect 12256 32444 12308 32496
rect 16212 32512 16264 32564
rect 17684 32512 17736 32564
rect 6184 32376 6236 32428
rect 14556 32419 14608 32428
rect 14556 32385 14565 32419
rect 14565 32385 14599 32419
rect 14599 32385 14608 32419
rect 14556 32376 14608 32385
rect 15936 32376 15988 32428
rect 17224 32419 17276 32428
rect 17224 32385 17233 32419
rect 17233 32385 17267 32419
rect 17267 32385 17276 32419
rect 17224 32376 17276 32385
rect 5448 32308 5500 32360
rect 7472 32308 7524 32360
rect 9864 32351 9916 32360
rect 9864 32317 9873 32351
rect 9873 32317 9907 32351
rect 9907 32317 9916 32351
rect 9864 32308 9916 32317
rect 11060 32308 11112 32360
rect 12164 32308 12216 32360
rect 11980 32240 12032 32292
rect 16212 32308 16264 32360
rect 17868 32308 17920 32360
rect 16304 32283 16356 32292
rect 16304 32249 16313 32283
rect 16313 32249 16347 32283
rect 16347 32249 16356 32283
rect 18696 32444 18748 32496
rect 21272 32512 21324 32564
rect 21916 32555 21968 32564
rect 21916 32521 21925 32555
rect 21925 32521 21959 32555
rect 21959 32521 21968 32555
rect 21916 32512 21968 32521
rect 24492 32512 24544 32564
rect 24768 32512 24820 32564
rect 18696 32351 18748 32360
rect 18696 32317 18705 32351
rect 18705 32317 18739 32351
rect 18739 32317 18748 32351
rect 18696 32308 18748 32317
rect 19524 32308 19576 32360
rect 21088 32419 21140 32428
rect 21088 32385 21097 32419
rect 21097 32385 21131 32419
rect 21131 32385 21140 32419
rect 21088 32376 21140 32385
rect 21640 32376 21692 32428
rect 24032 32444 24084 32496
rect 21548 32308 21600 32360
rect 23204 32308 23256 32360
rect 16304 32240 16356 32249
rect 10968 32172 11020 32224
rect 14556 32172 14608 32224
rect 15200 32172 15252 32224
rect 16856 32215 16908 32224
rect 16856 32181 16865 32215
rect 16865 32181 16899 32215
rect 16899 32181 16908 32215
rect 16856 32172 16908 32181
rect 17684 32172 17736 32224
rect 18604 32172 18656 32224
rect 20076 32215 20128 32224
rect 20076 32181 20085 32215
rect 20085 32181 20119 32215
rect 20119 32181 20128 32215
rect 20076 32172 20128 32181
rect 21364 32172 21416 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 8300 31968 8352 32020
rect 9680 32011 9732 32020
rect 9680 31977 9710 32011
rect 9710 31977 9732 32011
rect 9680 31968 9732 31977
rect 10140 31968 10192 32020
rect 8392 31900 8444 31952
rect 11152 32011 11204 32020
rect 11152 31977 11161 32011
rect 11161 31977 11195 32011
rect 11195 31977 11204 32011
rect 11152 31968 11204 31977
rect 11612 31968 11664 32020
rect 6184 31875 6236 31884
rect 6184 31841 6193 31875
rect 6193 31841 6227 31875
rect 6227 31841 6236 31875
rect 6184 31832 6236 31841
rect 6920 31832 6972 31884
rect 8484 31832 8536 31884
rect 5724 31628 5776 31680
rect 8484 31628 8536 31680
rect 9404 31807 9456 31816
rect 9404 31773 9413 31807
rect 9413 31773 9447 31807
rect 9447 31773 9456 31807
rect 9404 31764 9456 31773
rect 11060 31764 11112 31816
rect 11336 31764 11388 31816
rect 10968 31696 11020 31748
rect 11612 31764 11664 31816
rect 12072 31764 12124 31816
rect 13728 31832 13780 31884
rect 16580 31832 16632 31884
rect 21180 31968 21232 32020
rect 24216 31968 24268 32020
rect 25136 32011 25188 32020
rect 25136 31977 25145 32011
rect 25145 31977 25179 32011
rect 25179 31977 25188 32011
rect 25136 31968 25188 31977
rect 18420 31832 18472 31884
rect 17592 31696 17644 31748
rect 18880 31764 18932 31816
rect 18972 31764 19024 31816
rect 9772 31628 9824 31680
rect 13912 31671 13964 31680
rect 13912 31637 13921 31671
rect 13921 31637 13955 31671
rect 13955 31637 13964 31671
rect 13912 31628 13964 31637
rect 14832 31628 14884 31680
rect 16764 31671 16816 31680
rect 16764 31637 16773 31671
rect 16773 31637 16807 31671
rect 16807 31637 16816 31671
rect 16764 31628 16816 31637
rect 16948 31628 17000 31680
rect 18788 31628 18840 31680
rect 18972 31628 19024 31680
rect 19616 31832 19668 31884
rect 23388 31900 23440 31952
rect 21364 31832 21416 31884
rect 23480 31832 23532 31884
rect 20444 31764 20496 31816
rect 21824 31764 21876 31816
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 20536 31696 20588 31748
rect 21180 31696 21232 31748
rect 19156 31628 19208 31680
rect 20628 31671 20680 31680
rect 20628 31637 20637 31671
rect 20637 31637 20671 31671
rect 20671 31637 20680 31671
rect 20628 31628 20680 31637
rect 20904 31628 20956 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 7656 31424 7708 31476
rect 8668 31467 8720 31476
rect 8668 31433 8677 31467
rect 8677 31433 8711 31467
rect 8711 31433 8720 31467
rect 8668 31424 8720 31433
rect 9864 31424 9916 31476
rect 13360 31424 13412 31476
rect 13544 31424 13596 31476
rect 8392 31356 8444 31408
rect 15936 31424 15988 31476
rect 17592 31467 17644 31476
rect 17592 31433 17601 31467
rect 17601 31433 17635 31467
rect 17635 31433 17644 31467
rect 17592 31424 17644 31433
rect 18512 31424 18564 31476
rect 21456 31424 21508 31476
rect 21824 31424 21876 31476
rect 23296 31424 23348 31476
rect 1952 31288 2004 31340
rect 7840 31331 7892 31340
rect 7840 31297 7849 31331
rect 7849 31297 7883 31331
rect 7883 31297 7892 31331
rect 7840 31288 7892 31297
rect 1308 31220 1360 31272
rect 5632 31220 5684 31272
rect 8944 31288 8996 31340
rect 8116 31263 8168 31272
rect 8116 31229 8125 31263
rect 8125 31229 8159 31263
rect 8159 31229 8168 31263
rect 8116 31220 8168 31229
rect 8484 31220 8536 31272
rect 15108 31356 15160 31408
rect 9404 31220 9456 31272
rect 7380 31152 7432 31204
rect 13268 31220 13320 31272
rect 14372 31220 14424 31272
rect 18328 31288 18380 31340
rect 17776 31263 17828 31272
rect 17776 31229 17785 31263
rect 17785 31229 17819 31263
rect 17819 31229 17828 31263
rect 17776 31220 17828 31229
rect 19892 31399 19944 31408
rect 19892 31365 19901 31399
rect 19901 31365 19935 31399
rect 19935 31365 19944 31399
rect 19892 31356 19944 31365
rect 21640 31356 21692 31408
rect 24216 31356 24268 31408
rect 24400 31424 24452 31476
rect 25320 31331 25372 31340
rect 25320 31297 25329 31331
rect 25329 31297 25363 31331
rect 25363 31297 25372 31331
rect 25320 31288 25372 31297
rect 16488 31152 16540 31204
rect 19064 31220 19116 31272
rect 19984 31263 20036 31272
rect 19984 31229 19993 31263
rect 19993 31229 20027 31263
rect 20027 31229 20036 31263
rect 19984 31220 20036 31229
rect 20536 31220 20588 31272
rect 22100 31220 22152 31272
rect 22192 31263 22244 31272
rect 22192 31229 22201 31263
rect 22201 31229 22235 31263
rect 22235 31229 22244 31263
rect 22192 31220 22244 31229
rect 24952 31220 25004 31272
rect 14464 31084 14516 31136
rect 14648 31127 14700 31136
rect 14648 31093 14657 31127
rect 14657 31093 14691 31127
rect 14691 31093 14700 31127
rect 14648 31084 14700 31093
rect 17132 31127 17184 31136
rect 17132 31093 17141 31127
rect 17141 31093 17175 31127
rect 17175 31093 17184 31127
rect 17132 31084 17184 31093
rect 19892 31084 19944 31136
rect 22284 31084 22336 31136
rect 23572 31084 23624 31136
rect 24400 31127 24452 31136
rect 24400 31093 24409 31127
rect 24409 31093 24443 31127
rect 24443 31093 24452 31127
rect 24400 31084 24452 31093
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 8116 30880 8168 30932
rect 11612 30855 11664 30864
rect 1584 30744 1636 30796
rect 7840 30744 7892 30796
rect 9404 30744 9456 30796
rect 10600 30744 10652 30796
rect 11612 30821 11621 30855
rect 11621 30821 11655 30855
rect 11655 30821 11664 30855
rect 11612 30812 11664 30821
rect 12532 30880 12584 30932
rect 15936 30923 15988 30932
rect 15936 30889 15945 30923
rect 15945 30889 15979 30923
rect 15979 30889 15988 30923
rect 15936 30880 15988 30889
rect 15200 30744 15252 30796
rect 16948 30744 17000 30796
rect 11244 30676 11296 30728
rect 13544 30676 13596 30728
rect 18604 30880 18656 30932
rect 19248 30880 19300 30932
rect 20444 30923 20496 30932
rect 20444 30889 20453 30923
rect 20453 30889 20487 30923
rect 20487 30889 20496 30923
rect 20444 30880 20496 30889
rect 23480 30880 23532 30932
rect 23848 30880 23900 30932
rect 25320 30880 25372 30932
rect 19984 30787 20036 30796
rect 19984 30753 19993 30787
rect 19993 30753 20027 30787
rect 20027 30753 20036 30787
rect 19984 30744 20036 30753
rect 20168 30744 20220 30796
rect 20260 30676 20312 30728
rect 22284 30676 22336 30728
rect 22468 30676 22520 30728
rect 25504 30676 25556 30728
rect 3792 30608 3844 30660
rect 6276 30608 6328 30660
rect 16580 30608 16632 30660
rect 18512 30608 18564 30660
rect 18696 30608 18748 30660
rect 8484 30583 8536 30592
rect 8484 30549 8493 30583
rect 8493 30549 8527 30583
rect 8527 30549 8536 30583
rect 8484 30540 8536 30549
rect 11336 30583 11388 30592
rect 11336 30549 11345 30583
rect 11345 30549 11379 30583
rect 11379 30549 11388 30583
rect 11336 30540 11388 30549
rect 17868 30540 17920 30592
rect 19432 30583 19484 30592
rect 19432 30549 19441 30583
rect 19441 30549 19475 30583
rect 19475 30549 19484 30583
rect 19432 30540 19484 30549
rect 22284 30540 22336 30592
rect 23480 30540 23532 30592
rect 25044 30540 25096 30592
rect 25136 30583 25188 30592
rect 25136 30549 25145 30583
rect 25145 30549 25179 30583
rect 25179 30549 25188 30583
rect 25136 30540 25188 30549
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 11796 30336 11848 30388
rect 16948 30336 17000 30388
rect 18328 30336 18380 30388
rect 18696 30336 18748 30388
rect 20444 30336 20496 30388
rect 25136 30336 25188 30388
rect 8392 30268 8444 30320
rect 11244 30268 11296 30320
rect 16396 30268 16448 30320
rect 10048 30132 10100 30184
rect 10600 30132 10652 30184
rect 10692 30064 10744 30116
rect 10416 30039 10468 30048
rect 10416 30005 10425 30039
rect 10425 30005 10459 30039
rect 10459 30005 10468 30039
rect 10416 29996 10468 30005
rect 11888 29996 11940 30048
rect 14372 30200 14424 30252
rect 14464 30243 14516 30252
rect 14464 30209 14473 30243
rect 14473 30209 14507 30243
rect 14507 30209 14516 30243
rect 14464 30200 14516 30209
rect 15844 30200 15896 30252
rect 17408 30200 17460 30252
rect 17868 30200 17920 30252
rect 16212 30175 16264 30184
rect 16212 30141 16221 30175
rect 16221 30141 16255 30175
rect 16255 30141 16264 30175
rect 16212 30132 16264 30141
rect 17224 30132 17276 30184
rect 19064 30200 19116 30252
rect 23572 30268 23624 30320
rect 24216 30268 24268 30320
rect 22192 30200 22244 30252
rect 14372 29996 14424 30048
rect 17592 30039 17644 30048
rect 17592 30005 17601 30039
rect 17601 30005 17635 30039
rect 17635 30005 17644 30039
rect 17592 29996 17644 30005
rect 19800 30132 19852 30184
rect 23756 30132 23808 30184
rect 18328 30064 18380 30116
rect 21088 30064 21140 30116
rect 19064 29996 19116 30048
rect 19248 29996 19300 30048
rect 21824 29996 21876 30048
rect 24216 29996 24268 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 4252 29792 4304 29844
rect 7656 29792 7708 29844
rect 7748 29792 7800 29844
rect 9496 29835 9548 29844
rect 9496 29801 9505 29835
rect 9505 29801 9539 29835
rect 9539 29801 9548 29835
rect 9496 29792 9548 29801
rect 10416 29792 10468 29844
rect 12992 29792 13044 29844
rect 16028 29835 16080 29844
rect 16028 29801 16037 29835
rect 16037 29801 16071 29835
rect 16071 29801 16080 29835
rect 16028 29792 16080 29801
rect 16488 29792 16540 29844
rect 16580 29792 16632 29844
rect 21732 29792 21784 29844
rect 6368 29724 6420 29776
rect 9312 29724 9364 29776
rect 9588 29724 9640 29776
rect 11336 29724 11388 29776
rect 4068 29656 4120 29708
rect 6920 29656 6972 29708
rect 9680 29656 9732 29708
rect 7840 29588 7892 29640
rect 17316 29724 17368 29776
rect 17592 29724 17644 29776
rect 14924 29656 14976 29708
rect 18788 29699 18840 29708
rect 18788 29665 18797 29699
rect 18797 29665 18831 29699
rect 18831 29665 18840 29699
rect 18788 29656 18840 29665
rect 21180 29656 21232 29708
rect 11796 29631 11848 29640
rect 11796 29597 11805 29631
rect 11805 29597 11839 29631
rect 11839 29597 11848 29631
rect 11796 29588 11848 29597
rect 12808 29588 12860 29640
rect 13728 29631 13780 29640
rect 13728 29597 13737 29631
rect 13737 29597 13771 29631
rect 13771 29597 13780 29631
rect 13728 29588 13780 29597
rect 17040 29588 17092 29640
rect 20720 29588 20772 29640
rect 3884 29520 3936 29572
rect 6092 29563 6144 29572
rect 6092 29529 6101 29563
rect 6101 29529 6135 29563
rect 6135 29529 6144 29563
rect 6092 29520 6144 29529
rect 7104 29520 7156 29572
rect 7380 29452 7432 29504
rect 9588 29520 9640 29572
rect 9956 29563 10008 29572
rect 9956 29529 9965 29563
rect 9965 29529 9999 29563
rect 9999 29529 10008 29563
rect 9956 29520 10008 29529
rect 12992 29563 13044 29572
rect 12992 29529 13001 29563
rect 13001 29529 13035 29563
rect 13035 29529 13044 29563
rect 12992 29520 13044 29529
rect 14740 29563 14792 29572
rect 14740 29529 14749 29563
rect 14749 29529 14783 29563
rect 14783 29529 14792 29563
rect 14740 29520 14792 29529
rect 16396 29520 16448 29572
rect 7656 29452 7708 29504
rect 10692 29452 10744 29504
rect 10784 29452 10836 29504
rect 11888 29495 11940 29504
rect 11888 29461 11897 29495
rect 11897 29461 11931 29495
rect 11931 29461 11940 29495
rect 11888 29452 11940 29461
rect 15108 29452 15160 29504
rect 17592 29520 17644 29572
rect 19340 29520 19392 29572
rect 22560 29656 22612 29708
rect 23388 29699 23440 29708
rect 23388 29665 23397 29699
rect 23397 29665 23431 29699
rect 23431 29665 23440 29699
rect 23388 29656 23440 29665
rect 23756 29656 23808 29708
rect 22008 29588 22060 29640
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 21456 29520 21508 29572
rect 17500 29452 17552 29504
rect 19064 29452 19116 29504
rect 20352 29452 20404 29504
rect 20904 29495 20956 29504
rect 20904 29461 20913 29495
rect 20913 29461 20947 29495
rect 20947 29461 20956 29495
rect 20904 29452 20956 29461
rect 21548 29495 21600 29504
rect 21548 29461 21557 29495
rect 21557 29461 21591 29495
rect 21591 29461 21600 29495
rect 21548 29452 21600 29461
rect 21732 29520 21784 29572
rect 23848 29520 23900 29572
rect 22836 29452 22888 29504
rect 23296 29495 23348 29504
rect 23296 29461 23305 29495
rect 23305 29461 23339 29495
rect 23339 29461 23348 29495
rect 23296 29452 23348 29461
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 7656 29248 7708 29300
rect 9036 29180 9088 29232
rect 9772 29291 9824 29300
rect 9772 29257 9781 29291
rect 9781 29257 9815 29291
rect 9815 29257 9824 29291
rect 9772 29248 9824 29257
rect 11244 29248 11296 29300
rect 15660 29248 15712 29300
rect 17224 29291 17276 29300
rect 17224 29257 17233 29291
rect 17233 29257 17267 29291
rect 17267 29257 17276 29291
rect 17224 29248 17276 29257
rect 17500 29248 17552 29300
rect 17592 29248 17644 29300
rect 19524 29248 19576 29300
rect 6552 29044 6604 29096
rect 9404 29044 9456 29096
rect 9036 28976 9088 29028
rect 9772 29044 9824 29096
rect 13728 29112 13780 29164
rect 14096 29155 14148 29164
rect 14096 29121 14105 29155
rect 14105 29121 14139 29155
rect 14139 29121 14148 29155
rect 14096 29112 14148 29121
rect 14188 29155 14240 29164
rect 14188 29121 14197 29155
rect 14197 29121 14231 29155
rect 14231 29121 14240 29155
rect 14188 29112 14240 29121
rect 15568 29180 15620 29232
rect 16304 29180 16356 29232
rect 18328 29180 18380 29232
rect 20812 29248 20864 29300
rect 20904 29248 20956 29300
rect 23848 29248 23900 29300
rect 25320 29291 25372 29300
rect 25320 29257 25329 29291
rect 25329 29257 25363 29291
rect 25363 29257 25372 29291
rect 25320 29248 25372 29257
rect 25504 29291 25556 29300
rect 25504 29257 25513 29291
rect 25513 29257 25547 29291
rect 25547 29257 25556 29291
rect 25504 29248 25556 29257
rect 22468 29180 22520 29232
rect 24584 29180 24636 29232
rect 10876 28976 10928 29028
rect 13084 29044 13136 29096
rect 13268 29044 13320 29096
rect 13912 29044 13964 29096
rect 14280 29044 14332 29096
rect 14648 29044 14700 29096
rect 15200 29044 15252 29096
rect 16396 29112 16448 29164
rect 21456 29112 21508 29164
rect 24124 29155 24176 29164
rect 17408 29087 17460 29096
rect 17408 29053 17417 29087
rect 17417 29053 17451 29087
rect 17451 29053 17460 29087
rect 17408 29044 17460 29053
rect 17592 29044 17644 29096
rect 17776 29044 17828 29096
rect 13452 28976 13504 29028
rect 16028 28976 16080 29028
rect 16948 28976 17000 29028
rect 20168 29044 20220 29096
rect 24124 29121 24133 29155
rect 24133 29121 24167 29155
rect 24167 29121 24176 29155
rect 24124 29112 24176 29121
rect 23572 29044 23624 29096
rect 8668 28908 8720 28960
rect 16120 28908 16172 28960
rect 19064 28976 19116 29028
rect 19616 28976 19668 29028
rect 20812 28976 20864 29028
rect 20904 28976 20956 29028
rect 23296 28976 23348 29028
rect 23480 28976 23532 29028
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 14096 28704 14148 28756
rect 14740 28704 14792 28756
rect 21272 28704 21324 28756
rect 21456 28704 21508 28756
rect 24308 28704 24360 28756
rect 21180 28679 21232 28688
rect 21180 28645 21189 28679
rect 21189 28645 21223 28679
rect 21223 28645 21232 28679
rect 21180 28636 21232 28645
rect 1308 28568 1360 28620
rect 3424 28568 3476 28620
rect 5908 28611 5960 28620
rect 5908 28577 5917 28611
rect 5917 28577 5951 28611
rect 5951 28577 5960 28611
rect 5908 28568 5960 28577
rect 6552 28611 6604 28620
rect 6552 28577 6561 28611
rect 6561 28577 6595 28611
rect 6595 28577 6604 28611
rect 6552 28568 6604 28577
rect 1768 28543 1820 28552
rect 1768 28509 1777 28543
rect 1777 28509 1811 28543
rect 1811 28509 1820 28543
rect 1768 28500 1820 28509
rect 9864 28568 9916 28620
rect 11336 28568 11388 28620
rect 13360 28611 13412 28620
rect 13360 28577 13369 28611
rect 13369 28577 13403 28611
rect 13403 28577 13412 28611
rect 13360 28568 13412 28577
rect 13636 28568 13688 28620
rect 16212 28611 16264 28620
rect 16212 28577 16221 28611
rect 16221 28577 16255 28611
rect 16255 28577 16264 28611
rect 16212 28568 16264 28577
rect 17132 28568 17184 28620
rect 17776 28611 17828 28620
rect 17776 28577 17785 28611
rect 17785 28577 17819 28611
rect 17819 28577 17828 28611
rect 17776 28568 17828 28577
rect 22008 28568 22060 28620
rect 22836 28568 22888 28620
rect 9404 28500 9456 28552
rect 9956 28500 10008 28552
rect 15568 28500 15620 28552
rect 16028 28543 16080 28552
rect 16028 28509 16037 28543
rect 16037 28509 16071 28543
rect 16071 28509 16080 28543
rect 16028 28500 16080 28509
rect 16856 28500 16908 28552
rect 18604 28500 18656 28552
rect 3976 28432 4028 28484
rect 12532 28432 12584 28484
rect 13084 28432 13136 28484
rect 19800 28432 19852 28484
rect 21456 28475 21508 28484
rect 21456 28441 21465 28475
rect 21465 28441 21499 28475
rect 21499 28441 21508 28475
rect 21456 28432 21508 28441
rect 24216 28432 24268 28484
rect 24860 28432 24912 28484
rect 9036 28364 9088 28416
rect 9588 28364 9640 28416
rect 12808 28364 12860 28416
rect 13176 28407 13228 28416
rect 13176 28373 13185 28407
rect 13185 28373 13219 28407
rect 13219 28373 13228 28407
rect 13176 28364 13228 28373
rect 14004 28364 14056 28416
rect 14280 28407 14332 28416
rect 14280 28373 14289 28407
rect 14289 28373 14323 28407
rect 14323 28373 14332 28407
rect 14280 28364 14332 28373
rect 14740 28407 14792 28416
rect 14740 28373 14749 28407
rect 14749 28373 14783 28407
rect 14783 28373 14792 28407
rect 14740 28364 14792 28373
rect 15200 28364 15252 28416
rect 15752 28364 15804 28416
rect 16948 28364 17000 28416
rect 18420 28364 18472 28416
rect 24584 28407 24636 28416
rect 24584 28373 24593 28407
rect 24593 28373 24627 28407
rect 24627 28373 24636 28407
rect 24584 28364 24636 28373
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 1952 28160 2004 28212
rect 3792 28160 3844 28212
rect 5908 28160 5960 28212
rect 9036 28092 9088 28144
rect 13176 28160 13228 28212
rect 15660 28160 15712 28212
rect 15936 28203 15988 28212
rect 15936 28169 15945 28203
rect 15945 28169 15979 28203
rect 15979 28169 15988 28203
rect 15936 28160 15988 28169
rect 18328 28203 18380 28212
rect 18328 28169 18337 28203
rect 18337 28169 18371 28203
rect 18371 28169 18380 28203
rect 18328 28160 18380 28169
rect 20260 28160 20312 28212
rect 16120 28092 16172 28144
rect 3424 28024 3476 28076
rect 3608 28067 3660 28076
rect 3608 28033 3652 28067
rect 3652 28033 3660 28067
rect 3608 28024 3660 28033
rect 9588 28024 9640 28076
rect 12532 28024 12584 28076
rect 13360 28024 13412 28076
rect 15200 28024 15252 28076
rect 15844 28024 15896 28076
rect 15936 28024 15988 28076
rect 18512 28092 18564 28144
rect 18788 28092 18840 28144
rect 24308 28160 24360 28212
rect 24676 28135 24728 28144
rect 24676 28101 24685 28135
rect 24685 28101 24719 28135
rect 24719 28101 24728 28135
rect 24676 28092 24728 28101
rect 8576 27999 8628 28008
rect 8576 27965 8585 27999
rect 8585 27965 8619 27999
rect 8619 27965 8628 27999
rect 8576 27956 8628 27965
rect 8668 27956 8720 28008
rect 16028 27999 16080 28008
rect 16028 27965 16037 27999
rect 16037 27965 16071 27999
rect 16071 27965 16080 27999
rect 16028 27956 16080 27965
rect 11796 27888 11848 27940
rect 9956 27820 10008 27872
rect 12624 27820 12676 27872
rect 13084 27863 13136 27872
rect 13084 27829 13093 27863
rect 13093 27829 13127 27863
rect 13127 27829 13136 27863
rect 13084 27820 13136 27829
rect 13360 27863 13412 27872
rect 13360 27829 13369 27863
rect 13369 27829 13403 27863
rect 13403 27829 13412 27863
rect 13360 27820 13412 27829
rect 14740 27820 14792 27872
rect 15292 27888 15344 27940
rect 19524 28024 19576 28076
rect 22008 28067 22060 28076
rect 22008 28033 22017 28067
rect 22017 28033 22051 28067
rect 22051 28033 22060 28067
rect 22008 28024 22060 28033
rect 18512 27999 18564 28008
rect 18512 27965 18521 27999
rect 18521 27965 18555 27999
rect 18555 27965 18564 27999
rect 18512 27956 18564 27965
rect 18972 27956 19024 28008
rect 19064 27956 19116 28008
rect 19616 27956 19668 28008
rect 19984 27956 20036 28008
rect 24676 27956 24728 28008
rect 15568 27863 15620 27872
rect 15568 27829 15577 27863
rect 15577 27829 15611 27863
rect 15611 27829 15620 27863
rect 15568 27820 15620 27829
rect 16028 27820 16080 27872
rect 16396 27820 16448 27872
rect 21364 27888 21416 27940
rect 18972 27820 19024 27872
rect 19064 27863 19116 27872
rect 19064 27829 19073 27863
rect 19073 27829 19107 27863
rect 19107 27829 19116 27863
rect 19064 27820 19116 27829
rect 22100 27820 22152 27872
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 9864 27616 9916 27668
rect 18328 27616 18380 27668
rect 18788 27616 18840 27668
rect 7840 27548 7892 27600
rect 14188 27548 14240 27600
rect 15384 27548 15436 27600
rect 15844 27548 15896 27600
rect 16212 27548 16264 27600
rect 20996 27616 21048 27668
rect 24216 27659 24268 27668
rect 24216 27625 24225 27659
rect 24225 27625 24259 27659
rect 24259 27625 24268 27659
rect 24216 27616 24268 27625
rect 21088 27548 21140 27600
rect 24308 27548 24360 27600
rect 6552 27480 6604 27532
rect 7012 27480 7064 27532
rect 9036 27480 9088 27532
rect 12808 27480 12860 27532
rect 17868 27480 17920 27532
rect 9956 27412 10008 27464
rect 10968 27412 11020 27464
rect 13360 27412 13412 27464
rect 14556 27412 14608 27464
rect 7012 27344 7064 27396
rect 11428 27387 11480 27396
rect 11428 27353 11437 27387
rect 11437 27353 11471 27387
rect 11471 27353 11480 27387
rect 11428 27344 11480 27353
rect 13084 27344 13136 27396
rect 13912 27344 13964 27396
rect 15200 27344 15252 27396
rect 15384 27344 15436 27396
rect 17224 27344 17276 27396
rect 19524 27344 19576 27396
rect 11704 27276 11756 27328
rect 12900 27319 12952 27328
rect 12900 27285 12909 27319
rect 12909 27285 12943 27319
rect 12943 27285 12952 27319
rect 12900 27276 12952 27285
rect 13360 27276 13412 27328
rect 13544 27276 13596 27328
rect 15016 27276 15068 27328
rect 15844 27276 15896 27328
rect 18604 27276 18656 27328
rect 20536 27480 20588 27532
rect 21916 27523 21968 27532
rect 21916 27489 21925 27523
rect 21925 27489 21959 27523
rect 21959 27489 21968 27523
rect 21916 27480 21968 27489
rect 23388 27480 23440 27532
rect 20444 27412 20496 27464
rect 24492 27412 24544 27464
rect 22192 27387 22244 27396
rect 22192 27353 22201 27387
rect 22201 27353 22235 27387
rect 22235 27353 22244 27387
rect 22192 27344 22244 27353
rect 25228 27344 25280 27396
rect 23112 27276 23164 27328
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 3884 27072 3936 27124
rect 3332 26936 3384 26988
rect 3516 26936 3568 26988
rect 4344 26868 4396 26920
rect 7104 27004 7156 27056
rect 10508 27047 10560 27056
rect 10508 27013 10517 27047
rect 10517 27013 10551 27047
rect 10551 27013 10560 27047
rect 10508 27004 10560 27013
rect 6552 26979 6604 26988
rect 6552 26945 6561 26979
rect 6561 26945 6595 26979
rect 6595 26945 6604 26979
rect 6552 26936 6604 26945
rect 9128 26979 9180 26988
rect 9128 26945 9137 26979
rect 9137 26945 9171 26979
rect 9171 26945 9180 26979
rect 9128 26936 9180 26945
rect 7840 26868 7892 26920
rect 8944 26868 8996 26920
rect 9404 26911 9456 26920
rect 9404 26877 9413 26911
rect 9413 26877 9447 26911
rect 9447 26877 9456 26911
rect 9404 26868 9456 26877
rect 11060 27072 11112 27124
rect 11520 27072 11572 27124
rect 11612 27072 11664 27124
rect 12532 27072 12584 27124
rect 12900 27072 12952 27124
rect 11336 27004 11388 27056
rect 13084 27004 13136 27056
rect 15108 27072 15160 27124
rect 10968 26936 11020 26988
rect 13912 26936 13964 26988
rect 14556 26936 14608 26988
rect 11612 26868 11664 26920
rect 12808 26911 12860 26920
rect 12808 26877 12817 26911
rect 12817 26877 12851 26911
rect 12851 26877 12860 26911
rect 12808 26868 12860 26877
rect 13544 26868 13596 26920
rect 18420 27004 18472 27056
rect 18604 27004 18656 27056
rect 21732 27004 21784 27056
rect 17224 26936 17276 26988
rect 24584 27072 24636 27124
rect 23112 27047 23164 27056
rect 23112 27013 23121 27047
rect 23121 27013 23155 27047
rect 23155 27013 23164 27047
rect 23112 27004 23164 27013
rect 23388 27004 23440 27056
rect 25044 27004 25096 27056
rect 19340 26868 19392 26920
rect 19800 26868 19852 26920
rect 21180 26868 21232 26920
rect 22008 26868 22060 26920
rect 8300 26843 8352 26852
rect 8300 26809 8309 26843
rect 8309 26809 8343 26843
rect 8343 26809 8352 26843
rect 8300 26800 8352 26809
rect 9680 26800 9732 26852
rect 10232 26800 10284 26852
rect 17408 26800 17460 26852
rect 20536 26800 20588 26852
rect 23112 26868 23164 26920
rect 23204 26868 23256 26920
rect 3884 26732 3936 26784
rect 10508 26732 10560 26784
rect 11336 26732 11388 26784
rect 14372 26732 14424 26784
rect 17224 26775 17276 26784
rect 17224 26741 17233 26775
rect 17233 26741 17267 26775
rect 17267 26741 17276 26775
rect 17224 26732 17276 26741
rect 19524 26775 19576 26784
rect 19524 26741 19533 26775
rect 19533 26741 19567 26775
rect 19567 26741 19576 26775
rect 19524 26732 19576 26741
rect 23848 26732 23900 26784
rect 24584 26775 24636 26784
rect 24584 26741 24593 26775
rect 24593 26741 24627 26775
rect 24627 26741 24636 26775
rect 24584 26732 24636 26741
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 4068 26571 4120 26580
rect 4068 26537 4077 26571
rect 4077 26537 4111 26571
rect 4111 26537 4120 26571
rect 4068 26528 4120 26537
rect 8576 26528 8628 26580
rect 13636 26528 13688 26580
rect 16672 26528 16724 26580
rect 17776 26528 17828 26580
rect 22192 26528 22244 26580
rect 22652 26528 22704 26580
rect 24584 26528 24636 26580
rect 16764 26460 16816 26512
rect 18420 26460 18472 26512
rect 19708 26460 19760 26512
rect 6460 26435 6512 26444
rect 6460 26401 6469 26435
rect 6469 26401 6503 26435
rect 6503 26401 6512 26435
rect 6460 26392 6512 26401
rect 8300 26392 8352 26444
rect 9128 26435 9180 26444
rect 9128 26401 9137 26435
rect 9137 26401 9171 26435
rect 9171 26401 9180 26435
rect 9128 26392 9180 26401
rect 11704 26392 11756 26444
rect 11796 26392 11848 26444
rect 17592 26392 17644 26444
rect 18972 26392 19024 26444
rect 20260 26392 20312 26444
rect 22008 26460 22060 26512
rect 22560 26460 22612 26512
rect 23388 26460 23440 26512
rect 24952 26460 25004 26512
rect 22468 26392 22520 26444
rect 24584 26392 24636 26444
rect 2044 26324 2096 26376
rect 9956 26367 10008 26376
rect 9956 26333 9965 26367
rect 9965 26333 9999 26367
rect 9999 26333 10008 26367
rect 9956 26324 10008 26333
rect 11336 26324 11388 26376
rect 14280 26324 14332 26376
rect 15384 26367 15436 26376
rect 15384 26333 15393 26367
rect 15393 26333 15427 26367
rect 15427 26333 15436 26367
rect 15384 26324 15436 26333
rect 2780 26299 2832 26308
rect 2780 26265 2789 26299
rect 2789 26265 2823 26299
rect 2823 26265 2832 26299
rect 2780 26256 2832 26265
rect 8944 26256 8996 26308
rect 7104 26188 7156 26240
rect 7656 26188 7708 26240
rect 13728 26256 13780 26308
rect 12532 26231 12584 26240
rect 12532 26197 12541 26231
rect 12541 26197 12575 26231
rect 12575 26197 12584 26231
rect 12532 26188 12584 26197
rect 14556 26188 14608 26240
rect 17224 26188 17276 26240
rect 20628 26256 20680 26308
rect 21180 26256 21232 26308
rect 22284 26324 22336 26376
rect 24400 26324 24452 26376
rect 20996 26188 21048 26240
rect 23388 26256 23440 26308
rect 25044 26256 25096 26308
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 1768 25984 1820 26036
rect 7104 25984 7156 26036
rect 8852 25984 8904 26036
rect 3516 25916 3568 25968
rect 4068 25916 4120 25968
rect 10508 25984 10560 26036
rect 10876 26027 10928 26036
rect 10876 25993 10885 26027
rect 10885 25993 10919 26027
rect 10919 25993 10928 26027
rect 10876 25984 10928 25993
rect 2872 25848 2924 25900
rect 12532 25916 12584 25968
rect 2780 25780 2832 25832
rect 3608 25780 3660 25832
rect 4804 25848 4856 25900
rect 8484 25848 8536 25900
rect 6184 25780 6236 25832
rect 7840 25780 7892 25832
rect 9404 25848 9456 25900
rect 15384 25984 15436 26036
rect 15568 25984 15620 26036
rect 19340 26027 19392 26036
rect 19340 25993 19349 26027
rect 19349 25993 19383 26027
rect 19383 25993 19392 26027
rect 19340 25984 19392 25993
rect 19524 25984 19576 26036
rect 20352 26027 20404 26036
rect 20352 25993 20361 26027
rect 20361 25993 20395 26027
rect 20395 25993 20404 26027
rect 20352 25984 20404 25993
rect 22376 26027 22428 26036
rect 22376 25993 22385 26027
rect 22385 25993 22419 26027
rect 22419 25993 22428 26027
rect 22376 25984 22428 25993
rect 22744 25984 22796 26036
rect 14556 25916 14608 25968
rect 17500 25848 17552 25900
rect 20076 25916 20128 25968
rect 3424 25755 3476 25764
rect 3424 25721 3433 25755
rect 3433 25721 3467 25755
rect 3467 25721 3476 25755
rect 3424 25712 3476 25721
rect 8576 25712 8628 25764
rect 9864 25780 9916 25832
rect 11796 25780 11848 25832
rect 12348 25780 12400 25832
rect 12532 25780 12584 25832
rect 14372 25780 14424 25832
rect 12256 25712 12308 25764
rect 4252 25687 4304 25696
rect 4252 25653 4261 25687
rect 4261 25653 4295 25687
rect 4295 25653 4304 25687
rect 4252 25644 4304 25653
rect 11428 25644 11480 25696
rect 14924 25780 14976 25832
rect 16028 25823 16080 25832
rect 16028 25789 16037 25823
rect 16037 25789 16071 25823
rect 16071 25789 16080 25823
rect 16028 25780 16080 25789
rect 17868 25823 17920 25832
rect 17868 25789 17877 25823
rect 17877 25789 17911 25823
rect 17911 25789 17920 25823
rect 17868 25780 17920 25789
rect 18236 25780 18288 25832
rect 14556 25712 14608 25764
rect 17224 25712 17276 25764
rect 22192 25848 22244 25900
rect 23848 25848 23900 25900
rect 21640 25780 21692 25832
rect 22744 25780 22796 25832
rect 25136 25823 25188 25832
rect 25136 25789 25145 25823
rect 25145 25789 25179 25823
rect 25179 25789 25188 25823
rect 25136 25780 25188 25789
rect 23756 25712 23808 25764
rect 14924 25644 14976 25696
rect 18880 25644 18932 25696
rect 20996 25687 21048 25696
rect 20996 25653 21005 25687
rect 21005 25653 21039 25687
rect 21039 25653 21048 25687
rect 20996 25644 21048 25653
rect 21180 25644 21232 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 7472 25440 7524 25492
rect 7656 25440 7708 25492
rect 8852 25440 8904 25492
rect 13544 25440 13596 25492
rect 16764 25440 16816 25492
rect 12256 25372 12308 25424
rect 7656 25304 7708 25356
rect 8576 25347 8628 25356
rect 8576 25313 8585 25347
rect 8585 25313 8619 25347
rect 8619 25313 8628 25347
rect 8576 25304 8628 25313
rect 9404 25347 9456 25356
rect 9404 25313 9413 25347
rect 9413 25313 9447 25347
rect 9447 25313 9456 25347
rect 9404 25304 9456 25313
rect 9680 25304 9732 25356
rect 11428 25304 11480 25356
rect 12808 25304 12860 25356
rect 15384 25304 15436 25356
rect 16672 25304 16724 25356
rect 4068 25279 4120 25288
rect 4068 25245 4086 25279
rect 4086 25245 4120 25279
rect 4068 25236 4120 25245
rect 10784 25236 10836 25288
rect 11796 25279 11848 25288
rect 11796 25245 11805 25279
rect 11805 25245 11839 25279
rect 11839 25245 11848 25279
rect 11796 25236 11848 25245
rect 17224 25236 17276 25288
rect 18236 25440 18288 25492
rect 22836 25440 22888 25492
rect 24952 25440 25004 25492
rect 25504 25483 25556 25492
rect 25504 25449 25513 25483
rect 25513 25449 25547 25483
rect 25547 25449 25556 25483
rect 25504 25440 25556 25449
rect 24860 25372 24912 25424
rect 19064 25304 19116 25356
rect 20076 25347 20128 25356
rect 20076 25313 20085 25347
rect 20085 25313 20119 25347
rect 20119 25313 20128 25347
rect 20076 25304 20128 25313
rect 21088 25304 21140 25356
rect 22652 25347 22704 25356
rect 22652 25313 22661 25347
rect 22661 25313 22695 25347
rect 22695 25313 22704 25347
rect 22652 25304 22704 25313
rect 24032 25304 24084 25356
rect 18328 25236 18380 25288
rect 19432 25236 19484 25288
rect 21640 25236 21692 25288
rect 23940 25236 23992 25288
rect 7104 25168 7156 25220
rect 8392 25168 8444 25220
rect 12532 25168 12584 25220
rect 22376 25168 22428 25220
rect 3976 25100 4028 25152
rect 5540 25100 5592 25152
rect 11980 25100 12032 25152
rect 12624 25143 12676 25152
rect 12624 25109 12633 25143
rect 12633 25109 12667 25143
rect 12667 25109 12676 25143
rect 12624 25100 12676 25109
rect 12808 25100 12860 25152
rect 15108 25143 15160 25152
rect 15108 25109 15117 25143
rect 15117 25109 15151 25143
rect 15151 25109 15160 25143
rect 15108 25100 15160 25109
rect 16856 25100 16908 25152
rect 17040 25100 17092 25152
rect 17868 25100 17920 25152
rect 19524 25100 19576 25152
rect 22468 25100 22520 25152
rect 24032 25211 24084 25220
rect 24032 25177 24041 25211
rect 24041 25177 24075 25211
rect 24075 25177 24084 25211
rect 24032 25168 24084 25177
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 4252 24896 4304 24948
rect 7840 24896 7892 24948
rect 12624 24896 12676 24948
rect 16856 24939 16908 24948
rect 16856 24905 16865 24939
rect 16865 24905 16899 24939
rect 16899 24905 16908 24939
rect 16856 24896 16908 24905
rect 7104 24828 7156 24880
rect 7472 24828 7524 24880
rect 4988 24760 5040 24812
rect 7380 24803 7432 24812
rect 7380 24769 7389 24803
rect 7389 24769 7423 24803
rect 7423 24769 7432 24803
rect 7380 24760 7432 24769
rect 7748 24760 7800 24812
rect 13360 24828 13412 24880
rect 6000 24692 6052 24744
rect 8116 24735 8168 24744
rect 8116 24701 8125 24735
rect 8125 24701 8159 24735
rect 8159 24701 8168 24735
rect 8116 24692 8168 24701
rect 9312 24735 9364 24744
rect 9312 24701 9321 24735
rect 9321 24701 9355 24735
rect 9355 24701 9364 24735
rect 9312 24692 9364 24701
rect 9680 24692 9732 24744
rect 13636 24760 13688 24812
rect 13820 24803 13872 24812
rect 13820 24769 13829 24803
rect 13829 24769 13863 24803
rect 13863 24769 13872 24803
rect 13820 24760 13872 24769
rect 15016 24760 15068 24812
rect 16856 24760 16908 24812
rect 17776 24896 17828 24948
rect 18328 24896 18380 24948
rect 19340 24896 19392 24948
rect 19616 24896 19668 24948
rect 18420 24760 18472 24812
rect 22652 24828 22704 24880
rect 8392 24624 8444 24676
rect 3976 24556 4028 24608
rect 7472 24556 7524 24608
rect 12532 24624 12584 24676
rect 14096 24735 14148 24744
rect 14096 24701 14105 24735
rect 14105 24701 14139 24735
rect 14139 24701 14148 24735
rect 14096 24692 14148 24701
rect 14372 24692 14424 24744
rect 16580 24692 16632 24744
rect 17500 24735 17552 24744
rect 17500 24701 17509 24735
rect 17509 24701 17543 24735
rect 17543 24701 17552 24735
rect 17500 24692 17552 24701
rect 18604 24735 18656 24744
rect 18604 24701 18613 24735
rect 18613 24701 18647 24735
rect 18647 24701 18656 24735
rect 18604 24692 18656 24701
rect 18696 24692 18748 24744
rect 20720 24735 20772 24744
rect 20720 24701 20729 24735
rect 20729 24701 20763 24735
rect 20763 24701 20772 24735
rect 20720 24692 20772 24701
rect 22008 24760 22060 24812
rect 22100 24760 22152 24812
rect 24308 24760 24360 24812
rect 24952 24828 25004 24880
rect 25504 24760 25556 24812
rect 15108 24624 15160 24676
rect 11152 24556 11204 24608
rect 12440 24556 12492 24608
rect 12624 24556 12676 24608
rect 13360 24556 13412 24608
rect 17684 24624 17736 24676
rect 20168 24624 20220 24676
rect 20628 24624 20680 24676
rect 18512 24556 18564 24608
rect 22652 24624 22704 24676
rect 24676 24735 24728 24744
rect 24676 24701 24685 24735
rect 24685 24701 24719 24735
rect 24719 24701 24728 24735
rect 24676 24692 24728 24701
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 3332 24352 3384 24404
rect 4436 24352 4488 24404
rect 6184 24395 6236 24404
rect 6184 24361 6193 24395
rect 6193 24361 6227 24395
rect 6227 24361 6236 24395
rect 6184 24352 6236 24361
rect 8668 24352 8720 24404
rect 9312 24352 9364 24404
rect 6092 24284 6144 24336
rect 4252 24259 4304 24268
rect 4252 24225 4261 24259
rect 4261 24225 4295 24259
rect 4295 24225 4304 24259
rect 4252 24216 4304 24225
rect 4988 24216 5040 24268
rect 8300 24216 8352 24268
rect 13636 24352 13688 24404
rect 15476 24352 15528 24404
rect 16856 24352 16908 24404
rect 10048 24259 10100 24268
rect 10048 24225 10057 24259
rect 10057 24225 10091 24259
rect 10091 24225 10100 24259
rect 10048 24216 10100 24225
rect 2780 24148 2832 24200
rect 3516 24148 3568 24200
rect 3976 24191 4028 24200
rect 3976 24157 3985 24191
rect 3985 24157 4019 24191
rect 4019 24157 4028 24191
rect 3976 24148 4028 24157
rect 7012 24148 7064 24200
rect 8576 24148 8628 24200
rect 11244 24259 11296 24268
rect 11244 24225 11253 24259
rect 11253 24225 11287 24259
rect 11287 24225 11296 24259
rect 11244 24216 11296 24225
rect 24676 24284 24728 24336
rect 11152 24191 11204 24200
rect 11152 24157 11161 24191
rect 11161 24157 11195 24191
rect 11195 24157 11204 24191
rect 11152 24148 11204 24157
rect 12808 24216 12860 24268
rect 13820 24216 13872 24268
rect 16948 24216 17000 24268
rect 17040 24259 17092 24268
rect 17040 24225 17049 24259
rect 17049 24225 17083 24259
rect 17083 24225 17092 24259
rect 17040 24216 17092 24225
rect 22100 24216 22152 24268
rect 24952 24216 25004 24268
rect 4528 24080 4580 24132
rect 4988 24080 5040 24132
rect 10968 24080 11020 24132
rect 16764 24191 16816 24200
rect 16764 24157 16773 24191
rect 16773 24157 16807 24191
rect 16807 24157 16816 24191
rect 16764 24148 16816 24157
rect 17316 24148 17368 24200
rect 20996 24148 21048 24200
rect 21456 24148 21508 24200
rect 21548 24148 21600 24200
rect 11520 24080 11572 24132
rect 12164 24080 12216 24132
rect 14096 24080 14148 24132
rect 17500 24080 17552 24132
rect 18420 24080 18472 24132
rect 18604 24080 18656 24132
rect 19892 24080 19944 24132
rect 21824 24080 21876 24132
rect 22192 24123 22244 24132
rect 22192 24089 22201 24123
rect 22201 24089 22235 24123
rect 22235 24089 22244 24123
rect 22192 24080 22244 24089
rect 23480 24148 23532 24200
rect 1860 24012 1912 24064
rect 8760 24012 8812 24064
rect 9772 24055 9824 24064
rect 9772 24021 9781 24055
rect 9781 24021 9815 24055
rect 9815 24021 9824 24055
rect 9772 24012 9824 24021
rect 10508 24055 10560 24064
rect 10508 24021 10517 24055
rect 10517 24021 10551 24055
rect 10551 24021 10560 24055
rect 10508 24012 10560 24021
rect 11152 24012 11204 24064
rect 11980 24055 12032 24064
rect 11980 24021 11989 24055
rect 11989 24021 12023 24055
rect 12023 24021 12032 24055
rect 11980 24012 12032 24021
rect 13636 24012 13688 24064
rect 16672 24012 16724 24064
rect 17868 24012 17920 24064
rect 20260 24012 20312 24064
rect 22468 24012 22520 24064
rect 24860 24012 24912 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 6000 23851 6052 23860
rect 6000 23817 6009 23851
rect 6009 23817 6043 23851
rect 6043 23817 6052 23851
rect 6000 23808 6052 23817
rect 6828 23808 6880 23860
rect 9680 23808 9732 23860
rect 9772 23808 9824 23860
rect 10508 23808 10560 23860
rect 11244 23808 11296 23860
rect 11520 23808 11572 23860
rect 12440 23808 12492 23860
rect 12808 23808 12860 23860
rect 17500 23808 17552 23860
rect 7104 23740 7156 23792
rect 8208 23740 8260 23792
rect 11888 23740 11940 23792
rect 13912 23783 13964 23792
rect 13912 23749 13921 23783
rect 13921 23749 13955 23783
rect 13955 23749 13964 23783
rect 13912 23740 13964 23749
rect 17960 23740 18012 23792
rect 1768 23715 1820 23724
rect 1768 23681 1777 23715
rect 1777 23681 1811 23715
rect 1811 23681 1820 23715
rect 1768 23672 1820 23681
rect 20720 23808 20772 23860
rect 20628 23740 20680 23792
rect 23480 23740 23532 23792
rect 1308 23604 1360 23656
rect 3976 23604 4028 23656
rect 7564 23604 7616 23656
rect 7656 23647 7708 23656
rect 7656 23613 7665 23647
rect 7665 23613 7699 23647
rect 7699 23613 7708 23647
rect 7656 23604 7708 23613
rect 8576 23604 8628 23656
rect 11704 23604 11756 23656
rect 12072 23604 12124 23656
rect 14740 23604 14792 23656
rect 17040 23647 17092 23656
rect 17040 23613 17049 23647
rect 17049 23613 17083 23647
rect 17083 23613 17092 23647
rect 17040 23604 17092 23613
rect 18604 23604 18656 23656
rect 19800 23604 19852 23656
rect 22008 23672 22060 23724
rect 22100 23672 22152 23724
rect 24308 23672 24360 23724
rect 25320 23715 25372 23724
rect 25320 23681 25329 23715
rect 25329 23681 25363 23715
rect 25363 23681 25372 23715
rect 25320 23672 25372 23681
rect 5724 23468 5776 23520
rect 9956 23536 10008 23588
rect 11612 23579 11664 23588
rect 11612 23545 11621 23579
rect 11621 23545 11655 23579
rect 11655 23545 11664 23579
rect 11612 23536 11664 23545
rect 16488 23536 16540 23588
rect 11336 23468 11388 23520
rect 12072 23468 12124 23520
rect 12440 23511 12492 23520
rect 12440 23477 12449 23511
rect 12449 23477 12483 23511
rect 12483 23477 12492 23511
rect 12440 23468 12492 23477
rect 13360 23468 13412 23520
rect 20168 23468 20220 23520
rect 23572 23604 23624 23656
rect 24584 23604 24636 23656
rect 21456 23468 21508 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 2044 23307 2096 23316
rect 2044 23273 2053 23307
rect 2053 23273 2087 23307
rect 2087 23273 2096 23307
rect 2044 23264 2096 23273
rect 2872 23264 2924 23316
rect 7564 23307 7616 23316
rect 7564 23273 7573 23307
rect 7573 23273 7607 23307
rect 7607 23273 7616 23307
rect 7564 23264 7616 23273
rect 10876 23264 10928 23316
rect 12624 23264 12676 23316
rect 14556 23264 14608 23316
rect 16028 23307 16080 23316
rect 16028 23273 16037 23307
rect 16037 23273 16071 23307
rect 16071 23273 16080 23307
rect 16028 23264 16080 23273
rect 19432 23264 19484 23316
rect 20076 23264 20128 23316
rect 20444 23264 20496 23316
rect 9680 23196 9732 23248
rect 12440 23196 12492 23248
rect 23664 23196 23716 23248
rect 24584 23196 24636 23248
rect 2872 23128 2924 23180
rect 3332 23128 3384 23180
rect 5724 23128 5776 23180
rect 6460 23128 6512 23180
rect 7104 23128 7156 23180
rect 3792 22992 3844 23044
rect 3976 23060 4028 23112
rect 4344 23060 4396 23112
rect 11888 23171 11940 23180
rect 11888 23137 11897 23171
rect 11897 23137 11931 23171
rect 11931 23137 11940 23171
rect 11888 23128 11940 23137
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 14280 23171 14332 23180
rect 14280 23137 14289 23171
rect 14289 23137 14323 23171
rect 14323 23137 14332 23171
rect 14280 23128 14332 23137
rect 15292 23128 15344 23180
rect 18604 23128 18656 23180
rect 7656 23060 7708 23112
rect 9312 23060 9364 23112
rect 11612 23060 11664 23112
rect 11704 23103 11756 23112
rect 11704 23069 11713 23103
rect 11713 23069 11747 23103
rect 11747 23069 11756 23103
rect 11704 23060 11756 23069
rect 13912 23060 13964 23112
rect 16396 23060 16448 23112
rect 23296 23060 23348 23112
rect 23848 23103 23900 23112
rect 23848 23069 23857 23103
rect 23857 23069 23891 23103
rect 23891 23069 23900 23103
rect 23848 23060 23900 23069
rect 5080 22992 5132 23044
rect 7748 22992 7800 23044
rect 9956 22924 10008 22976
rect 10784 22992 10836 23044
rect 12072 22924 12124 22976
rect 15936 22992 15988 23044
rect 15844 22924 15896 22976
rect 16396 22924 16448 22976
rect 19432 22992 19484 23044
rect 19984 22992 20036 23044
rect 22652 22992 22704 23044
rect 21456 22967 21508 22976
rect 21456 22933 21465 22967
rect 21465 22933 21499 22967
rect 21499 22933 21508 22967
rect 21456 22924 21508 22933
rect 23480 22924 23532 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 1768 22720 1820 22772
rect 8760 22720 8812 22772
rect 9312 22763 9364 22772
rect 9312 22729 9321 22763
rect 9321 22729 9355 22763
rect 9355 22729 9364 22763
rect 9312 22720 9364 22729
rect 9864 22720 9916 22772
rect 10876 22763 10928 22772
rect 10876 22729 10885 22763
rect 10885 22729 10919 22763
rect 10919 22729 10928 22763
rect 10876 22720 10928 22729
rect 12532 22720 12584 22772
rect 14924 22720 14976 22772
rect 16396 22720 16448 22772
rect 16580 22720 16632 22772
rect 17500 22763 17552 22772
rect 17500 22729 17509 22763
rect 17509 22729 17543 22763
rect 17543 22729 17552 22763
rect 17500 22720 17552 22729
rect 11612 22652 11664 22704
rect 12164 22652 12216 22704
rect 2872 22584 2924 22636
rect 6920 22584 6972 22636
rect 15660 22652 15712 22704
rect 20352 22720 20404 22772
rect 23572 22720 23624 22772
rect 24308 22763 24360 22772
rect 18604 22695 18656 22704
rect 18604 22661 18613 22695
rect 18613 22661 18647 22695
rect 18647 22661 18656 22695
rect 18604 22652 18656 22661
rect 19708 22695 19760 22704
rect 19708 22661 19717 22695
rect 19717 22661 19751 22695
rect 19751 22661 19760 22695
rect 19708 22652 19760 22661
rect 24308 22729 24317 22763
rect 24317 22729 24351 22763
rect 24351 22729 24360 22763
rect 24308 22720 24360 22729
rect 25320 22720 25372 22772
rect 6000 22516 6052 22568
rect 7288 22559 7340 22568
rect 7288 22525 7297 22559
rect 7297 22525 7331 22559
rect 7331 22525 7340 22559
rect 7288 22516 7340 22525
rect 7564 22516 7616 22568
rect 8852 22559 8904 22568
rect 8852 22525 8861 22559
rect 8861 22525 8895 22559
rect 8895 22525 8904 22559
rect 8852 22516 8904 22525
rect 10968 22559 11020 22568
rect 10968 22525 10977 22559
rect 10977 22525 11011 22559
rect 11011 22525 11020 22559
rect 10968 22516 11020 22525
rect 13820 22584 13872 22636
rect 16580 22584 16632 22636
rect 16856 22584 16908 22636
rect 19616 22627 19668 22636
rect 19616 22593 19625 22627
rect 19625 22593 19659 22627
rect 19659 22593 19668 22627
rect 19616 22584 19668 22593
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 23572 22584 23624 22636
rect 9404 22448 9456 22500
rect 13636 22448 13688 22500
rect 13912 22559 13964 22568
rect 13912 22525 13921 22559
rect 13921 22525 13955 22559
rect 13955 22525 13964 22559
rect 13912 22516 13964 22525
rect 15936 22516 15988 22568
rect 19800 22559 19852 22568
rect 19800 22525 19809 22559
rect 19809 22525 19843 22559
rect 19843 22525 19852 22559
rect 19800 22516 19852 22525
rect 21640 22516 21692 22568
rect 15844 22448 15896 22500
rect 4252 22380 4304 22432
rect 6276 22380 6328 22432
rect 11612 22423 11664 22432
rect 11612 22389 11621 22423
rect 11621 22389 11655 22423
rect 11655 22389 11664 22423
rect 11612 22380 11664 22389
rect 12532 22380 12584 22432
rect 12808 22380 12860 22432
rect 15568 22380 15620 22432
rect 19248 22423 19300 22432
rect 19248 22389 19257 22423
rect 19257 22389 19291 22423
rect 19291 22389 19300 22423
rect 19248 22380 19300 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 16028 22176 16080 22228
rect 16396 22219 16448 22228
rect 16396 22185 16405 22219
rect 16405 22185 16439 22219
rect 16439 22185 16448 22219
rect 16396 22176 16448 22185
rect 10692 22040 10744 22092
rect 12164 22040 12216 22092
rect 14280 22083 14332 22092
rect 14280 22049 14289 22083
rect 14289 22049 14323 22083
rect 14323 22049 14332 22083
rect 14280 22040 14332 22049
rect 16120 22040 16172 22092
rect 18420 22108 18472 22160
rect 10600 21904 10652 21956
rect 13360 21972 13412 22024
rect 17040 21972 17092 22024
rect 18512 22083 18564 22092
rect 18512 22049 18521 22083
rect 18521 22049 18555 22083
rect 18555 22049 18564 22083
rect 18512 22040 18564 22049
rect 20260 22176 20312 22228
rect 21456 22151 21508 22160
rect 21456 22117 21465 22151
rect 21465 22117 21499 22151
rect 21499 22117 21508 22151
rect 21456 22108 21508 22117
rect 22008 22083 22060 22092
rect 22008 22049 22017 22083
rect 22017 22049 22051 22083
rect 22051 22049 22060 22083
rect 22008 22040 22060 22049
rect 22652 22040 22704 22092
rect 22836 22040 22888 22092
rect 19340 21972 19392 22024
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 23572 21972 23624 22024
rect 4528 21836 4580 21888
rect 10692 21836 10744 21888
rect 13360 21836 13412 21888
rect 14188 21904 14240 21956
rect 14556 21947 14608 21956
rect 14556 21913 14565 21947
rect 14565 21913 14599 21947
rect 14599 21913 14608 21947
rect 14556 21904 14608 21913
rect 16028 21904 16080 21956
rect 15936 21836 15988 21888
rect 21456 21904 21508 21956
rect 19616 21836 19668 21888
rect 19892 21836 19944 21888
rect 21732 21836 21784 21888
rect 24216 21836 24268 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 7012 21632 7064 21684
rect 9680 21632 9732 21684
rect 11980 21632 12032 21684
rect 13820 21632 13872 21684
rect 13912 21675 13964 21684
rect 13912 21641 13921 21675
rect 13921 21641 13955 21675
rect 13955 21641 13964 21675
rect 13912 21632 13964 21641
rect 21088 21632 21140 21684
rect 23480 21632 23532 21684
rect 23572 21632 23624 21684
rect 7656 21564 7708 21616
rect 1860 21496 1912 21548
rect 4160 21496 4212 21548
rect 4528 21539 4580 21548
rect 4528 21505 4537 21539
rect 4537 21505 4571 21539
rect 4571 21505 4580 21539
rect 4528 21496 4580 21505
rect 8944 21496 8996 21548
rect 1308 21428 1360 21480
rect 3608 21471 3660 21480
rect 3608 21437 3617 21471
rect 3617 21437 3651 21471
rect 3651 21437 3660 21471
rect 3608 21428 3660 21437
rect 4068 21428 4120 21480
rect 7656 21471 7708 21480
rect 7656 21437 7665 21471
rect 7665 21437 7699 21471
rect 7699 21437 7708 21471
rect 7656 21428 7708 21437
rect 8760 21471 8812 21480
rect 8760 21437 8769 21471
rect 8769 21437 8803 21471
rect 8803 21437 8812 21471
rect 8760 21428 8812 21437
rect 9128 21428 9180 21480
rect 13636 21564 13688 21616
rect 13820 21496 13872 21548
rect 3792 21403 3844 21412
rect 3792 21369 3801 21403
rect 3801 21369 3835 21403
rect 3835 21369 3844 21403
rect 3792 21360 3844 21369
rect 6920 21360 6972 21412
rect 11888 21428 11940 21480
rect 13728 21428 13780 21480
rect 15200 21539 15252 21548
rect 15200 21505 15209 21539
rect 15209 21505 15243 21539
rect 15243 21505 15252 21539
rect 15200 21496 15252 21505
rect 22008 21564 22060 21616
rect 14188 21471 14240 21480
rect 14188 21437 14197 21471
rect 14197 21437 14231 21471
rect 14231 21437 14240 21471
rect 14188 21428 14240 21437
rect 14464 21428 14516 21480
rect 15108 21428 15160 21480
rect 15476 21471 15528 21480
rect 15476 21437 15485 21471
rect 15485 21437 15519 21471
rect 15519 21437 15528 21471
rect 15476 21428 15528 21437
rect 11520 21360 11572 21412
rect 12348 21360 12400 21412
rect 17408 21496 17460 21548
rect 19984 21496 20036 21548
rect 22836 21496 22888 21548
rect 23664 21607 23716 21616
rect 23664 21573 23673 21607
rect 23673 21573 23707 21607
rect 23707 21573 23716 21607
rect 23664 21564 23716 21573
rect 17592 21428 17644 21480
rect 17776 21428 17828 21480
rect 18696 21360 18748 21412
rect 20168 21428 20220 21480
rect 20444 21428 20496 21480
rect 22560 21471 22612 21480
rect 22560 21437 22569 21471
rect 22569 21437 22603 21471
rect 22603 21437 22612 21471
rect 22560 21428 22612 21437
rect 22652 21428 22704 21480
rect 20260 21360 20312 21412
rect 20904 21360 20956 21412
rect 5816 21292 5868 21344
rect 10324 21292 10376 21344
rect 10876 21292 10928 21344
rect 13452 21292 13504 21344
rect 15292 21292 15344 21344
rect 15476 21292 15528 21344
rect 19064 21292 19116 21344
rect 20444 21335 20496 21344
rect 20444 21301 20453 21335
rect 20453 21301 20487 21335
rect 20487 21301 20496 21335
rect 20444 21292 20496 21301
rect 22284 21292 22336 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 2872 21088 2924 21140
rect 7288 21088 7340 21140
rect 12072 21088 12124 21140
rect 14464 21088 14516 21140
rect 16580 21088 16632 21140
rect 15200 21020 15252 21072
rect 19984 21088 20036 21140
rect 21548 21088 21600 21140
rect 19340 21020 19392 21072
rect 21456 21020 21508 21072
rect 22560 21020 22612 21072
rect 7840 20952 7892 21004
rect 10048 20952 10100 21004
rect 11888 20952 11940 21004
rect 4068 20884 4120 20936
rect 4252 20927 4304 20936
rect 4252 20893 4261 20927
rect 4261 20893 4295 20927
rect 4295 20893 4304 20927
rect 4252 20884 4304 20893
rect 1768 20748 1820 20800
rect 2780 20748 2832 20800
rect 5448 20748 5500 20800
rect 8668 20816 8720 20868
rect 11336 20884 11388 20936
rect 9956 20816 10008 20868
rect 10324 20816 10376 20868
rect 14280 20884 14332 20936
rect 17776 20952 17828 21004
rect 15752 20927 15804 20936
rect 15752 20893 15761 20927
rect 15761 20893 15795 20927
rect 15795 20893 15804 20927
rect 15752 20884 15804 20893
rect 17592 20927 17644 20936
rect 17592 20893 17601 20927
rect 17601 20893 17635 20927
rect 17635 20893 17644 20927
rect 17592 20884 17644 20893
rect 17684 20884 17736 20936
rect 14832 20859 14884 20868
rect 10416 20748 10468 20800
rect 10968 20748 11020 20800
rect 14832 20825 14841 20859
rect 14841 20825 14875 20859
rect 14875 20825 14884 20859
rect 14832 20816 14884 20825
rect 15384 20816 15436 20868
rect 16764 20816 16816 20868
rect 19432 20952 19484 21004
rect 20720 20952 20772 21004
rect 24860 20952 24912 21004
rect 21456 20884 21508 20936
rect 22192 20884 22244 20936
rect 20168 20859 20220 20868
rect 20168 20825 20177 20859
rect 20177 20825 20211 20859
rect 20211 20825 20220 20859
rect 20168 20816 20220 20825
rect 13912 20791 13964 20800
rect 13912 20757 13921 20791
rect 13921 20757 13955 20791
rect 13955 20757 13964 20791
rect 13912 20748 13964 20757
rect 14372 20791 14424 20800
rect 14372 20757 14381 20791
rect 14381 20757 14415 20791
rect 14415 20757 14424 20791
rect 14372 20748 14424 20757
rect 15476 20748 15528 20800
rect 16580 20748 16632 20800
rect 24860 20816 24912 20868
rect 21640 20791 21692 20800
rect 21640 20757 21649 20791
rect 21649 20757 21683 20791
rect 21683 20757 21692 20791
rect 21640 20748 21692 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 6552 20544 6604 20596
rect 8852 20544 8904 20596
rect 8944 20544 8996 20596
rect 4344 20476 4396 20528
rect 7104 20476 7156 20528
rect 6552 20451 6604 20460
rect 6552 20417 6561 20451
rect 6561 20417 6595 20451
rect 6595 20417 6604 20451
rect 6552 20408 6604 20417
rect 5724 20340 5776 20392
rect 8944 20408 8996 20460
rect 11980 20544 12032 20596
rect 13636 20544 13688 20596
rect 14004 20544 14056 20596
rect 17316 20587 17368 20596
rect 17316 20553 17325 20587
rect 17325 20553 17359 20587
rect 17359 20553 17368 20587
rect 17316 20544 17368 20553
rect 10968 20476 11020 20528
rect 12256 20476 12308 20528
rect 19340 20587 19392 20596
rect 19340 20553 19349 20587
rect 19349 20553 19383 20587
rect 19383 20553 19392 20587
rect 19340 20544 19392 20553
rect 19524 20544 19576 20596
rect 11704 20408 11756 20460
rect 23388 20476 23440 20528
rect 19156 20408 19208 20460
rect 22376 20408 22428 20460
rect 25044 20408 25096 20460
rect 8760 20315 8812 20324
rect 8760 20281 8769 20315
rect 8769 20281 8803 20315
rect 8803 20281 8812 20315
rect 8760 20272 8812 20281
rect 9588 20340 9640 20392
rect 11152 20340 11204 20392
rect 11612 20272 11664 20324
rect 12716 20383 12768 20392
rect 12716 20349 12725 20383
rect 12725 20349 12759 20383
rect 12759 20349 12768 20383
rect 12716 20340 12768 20349
rect 21640 20340 21692 20392
rect 23296 20340 23348 20392
rect 17040 20272 17092 20324
rect 5816 20204 5868 20256
rect 8300 20247 8352 20256
rect 8300 20213 8309 20247
rect 8309 20213 8343 20247
rect 8343 20213 8352 20247
rect 8300 20204 8352 20213
rect 9128 20204 9180 20256
rect 9588 20204 9640 20256
rect 12072 20247 12124 20256
rect 12072 20213 12081 20247
rect 12081 20213 12115 20247
rect 12115 20213 12124 20247
rect 12072 20204 12124 20213
rect 13636 20204 13688 20256
rect 15108 20204 15160 20256
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 16856 20204 16908 20256
rect 18420 20204 18472 20256
rect 19800 20204 19852 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 5080 20043 5132 20052
rect 5080 20009 5089 20043
rect 5089 20009 5123 20043
rect 5123 20009 5132 20043
rect 5080 20000 5132 20009
rect 5724 20000 5776 20052
rect 6552 20000 6604 20052
rect 11704 20043 11756 20052
rect 11704 20009 11713 20043
rect 11713 20009 11747 20043
rect 11747 20009 11756 20043
rect 11704 20000 11756 20009
rect 11980 20000 12032 20052
rect 12256 20000 12308 20052
rect 13820 20000 13872 20052
rect 20812 20000 20864 20052
rect 12164 19932 12216 19984
rect 12624 19932 12676 19984
rect 8300 19864 8352 19916
rect 8852 19864 8904 19916
rect 12256 19907 12308 19916
rect 12256 19873 12265 19907
rect 12265 19873 12299 19907
rect 12299 19873 12308 19907
rect 12256 19864 12308 19873
rect 14188 19864 14240 19916
rect 7104 19796 7156 19848
rect 7748 19839 7800 19848
rect 7748 19805 7757 19839
rect 7757 19805 7791 19839
rect 7791 19805 7800 19839
rect 7748 19796 7800 19805
rect 8208 19796 8260 19848
rect 9036 19796 9088 19848
rect 12440 19796 12492 19848
rect 18788 19932 18840 19984
rect 20260 19932 20312 19984
rect 17868 19864 17920 19916
rect 17776 19839 17828 19848
rect 17776 19805 17785 19839
rect 17785 19805 17819 19839
rect 17819 19805 17828 19839
rect 17776 19796 17828 19805
rect 18880 19796 18932 19848
rect 24952 19864 25004 19916
rect 25228 19796 25280 19848
rect 7288 19660 7340 19712
rect 7656 19728 7708 19780
rect 8852 19660 8904 19712
rect 9036 19660 9088 19712
rect 11428 19728 11480 19780
rect 17316 19771 17368 19780
rect 17316 19737 17325 19771
rect 17325 19737 17359 19771
rect 17359 19737 17368 19771
rect 17316 19728 17368 19737
rect 18788 19728 18840 19780
rect 23848 19728 23900 19780
rect 13728 19660 13780 19712
rect 18512 19703 18564 19712
rect 18512 19669 18521 19703
rect 18521 19669 18555 19703
rect 18555 19669 18564 19703
rect 18512 19660 18564 19669
rect 19340 19703 19392 19712
rect 19340 19669 19349 19703
rect 19349 19669 19383 19703
rect 19383 19669 19392 19703
rect 19340 19660 19392 19669
rect 19432 19660 19484 19712
rect 21548 19660 21600 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 1492 19456 1544 19508
rect 4160 19456 4212 19508
rect 7840 19456 7892 19508
rect 9404 19456 9456 19508
rect 11612 19456 11664 19508
rect 7104 19388 7156 19440
rect 17224 19456 17276 19508
rect 17316 19456 17368 19508
rect 19432 19499 19484 19508
rect 19432 19465 19441 19499
rect 19441 19465 19475 19499
rect 19475 19465 19484 19499
rect 19432 19456 19484 19465
rect 19524 19456 19576 19508
rect 20812 19456 20864 19508
rect 21180 19499 21232 19508
rect 21180 19465 21189 19499
rect 21189 19465 21223 19499
rect 21223 19465 21232 19499
rect 21180 19456 21232 19465
rect 21824 19456 21876 19508
rect 14924 19388 14976 19440
rect 19248 19388 19300 19440
rect 3608 19320 3660 19372
rect 6276 19320 6328 19372
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 8392 19320 8444 19372
rect 8576 19320 8628 19372
rect 13360 19320 13412 19372
rect 13544 19320 13596 19372
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 9220 19252 9272 19304
rect 11060 19252 11112 19304
rect 12992 19252 13044 19304
rect 14096 19320 14148 19372
rect 14740 19320 14792 19372
rect 17040 19363 17092 19372
rect 17040 19329 17049 19363
rect 17049 19329 17083 19363
rect 17083 19329 17092 19363
rect 17040 19320 17092 19329
rect 20536 19388 20588 19440
rect 22560 19388 22612 19440
rect 14188 19295 14240 19304
rect 7564 19116 7616 19168
rect 10876 19159 10928 19168
rect 10876 19125 10885 19159
rect 10885 19125 10919 19159
rect 10919 19125 10928 19159
rect 10876 19116 10928 19125
rect 11060 19159 11112 19168
rect 11060 19125 11069 19159
rect 11069 19125 11103 19159
rect 11103 19125 11112 19159
rect 11060 19116 11112 19125
rect 11152 19116 11204 19168
rect 11336 19116 11388 19168
rect 11704 19116 11756 19168
rect 13084 19184 13136 19236
rect 13268 19184 13320 19236
rect 12440 19116 12492 19168
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 14556 19295 14608 19304
rect 14556 19261 14565 19295
rect 14565 19261 14599 19295
rect 14599 19261 14608 19295
rect 14556 19252 14608 19261
rect 14004 19184 14056 19236
rect 19340 19252 19392 19304
rect 19248 19184 19300 19236
rect 21272 19252 21324 19304
rect 21824 19252 21876 19304
rect 22008 19295 22060 19304
rect 22008 19261 22017 19295
rect 22017 19261 22051 19295
rect 22051 19261 22060 19295
rect 22008 19252 22060 19261
rect 22744 19252 22796 19304
rect 17132 19116 17184 19168
rect 17776 19116 17828 19168
rect 18880 19159 18932 19168
rect 18880 19125 18889 19159
rect 18889 19125 18923 19159
rect 18923 19125 18932 19159
rect 18880 19116 18932 19125
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 22652 19116 22704 19168
rect 24400 19116 24452 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 8300 18912 8352 18964
rect 11152 18912 11204 18964
rect 12164 18955 12216 18964
rect 12164 18921 12173 18955
rect 12173 18921 12207 18955
rect 12207 18921 12216 18955
rect 12164 18912 12216 18921
rect 13728 18912 13780 18964
rect 1308 18776 1360 18828
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 6552 18708 6604 18760
rect 9312 18708 9364 18760
rect 12716 18844 12768 18896
rect 13452 18819 13504 18828
rect 13452 18785 13461 18819
rect 13461 18785 13495 18819
rect 13495 18785 13504 18819
rect 13452 18776 13504 18785
rect 13820 18844 13872 18896
rect 14004 18844 14056 18896
rect 14188 18776 14240 18828
rect 14556 18776 14608 18828
rect 14832 18819 14884 18828
rect 14832 18785 14841 18819
rect 14841 18785 14875 18819
rect 14875 18785 14884 18819
rect 14832 18776 14884 18785
rect 8576 18615 8628 18624
rect 8576 18581 8585 18615
rect 8585 18581 8619 18615
rect 8619 18581 8628 18615
rect 8576 18572 8628 18581
rect 9128 18572 9180 18624
rect 12256 18640 12308 18692
rect 17776 18912 17828 18964
rect 18972 18955 19024 18964
rect 18972 18921 18981 18955
rect 18981 18921 19015 18955
rect 19015 18921 19024 18955
rect 18972 18912 19024 18921
rect 22744 18912 22796 18964
rect 24400 18955 24452 18964
rect 24400 18921 24409 18955
rect 24409 18921 24443 18955
rect 24443 18921 24452 18955
rect 24400 18912 24452 18921
rect 18512 18844 18564 18896
rect 15844 18776 15896 18828
rect 16212 18751 16264 18760
rect 16212 18717 16221 18751
rect 16221 18717 16255 18751
rect 16255 18717 16264 18751
rect 16212 18708 16264 18717
rect 20628 18844 20680 18896
rect 18972 18708 19024 18760
rect 20444 18708 20496 18760
rect 12808 18640 12860 18692
rect 13728 18640 13780 18692
rect 11060 18572 11112 18624
rect 11796 18572 11848 18624
rect 11980 18572 12032 18624
rect 13360 18615 13412 18624
rect 13360 18581 13369 18615
rect 13369 18581 13403 18615
rect 13403 18581 13412 18615
rect 13360 18572 13412 18581
rect 21732 18640 21784 18692
rect 22008 18640 22060 18692
rect 22560 18683 22612 18692
rect 22560 18649 22569 18683
rect 22569 18649 22603 18683
rect 22603 18649 22612 18683
rect 22560 18640 22612 18649
rect 22652 18640 22704 18692
rect 18972 18572 19024 18624
rect 19708 18615 19760 18624
rect 19708 18581 19717 18615
rect 19717 18581 19751 18615
rect 19751 18581 19760 18615
rect 19708 18572 19760 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 7472 18368 7524 18420
rect 10416 18411 10468 18420
rect 10416 18377 10425 18411
rect 10425 18377 10459 18411
rect 10459 18377 10468 18411
rect 10416 18368 10468 18377
rect 12164 18368 12216 18420
rect 13360 18368 13412 18420
rect 18328 18368 18380 18420
rect 9312 18343 9364 18352
rect 9312 18309 9321 18343
rect 9321 18309 9355 18343
rect 9355 18309 9364 18343
rect 9312 18300 9364 18309
rect 11704 18300 11756 18352
rect 13728 18300 13780 18352
rect 16304 18300 16356 18352
rect 16488 18300 16540 18352
rect 17500 18343 17552 18352
rect 17500 18309 17509 18343
rect 17509 18309 17543 18343
rect 17543 18309 17552 18343
rect 17500 18300 17552 18309
rect 19340 18368 19392 18420
rect 20628 18300 20680 18352
rect 4896 18096 4948 18148
rect 9772 18232 9824 18284
rect 10324 18232 10376 18284
rect 11888 18232 11940 18284
rect 7564 18164 7616 18216
rect 4160 18028 4212 18080
rect 5540 18028 5592 18080
rect 8668 18028 8720 18080
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 9864 18028 9916 18080
rect 11060 18207 11112 18216
rect 11060 18173 11069 18207
rect 11069 18173 11103 18207
rect 11103 18173 11112 18207
rect 11060 18164 11112 18173
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 12440 18164 12492 18216
rect 11520 18096 11572 18148
rect 12348 18096 12400 18148
rect 15016 18232 15068 18284
rect 12624 18028 12676 18080
rect 13268 18028 13320 18080
rect 15292 18164 15344 18216
rect 15936 18164 15988 18216
rect 16212 18164 16264 18216
rect 16488 18164 16540 18216
rect 19156 18164 19208 18216
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 24032 18275 24084 18284
rect 24032 18241 24041 18275
rect 24041 18241 24075 18275
rect 24075 18241 24084 18275
rect 24032 18232 24084 18241
rect 23388 18164 23440 18216
rect 24768 18207 24820 18216
rect 24768 18173 24777 18207
rect 24777 18173 24811 18207
rect 24811 18173 24820 18207
rect 24768 18164 24820 18173
rect 22192 18096 22244 18148
rect 14924 18028 14976 18080
rect 18880 18028 18932 18080
rect 20168 18028 20220 18080
rect 22100 18028 22152 18080
rect 22744 18028 22796 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 6276 17867 6328 17876
rect 6276 17833 6285 17867
rect 6285 17833 6319 17867
rect 6319 17833 6328 17867
rect 6276 17824 6328 17833
rect 7288 17824 7340 17876
rect 8300 17756 8352 17808
rect 6920 17688 6972 17740
rect 7840 17688 7892 17740
rect 8392 17688 8444 17740
rect 9404 17688 9456 17740
rect 9772 17688 9824 17740
rect 17500 17824 17552 17876
rect 21272 17824 21324 17876
rect 12716 17799 12768 17808
rect 12716 17765 12725 17799
rect 12725 17765 12759 17799
rect 12759 17765 12768 17799
rect 12716 17756 12768 17765
rect 7288 17484 7340 17536
rect 9312 17552 9364 17604
rect 7840 17527 7892 17536
rect 7840 17493 7849 17527
rect 7849 17493 7883 17527
rect 7883 17493 7892 17527
rect 7840 17484 7892 17493
rect 9496 17527 9548 17536
rect 9496 17493 9505 17527
rect 9505 17493 9539 17527
rect 9539 17493 9548 17527
rect 9496 17484 9548 17493
rect 9588 17527 9640 17536
rect 9588 17493 9597 17527
rect 9597 17493 9631 17527
rect 9631 17493 9640 17527
rect 9588 17484 9640 17493
rect 11336 17595 11388 17604
rect 11336 17561 11345 17595
rect 11345 17561 11379 17595
rect 11379 17561 11388 17595
rect 11336 17552 11388 17561
rect 11612 17552 11664 17604
rect 14004 17688 14056 17740
rect 14280 17688 14332 17740
rect 14740 17731 14792 17740
rect 14740 17697 14749 17731
rect 14749 17697 14783 17731
rect 14783 17697 14792 17731
rect 14740 17688 14792 17697
rect 14832 17731 14884 17740
rect 14832 17697 14841 17731
rect 14841 17697 14875 17731
rect 14875 17697 14884 17731
rect 14832 17688 14884 17697
rect 16396 17688 16448 17740
rect 17132 17688 17184 17740
rect 21732 17688 21784 17740
rect 22560 17824 22612 17876
rect 22744 17824 22796 17876
rect 14924 17620 14976 17672
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 19524 17620 19576 17672
rect 24860 17663 24912 17672
rect 24860 17629 24869 17663
rect 24869 17629 24903 17663
rect 24903 17629 24912 17663
rect 24860 17620 24912 17629
rect 15384 17552 15436 17604
rect 12716 17484 12768 17536
rect 14280 17527 14332 17536
rect 14280 17493 14289 17527
rect 14289 17493 14323 17527
rect 14323 17493 14332 17527
rect 14280 17484 14332 17493
rect 15568 17484 15620 17536
rect 18880 17552 18932 17604
rect 20168 17595 20220 17604
rect 20168 17561 20177 17595
rect 20177 17561 20211 17595
rect 20211 17561 20220 17595
rect 20168 17552 20220 17561
rect 20628 17552 20680 17604
rect 22652 17552 22704 17604
rect 16580 17527 16632 17536
rect 16580 17493 16589 17527
rect 16589 17493 16623 17527
rect 16623 17493 16632 17527
rect 16580 17484 16632 17493
rect 22836 17552 22888 17604
rect 24308 17484 24360 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 4528 17280 4580 17332
rect 8300 17212 8352 17264
rect 9496 17280 9548 17332
rect 12072 17280 12124 17332
rect 14188 17280 14240 17332
rect 14832 17323 14884 17332
rect 14832 17289 14841 17323
rect 14841 17289 14875 17323
rect 14875 17289 14884 17323
rect 14832 17280 14884 17289
rect 12808 17212 12860 17264
rect 13360 17212 13412 17264
rect 19524 17280 19576 17332
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 9036 17187 9088 17196
rect 9036 17153 9045 17187
rect 9045 17153 9079 17187
rect 9079 17153 9088 17187
rect 9036 17144 9088 17153
rect 16672 17144 16724 17196
rect 17960 17212 18012 17264
rect 21088 17212 21140 17264
rect 20628 17144 20680 17196
rect 6920 17076 6972 17128
rect 10324 17076 10376 17128
rect 10508 17119 10560 17128
rect 10508 17085 10517 17119
rect 10517 17085 10551 17119
rect 10551 17085 10560 17119
rect 10508 17076 10560 17085
rect 10876 17076 10928 17128
rect 11336 17076 11388 17128
rect 13268 17076 13320 17128
rect 13360 17076 13412 17128
rect 11520 17008 11572 17060
rect 18604 17076 18656 17128
rect 18696 17076 18748 17128
rect 19340 17076 19392 17128
rect 20444 17119 20496 17128
rect 20444 17085 20453 17119
rect 20453 17085 20487 17119
rect 20487 17085 20496 17119
rect 20444 17076 20496 17085
rect 23756 17144 23808 17196
rect 24676 17119 24728 17128
rect 24676 17085 24685 17119
rect 24685 17085 24719 17119
rect 24719 17085 24728 17119
rect 24676 17076 24728 17085
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 10324 16940 10376 16992
rect 10784 16940 10836 16992
rect 15016 16940 15068 16992
rect 16580 16940 16632 16992
rect 17316 16940 17368 16992
rect 22652 17008 22704 17060
rect 23296 17008 23348 17060
rect 17960 16940 18012 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 6920 16736 6972 16788
rect 7472 16779 7524 16788
rect 7472 16745 7481 16779
rect 7481 16745 7515 16779
rect 7515 16745 7524 16779
rect 7472 16736 7524 16745
rect 8300 16736 8352 16788
rect 9036 16736 9088 16788
rect 8392 16668 8444 16720
rect 6368 16600 6420 16652
rect 8300 16600 8352 16652
rect 9220 16600 9272 16652
rect 12624 16736 12676 16788
rect 21824 16736 21876 16788
rect 10876 16668 10928 16720
rect 14372 16668 14424 16720
rect 12624 16600 12676 16652
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 15936 16643 15988 16652
rect 15936 16609 15945 16643
rect 15945 16609 15979 16643
rect 15979 16609 15988 16643
rect 15936 16600 15988 16609
rect 20168 16600 20220 16652
rect 23020 16600 23072 16652
rect 1492 16532 1544 16584
rect 9312 16532 9364 16584
rect 9588 16532 9640 16584
rect 11980 16532 12032 16584
rect 12716 16532 12768 16584
rect 20444 16575 20496 16584
rect 20444 16541 20453 16575
rect 20453 16541 20487 16575
rect 20487 16541 20496 16575
rect 20444 16532 20496 16541
rect 20536 16575 20588 16584
rect 20536 16541 20545 16575
rect 20545 16541 20579 16575
rect 20579 16541 20588 16575
rect 20536 16532 20588 16541
rect 21732 16575 21784 16584
rect 21732 16541 21741 16575
rect 21741 16541 21775 16575
rect 21775 16541 21784 16575
rect 21732 16532 21784 16541
rect 23388 16600 23440 16652
rect 1308 16464 1360 16516
rect 7472 16464 7524 16516
rect 7840 16464 7892 16516
rect 10232 16396 10284 16448
rect 19524 16464 19576 16516
rect 11704 16396 11756 16448
rect 11796 16439 11848 16448
rect 11796 16405 11805 16439
rect 11805 16405 11839 16439
rect 11839 16405 11848 16439
rect 11796 16396 11848 16405
rect 14648 16396 14700 16448
rect 16304 16396 16356 16448
rect 17500 16396 17552 16448
rect 20076 16439 20128 16448
rect 20076 16405 20085 16439
rect 20085 16405 20119 16439
rect 20119 16405 20128 16439
rect 20076 16396 20128 16405
rect 21180 16396 21232 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 7288 16192 7340 16244
rect 10508 16192 10560 16244
rect 10600 16235 10652 16244
rect 10600 16201 10609 16235
rect 10609 16201 10643 16235
rect 10643 16201 10652 16235
rect 10600 16192 10652 16201
rect 10968 16192 11020 16244
rect 12532 16192 12584 16244
rect 13452 16192 13504 16244
rect 16396 16235 16448 16244
rect 16396 16201 16405 16235
rect 16405 16201 16439 16235
rect 16439 16201 16448 16235
rect 16396 16192 16448 16201
rect 2504 16167 2556 16176
rect 2504 16133 2513 16167
rect 2513 16133 2547 16167
rect 2547 16133 2556 16167
rect 2504 16124 2556 16133
rect 7472 16124 7524 16176
rect 11796 16124 11848 16176
rect 14280 16124 14332 16176
rect 6552 16056 6604 16108
rect 8300 15988 8352 16040
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 10416 16056 10468 16108
rect 12808 16056 12860 16108
rect 14188 16099 14240 16108
rect 14188 16065 14197 16099
rect 14197 16065 14231 16099
rect 14231 16065 14240 16099
rect 14188 16056 14240 16065
rect 15752 16056 15804 16108
rect 16304 16056 16356 16108
rect 17132 16167 17184 16176
rect 17132 16133 17141 16167
rect 17141 16133 17175 16167
rect 17175 16133 17184 16167
rect 17132 16124 17184 16133
rect 17868 16124 17920 16176
rect 18604 16235 18656 16244
rect 18604 16201 18613 16235
rect 18613 16201 18647 16235
rect 18647 16201 18656 16235
rect 18604 16192 18656 16201
rect 19248 16235 19300 16244
rect 19248 16201 19257 16235
rect 19257 16201 19291 16235
rect 19291 16201 19300 16235
rect 19248 16192 19300 16201
rect 20076 16192 20128 16244
rect 22836 16192 22888 16244
rect 16580 16056 16632 16108
rect 18144 16056 18196 16108
rect 1768 15852 1820 15904
rect 10232 15988 10284 16040
rect 11888 15988 11940 16040
rect 15476 15988 15528 16040
rect 10968 15920 11020 15972
rect 14004 15920 14056 15972
rect 22100 16124 22152 16176
rect 22468 16124 22520 16176
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 24216 16056 24268 16108
rect 21548 15988 21600 16040
rect 22744 15988 22796 16040
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 22560 15920 22612 15972
rect 12348 15852 12400 15904
rect 12624 15852 12676 15904
rect 14280 15895 14332 15904
rect 14280 15861 14289 15895
rect 14289 15861 14323 15895
rect 14323 15861 14332 15895
rect 14280 15852 14332 15861
rect 15200 15852 15252 15904
rect 21916 15852 21968 15904
rect 22100 15852 22152 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 7472 15648 7524 15700
rect 9312 15648 9364 15700
rect 11704 15648 11756 15700
rect 17224 15648 17276 15700
rect 20812 15648 20864 15700
rect 20996 15648 21048 15700
rect 22100 15648 22152 15700
rect 12440 15580 12492 15632
rect 19892 15580 19944 15632
rect 19984 15580 20036 15632
rect 11336 15512 11388 15564
rect 14096 15512 14148 15564
rect 17408 15512 17460 15564
rect 21180 15512 21232 15564
rect 12624 15444 12676 15496
rect 13452 15487 13504 15496
rect 13452 15453 13461 15487
rect 13461 15453 13495 15487
rect 13495 15453 13504 15487
rect 13452 15444 13504 15453
rect 14648 15487 14700 15496
rect 14648 15453 14657 15487
rect 14657 15453 14691 15487
rect 14691 15453 14700 15487
rect 14648 15444 14700 15453
rect 16120 15444 16172 15496
rect 19984 15444 20036 15496
rect 22284 15444 22336 15496
rect 24308 15444 24360 15496
rect 10968 15376 11020 15428
rect 10232 15308 10284 15360
rect 14096 15376 14148 15428
rect 12716 15308 12768 15360
rect 15660 15308 15712 15360
rect 16672 15308 16724 15360
rect 18696 15351 18748 15360
rect 18696 15317 18705 15351
rect 18705 15317 18739 15351
rect 18739 15317 18748 15351
rect 18696 15308 18748 15317
rect 21272 15376 21324 15428
rect 19616 15308 19668 15360
rect 20628 15351 20680 15360
rect 20628 15317 20637 15351
rect 20637 15317 20671 15351
rect 20671 15317 20680 15351
rect 20628 15308 20680 15317
rect 20812 15308 20864 15360
rect 24952 15376 25004 15428
rect 21548 15308 21600 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 2688 15104 2740 15156
rect 8576 15104 8628 15156
rect 9312 15104 9364 15156
rect 9404 15079 9456 15088
rect 9404 15045 9413 15079
rect 9413 15045 9447 15079
rect 9447 15045 9456 15079
rect 9404 15036 9456 15045
rect 9772 15104 9824 15156
rect 10968 15036 11020 15088
rect 12164 15104 12216 15156
rect 17040 15104 17092 15156
rect 18696 15104 18748 15156
rect 18880 15147 18932 15156
rect 18880 15113 18889 15147
rect 18889 15113 18923 15147
rect 18923 15113 18932 15147
rect 18880 15104 18932 15113
rect 22376 15104 22428 15156
rect 11980 15036 12032 15088
rect 12624 15036 12676 15088
rect 13452 15079 13504 15088
rect 13452 15045 13461 15079
rect 13461 15045 13495 15079
rect 13495 15045 13504 15079
rect 13452 15036 13504 15045
rect 16672 15036 16724 15088
rect 16764 15036 16816 15088
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 13820 14900 13872 14952
rect 14832 14943 14884 14952
rect 14832 14909 14841 14943
rect 14841 14909 14875 14943
rect 14875 14909 14884 14943
rect 14832 14900 14884 14909
rect 16028 14968 16080 15020
rect 18604 14968 18656 15020
rect 16120 14900 16172 14952
rect 19800 15011 19852 15020
rect 19800 14977 19809 15011
rect 19809 14977 19843 15011
rect 19843 14977 19852 15011
rect 19800 14968 19852 14977
rect 23848 14968 23900 15020
rect 24676 14943 24728 14952
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 16856 14832 16908 14884
rect 17500 14832 17552 14884
rect 20812 14832 20864 14884
rect 9956 14764 10008 14816
rect 13268 14764 13320 14816
rect 13728 14764 13780 14816
rect 16672 14764 16724 14816
rect 19340 14764 19392 14816
rect 20444 14764 20496 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 9864 14560 9916 14612
rect 10784 14560 10836 14612
rect 11336 14492 11388 14544
rect 11980 14535 12032 14544
rect 11980 14501 11989 14535
rect 11989 14501 12023 14535
rect 12023 14501 12032 14535
rect 11980 14492 12032 14501
rect 12808 14560 12860 14612
rect 15292 14560 15344 14612
rect 14556 14492 14608 14544
rect 17132 14603 17184 14612
rect 17132 14569 17141 14603
rect 17141 14569 17175 14603
rect 17175 14569 17184 14603
rect 17132 14560 17184 14569
rect 19432 14492 19484 14544
rect 9956 14467 10008 14476
rect 9956 14433 9965 14467
rect 9965 14433 9999 14467
rect 9999 14433 10008 14467
rect 9956 14424 10008 14433
rect 12624 14424 12676 14476
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 14740 14424 14792 14476
rect 15384 14467 15436 14476
rect 15384 14433 15393 14467
rect 15393 14433 15427 14467
rect 15427 14433 15436 14467
rect 15384 14424 15436 14433
rect 16396 14424 16448 14476
rect 21180 14467 21232 14476
rect 21180 14433 21189 14467
rect 21189 14433 21223 14467
rect 21223 14433 21232 14467
rect 21180 14424 21232 14433
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 19524 14356 19576 14408
rect 10232 14331 10284 14340
rect 10232 14297 10241 14331
rect 10241 14297 10275 14331
rect 10275 14297 10284 14331
rect 10232 14288 10284 14297
rect 13360 14331 13412 14340
rect 13360 14297 13369 14331
rect 13369 14297 13403 14331
rect 13403 14297 13412 14331
rect 13360 14288 13412 14297
rect 9864 14220 9916 14272
rect 10876 14220 10928 14272
rect 15936 14288 15988 14340
rect 15568 14220 15620 14272
rect 16396 14220 16448 14272
rect 16488 14220 16540 14272
rect 21088 14288 21140 14340
rect 23388 14288 23440 14340
rect 18512 14220 18564 14272
rect 19432 14263 19484 14272
rect 19432 14229 19441 14263
rect 19441 14229 19475 14263
rect 19475 14229 19484 14263
rect 19432 14220 19484 14229
rect 19984 14263 20036 14272
rect 19984 14229 19993 14263
rect 19993 14229 20027 14263
rect 20027 14229 20036 14263
rect 19984 14220 20036 14229
rect 20260 14220 20312 14272
rect 21824 14220 21876 14272
rect 22928 14263 22980 14272
rect 22928 14229 22937 14263
rect 22937 14229 22971 14263
rect 22971 14229 22980 14263
rect 22928 14220 22980 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 9956 14016 10008 14068
rect 10140 14016 10192 14068
rect 10784 14016 10836 14068
rect 12164 14016 12216 14068
rect 13728 14016 13780 14068
rect 17592 14016 17644 14068
rect 19616 14016 19668 14068
rect 21180 14016 21232 14068
rect 21456 14016 21508 14068
rect 23388 14016 23440 14068
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 1860 13880 1912 13932
rect 5448 13880 5500 13932
rect 9772 13948 9824 14000
rect 11244 13948 11296 14000
rect 17408 13991 17460 14000
rect 17408 13957 17417 13991
rect 17417 13957 17451 13991
rect 17451 13957 17460 13991
rect 17408 13948 17460 13957
rect 19984 13948 20036 14000
rect 20720 13948 20772 14000
rect 9588 13880 9640 13932
rect 10416 13880 10468 13932
rect 16580 13880 16632 13932
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 18512 13880 18564 13932
rect 1308 13812 1360 13864
rect 9496 13812 9548 13864
rect 11796 13744 11848 13796
rect 13452 13812 13504 13864
rect 19156 13812 19208 13864
rect 20352 13880 20404 13932
rect 21180 13923 21232 13932
rect 21180 13889 21189 13923
rect 21189 13889 21223 13923
rect 21223 13889 21232 13923
rect 21180 13880 21232 13889
rect 21732 13948 21784 14000
rect 22192 13948 22244 14000
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 20168 13812 20220 13864
rect 20536 13812 20588 13864
rect 21364 13812 21416 13864
rect 23756 13812 23808 13864
rect 9864 13676 9916 13728
rect 22008 13676 22060 13728
rect 22928 13676 22980 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 5816 13472 5868 13524
rect 6552 13336 6604 13388
rect 6828 13379 6880 13388
rect 6828 13345 6837 13379
rect 6837 13345 6871 13379
rect 6871 13345 6880 13379
rect 6828 13336 6880 13345
rect 7104 13379 7156 13388
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 7564 13336 7616 13388
rect 9772 13404 9824 13456
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 11520 13472 11572 13524
rect 11980 13515 12032 13524
rect 11980 13481 11989 13515
rect 11989 13481 12023 13515
rect 12023 13481 12032 13515
rect 11980 13472 12032 13481
rect 12348 13515 12400 13524
rect 12348 13481 12357 13515
rect 12357 13481 12391 13515
rect 12391 13481 12400 13515
rect 12348 13472 12400 13481
rect 13728 13472 13780 13524
rect 12716 13336 12768 13388
rect 15384 13336 15436 13388
rect 15936 13472 15988 13524
rect 20352 13472 20404 13524
rect 18328 13404 18380 13456
rect 18880 13404 18932 13456
rect 19156 13404 19208 13456
rect 6460 13132 6512 13184
rect 18512 13336 18564 13388
rect 19892 13379 19944 13388
rect 19892 13345 19901 13379
rect 19901 13345 19935 13379
rect 19935 13345 19944 13379
rect 19892 13336 19944 13345
rect 11612 13200 11664 13252
rect 11980 13200 12032 13252
rect 14464 13200 14516 13252
rect 8760 13132 8812 13184
rect 19432 13268 19484 13320
rect 22652 13311 22704 13320
rect 22652 13277 22661 13311
rect 22661 13277 22695 13311
rect 22695 13277 22704 13311
rect 22652 13268 22704 13277
rect 14832 13243 14884 13252
rect 14832 13209 14841 13243
rect 14841 13209 14875 13243
rect 14875 13209 14884 13243
rect 14832 13200 14884 13209
rect 16488 13200 16540 13252
rect 18328 13200 18380 13252
rect 25688 13200 25740 13252
rect 15476 13132 15528 13184
rect 17224 13132 17276 13184
rect 17776 13175 17828 13184
rect 17776 13141 17785 13175
rect 17785 13141 17819 13175
rect 17819 13141 17828 13175
rect 17776 13132 17828 13141
rect 19800 13132 19852 13184
rect 21364 13132 21416 13184
rect 22008 13132 22060 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 8668 12971 8720 12980
rect 8668 12937 8677 12971
rect 8677 12937 8711 12971
rect 8711 12937 8720 12971
rect 8668 12928 8720 12937
rect 11796 12928 11848 12980
rect 12532 12928 12584 12980
rect 12716 12928 12768 12980
rect 15752 12928 15804 12980
rect 16488 12971 16540 12980
rect 16488 12937 16497 12971
rect 16497 12937 16531 12971
rect 16531 12937 16540 12971
rect 16488 12928 16540 12937
rect 17224 12971 17276 12980
rect 17224 12937 17233 12971
rect 17233 12937 17267 12971
rect 17267 12937 17276 12971
rect 17224 12928 17276 12937
rect 18512 12928 18564 12980
rect 6552 12792 6604 12844
rect 9680 12860 9732 12912
rect 9956 12860 10008 12912
rect 11612 12903 11664 12912
rect 11612 12869 11621 12903
rect 11621 12869 11655 12903
rect 11655 12869 11664 12903
rect 11612 12860 11664 12869
rect 14372 12860 14424 12912
rect 17040 12860 17092 12912
rect 18880 12860 18932 12912
rect 21364 12860 21416 12912
rect 13636 12792 13688 12844
rect 13820 12792 13872 12844
rect 15936 12792 15988 12844
rect 8760 12767 8812 12776
rect 8760 12733 8769 12767
rect 8769 12733 8803 12767
rect 8803 12733 8812 12767
rect 22836 12835 22888 12844
rect 22836 12801 22845 12835
rect 22845 12801 22879 12835
rect 22879 12801 22888 12835
rect 22836 12792 22888 12801
rect 23296 12792 23348 12844
rect 8760 12724 8812 12733
rect 19524 12724 19576 12776
rect 21824 12724 21876 12776
rect 22008 12767 22060 12776
rect 22008 12733 22017 12767
rect 22017 12733 22051 12767
rect 22051 12733 22060 12767
rect 22008 12724 22060 12733
rect 24768 12767 24820 12776
rect 24768 12733 24777 12767
rect 24777 12733 24811 12767
rect 24811 12733 24820 12767
rect 24768 12724 24820 12733
rect 14372 12656 14424 12708
rect 14648 12699 14700 12708
rect 14648 12665 14657 12699
rect 14657 12665 14691 12699
rect 14691 12665 14700 12699
rect 14648 12656 14700 12665
rect 16212 12656 16264 12708
rect 10968 12588 11020 12640
rect 17684 12588 17736 12640
rect 18604 12631 18656 12640
rect 18604 12597 18613 12631
rect 18613 12597 18647 12631
rect 18647 12597 18656 12631
rect 18604 12588 18656 12597
rect 24584 12588 24636 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 8944 12384 8996 12436
rect 10140 12384 10192 12436
rect 12164 12384 12216 12436
rect 12348 12384 12400 12436
rect 13820 12384 13872 12436
rect 14464 12427 14516 12436
rect 14464 12393 14473 12427
rect 14473 12393 14507 12427
rect 14507 12393 14516 12427
rect 14464 12384 14516 12393
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 15660 12384 15712 12393
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 14004 12248 14056 12300
rect 15660 12248 15712 12300
rect 9680 12180 9732 12232
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 17408 12384 17460 12436
rect 17500 12384 17552 12436
rect 23296 12316 23348 12368
rect 16120 12248 16172 12300
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 19984 12248 20036 12300
rect 21272 12248 21324 12300
rect 21824 12248 21876 12300
rect 21916 12248 21968 12300
rect 19340 12180 19392 12232
rect 22008 12180 22060 12232
rect 10232 12112 10284 12164
rect 12072 12112 12124 12164
rect 14188 12112 14240 12164
rect 17316 12112 17368 12164
rect 3516 12044 3568 12096
rect 9588 12044 9640 12096
rect 13176 12044 13228 12096
rect 14924 12087 14976 12096
rect 14924 12053 14933 12087
rect 14933 12053 14967 12087
rect 14967 12053 14976 12087
rect 14924 12044 14976 12053
rect 15292 12044 15344 12096
rect 15384 12044 15436 12096
rect 18328 12044 18380 12096
rect 19892 12044 19944 12096
rect 21088 12087 21140 12096
rect 21088 12053 21097 12087
rect 21097 12053 21131 12087
rect 21131 12053 21140 12087
rect 21088 12044 21140 12053
rect 24860 12044 24912 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 12348 11840 12400 11892
rect 5172 11772 5224 11824
rect 10692 11772 10744 11824
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 11520 11704 11572 11756
rect 14188 11704 14240 11756
rect 14740 11704 14792 11756
rect 16488 11840 16540 11892
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 19524 11840 19576 11892
rect 19984 11883 20036 11892
rect 19984 11849 19993 11883
rect 19993 11849 20027 11883
rect 20027 11849 20036 11883
rect 19984 11840 20036 11849
rect 18512 11815 18564 11824
rect 18512 11781 18521 11815
rect 18521 11781 18555 11815
rect 18555 11781 18564 11815
rect 18512 11772 18564 11781
rect 20720 11772 20772 11824
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 13176 11636 13228 11688
rect 19892 11704 19944 11756
rect 17408 11636 17460 11688
rect 20444 11636 20496 11688
rect 15752 11500 15804 11552
rect 16764 11500 16816 11552
rect 22560 11704 22612 11756
rect 22100 11568 22152 11620
rect 21364 11500 21416 11552
rect 24492 11500 24544 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 15476 11339 15528 11348
rect 15476 11305 15485 11339
rect 15485 11305 15519 11339
rect 15519 11305 15528 11339
rect 15476 11296 15528 11305
rect 16672 11296 16724 11348
rect 16856 11296 16908 11348
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 15660 11160 15712 11212
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 17592 11092 17644 11144
rect 20628 11024 20680 11076
rect 20812 11067 20864 11076
rect 20812 11033 20821 11067
rect 20821 11033 20855 11067
rect 20855 11033 20864 11067
rect 20812 11024 20864 11033
rect 23848 11024 23900 11076
rect 19616 10999 19668 11008
rect 19616 10965 19625 10999
rect 19625 10965 19659 10999
rect 19659 10965 19668 10999
rect 19616 10956 19668 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 19616 10752 19668 10804
rect 10968 10684 11020 10736
rect 12072 10659 12124 10668
rect 12072 10625 12081 10659
rect 12081 10625 12115 10659
rect 12115 10625 12124 10659
rect 12072 10616 12124 10625
rect 17684 10684 17736 10736
rect 15752 10616 15804 10668
rect 17776 10548 17828 10600
rect 19984 10548 20036 10600
rect 21548 10548 21600 10600
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 12532 10480 12584 10532
rect 20812 10480 20864 10532
rect 5264 10412 5316 10464
rect 9864 10412 9916 10464
rect 18236 10455 18288 10464
rect 18236 10421 18245 10455
rect 18245 10421 18279 10455
rect 18279 10421 18288 10455
rect 18236 10412 18288 10421
rect 21732 10412 21784 10464
rect 23940 10412 23992 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 22560 10140 22612 10192
rect 18236 10072 18288 10124
rect 13636 10004 13688 10056
rect 19432 10004 19484 10056
rect 19800 10004 19852 10056
rect 18420 9936 18472 9988
rect 24952 10004 25004 10056
rect 16856 9911 16908 9920
rect 16856 9877 16865 9911
rect 16865 9877 16899 9911
rect 16899 9877 16908 9911
rect 16856 9868 16908 9877
rect 23296 9936 23348 9988
rect 24032 9868 24084 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 9496 9596 9548 9648
rect 13912 9596 13964 9648
rect 15568 9596 15620 9648
rect 18696 9596 18748 9648
rect 21088 9528 21140 9580
rect 23848 9528 23900 9580
rect 5540 9460 5592 9512
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 24676 9503 24728 9512
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 6552 9435 6604 9444
rect 6552 9401 6561 9435
rect 6561 9401 6595 9435
rect 6595 9401 6604 9435
rect 6552 9392 6604 9401
rect 17684 9392 17736 9444
rect 23848 9392 23900 9444
rect 7104 9324 7156 9376
rect 11704 9324 11756 9376
rect 22744 9367 22796 9376
rect 22744 9333 22753 9367
rect 22753 9333 22787 9367
rect 22787 9333 22796 9367
rect 22744 9324 22796 9333
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 3056 9120 3108 9172
rect 5908 9120 5960 9172
rect 22836 9052 22888 9104
rect 7748 8916 7800 8968
rect 15016 8916 15068 8968
rect 21732 8959 21784 8968
rect 21732 8925 21741 8959
rect 21741 8925 21775 8959
rect 21775 8925 21784 8959
rect 21732 8916 21784 8925
rect 23388 8916 23440 8968
rect 24584 8916 24636 8968
rect 23296 8780 23348 8832
rect 23480 8780 23532 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18880 8508 18932 8560
rect 20904 8508 20956 8560
rect 25136 8551 25188 8560
rect 25136 8517 25145 8551
rect 25145 8517 25179 8551
rect 25179 8517 25188 8551
rect 25136 8508 25188 8517
rect 21272 8372 21324 8424
rect 22376 8372 22428 8424
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 24952 8372 25004 8424
rect 11612 8304 11664 8356
rect 18420 8304 18472 8356
rect 22008 8304 22060 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 6460 8075 6512 8084
rect 6460 8041 6469 8075
rect 6469 8041 6503 8075
rect 6503 8041 6512 8075
rect 6460 8032 6512 8041
rect 11888 8032 11940 8084
rect 12716 8032 12768 8084
rect 6828 7896 6880 7948
rect 23388 7939 23440 7948
rect 23388 7905 23397 7939
rect 23397 7905 23431 7939
rect 23431 7905 23440 7939
rect 23388 7896 23440 7905
rect 6460 7828 6512 7880
rect 20444 7871 20496 7880
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 20628 7828 20680 7880
rect 23480 7828 23532 7880
rect 24860 7871 24912 7880
rect 24860 7837 24869 7871
rect 24869 7837 24903 7871
rect 24903 7837 24912 7871
rect 24860 7828 24912 7837
rect 2780 7760 2832 7812
rect 9128 7760 9180 7812
rect 20812 7692 20864 7744
rect 21088 7735 21140 7744
rect 21088 7701 21097 7735
rect 21097 7701 21131 7735
rect 21131 7701 21140 7735
rect 21088 7692 21140 7701
rect 24124 7692 24176 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 17316 7420 17368 7472
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 20904 7352 20956 7404
rect 22008 7352 22060 7404
rect 23940 7395 23992 7404
rect 23940 7361 23949 7395
rect 23949 7361 23983 7395
rect 23983 7361 23992 7395
rect 23940 7352 23992 7361
rect 22192 7284 22244 7336
rect 22284 7284 22336 7336
rect 20628 7216 20680 7268
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 16488 6740 16540 6792
rect 20812 6783 20864 6792
rect 20812 6749 20821 6783
rect 20821 6749 20855 6783
rect 20855 6749 20864 6783
rect 20812 6740 20864 6749
rect 22836 6783 22888 6792
rect 22836 6749 22845 6783
rect 22845 6749 22879 6783
rect 22879 6749 22888 6783
rect 22836 6740 22888 6749
rect 3056 6672 3108 6724
rect 6000 6672 6052 6724
rect 22008 6715 22060 6724
rect 22008 6681 22017 6715
rect 22017 6681 22051 6715
rect 22051 6681 22060 6715
rect 22008 6672 22060 6681
rect 24952 6672 25004 6724
rect 18512 6604 18564 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 11244 6332 11296 6384
rect 16396 6332 16448 6384
rect 22652 6332 22704 6384
rect 25136 6375 25188 6384
rect 25136 6341 25145 6375
rect 25145 6341 25179 6375
rect 25179 6341 25188 6375
rect 25136 6332 25188 6341
rect 18420 6307 18472 6316
rect 18420 6273 18429 6307
rect 18429 6273 18463 6307
rect 18463 6273 18472 6307
rect 18420 6264 18472 6273
rect 21088 6264 21140 6316
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 24032 6307 24084 6316
rect 24032 6273 24041 6307
rect 24041 6273 24075 6307
rect 24075 6273 24084 6307
rect 24032 6264 24084 6273
rect 21916 6196 21968 6248
rect 22836 6128 22888 6180
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 20904 5856 20956 5908
rect 20720 5720 20772 5772
rect 21548 5720 21600 5772
rect 2596 5652 2648 5704
rect 8760 5652 8812 5704
rect 20536 5695 20588 5704
rect 20536 5661 20545 5695
rect 20545 5661 20579 5695
rect 20579 5661 20588 5695
rect 20536 5652 20588 5661
rect 20628 5652 20680 5704
rect 22560 5652 22612 5704
rect 10048 5584 10100 5636
rect 15108 5584 15160 5636
rect 9312 5516 9364 5568
rect 11428 5516 11480 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 19616 5244 19668 5296
rect 17776 5219 17828 5228
rect 17776 5185 17785 5219
rect 17785 5185 17819 5219
rect 17819 5185 17828 5219
rect 17776 5176 17828 5185
rect 19524 5219 19576 5228
rect 19524 5185 19533 5219
rect 19533 5185 19567 5219
rect 19567 5185 19576 5219
rect 19524 5176 19576 5185
rect 21824 5176 21876 5228
rect 24124 5219 24176 5228
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 19340 5108 19392 5160
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 22468 5108 22520 5117
rect 24768 5151 24820 5160
rect 24768 5117 24777 5151
rect 24777 5117 24811 5151
rect 24811 5117 24820 5151
rect 24768 5108 24820 5117
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 17776 4700 17828 4752
rect 19892 4675 19944 4684
rect 19892 4641 19901 4675
rect 19901 4641 19935 4675
rect 19935 4641 19944 4675
rect 19892 4632 19944 4641
rect 18512 4564 18564 4616
rect 18604 4564 18656 4616
rect 19708 4564 19760 4616
rect 22744 4632 22796 4684
rect 24860 4743 24912 4752
rect 24860 4709 24869 4743
rect 24869 4709 24903 4743
rect 24903 4709 24912 4743
rect 24860 4700 24912 4709
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 23296 4564 23348 4616
rect 20628 4496 20680 4548
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 8208 4156 8260 4208
rect 10324 4156 10376 4208
rect 12624 4156 12676 4208
rect 14188 4156 14240 4208
rect 13452 4088 13504 4140
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 16672 4088 16724 4140
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 22100 4131 22152 4140
rect 22100 4097 22109 4131
rect 22109 4097 22143 4131
rect 22143 4097 22152 4131
rect 22100 4088 22152 4097
rect 23848 4131 23900 4140
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 3148 4020 3200 4072
rect 6184 4020 6236 4072
rect 11612 4020 11664 4072
rect 2780 3952 2832 4004
rect 9036 3952 9088 4004
rect 2872 3884 2924 3936
rect 6092 3884 6144 3936
rect 9404 3884 9456 3936
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 10508 3884 10560 3936
rect 16396 4020 16448 4072
rect 17500 4020 17552 4072
rect 20076 4020 20128 4072
rect 13452 3952 13504 4004
rect 16304 3995 16356 4004
rect 16304 3961 16313 3995
rect 16313 3961 16347 3995
rect 16347 3961 16356 3995
rect 16304 3952 16356 3961
rect 21180 3952 21232 4004
rect 15936 3884 15988 3936
rect 19616 3884 19668 3936
rect 22376 3884 22428 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 6736 3723 6788 3732
rect 6736 3689 6745 3723
rect 6745 3689 6779 3723
rect 6779 3689 6788 3723
rect 6736 3680 6788 3689
rect 8208 3723 8260 3732
rect 8208 3689 8217 3723
rect 8217 3689 8251 3723
rect 8251 3689 8260 3723
rect 8208 3680 8260 3689
rect 9496 3680 9548 3732
rect 10048 3723 10100 3732
rect 10048 3689 10057 3723
rect 10057 3689 10091 3723
rect 10091 3689 10100 3723
rect 10048 3680 10100 3689
rect 22836 3680 22888 3732
rect 24952 3680 25004 3732
rect 5540 3612 5592 3664
rect 16120 3612 16172 3664
rect 16580 3612 16632 3664
rect 8300 3544 8352 3596
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 12716 3544 12768 3596
rect 14924 3544 14976 3596
rect 16028 3544 16080 3596
rect 1676 3476 1728 3528
rect 3332 3408 3384 3460
rect 6092 3519 6144 3528
rect 6092 3485 6101 3519
rect 6101 3485 6135 3519
rect 6135 3485 6144 3519
rect 6092 3476 6144 3485
rect 6460 3476 6512 3528
rect 9404 3476 9456 3528
rect 9772 3476 9824 3528
rect 10876 3476 10928 3528
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 15108 3519 15160 3528
rect 15108 3485 15117 3519
rect 15117 3485 15151 3519
rect 15151 3485 15160 3519
rect 15108 3476 15160 3485
rect 16212 3476 16264 3528
rect 17868 3544 17920 3596
rect 20996 3476 21048 3528
rect 18972 3408 19024 3460
rect 2044 3340 2096 3392
rect 2780 3340 2832 3392
rect 3424 3340 3476 3392
rect 3884 3340 3936 3392
rect 4988 3340 5040 3392
rect 6828 3340 6880 3392
rect 7840 3340 7892 3392
rect 8668 3383 8720 3392
rect 8668 3349 8677 3383
rect 8677 3349 8711 3383
rect 8711 3349 8720 3383
rect 8668 3340 8720 3349
rect 11244 3340 11296 3392
rect 22008 3340 22060 3392
rect 22836 3340 22888 3392
rect 23572 3340 23624 3392
rect 24124 3340 24176 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 2688 3179 2740 3188
rect 2688 3145 2697 3179
rect 2697 3145 2731 3179
rect 2731 3145 2740 3179
rect 2688 3136 2740 3145
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 5908 3179 5960 3188
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 7196 3136 7248 3188
rect 8484 3179 8536 3188
rect 8484 3145 8493 3179
rect 8493 3145 8527 3179
rect 8527 3145 8536 3179
rect 8484 3136 8536 3145
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 24676 3136 24728 3188
rect 2044 3000 2096 3052
rect 2780 3000 2832 3052
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 5356 3000 5408 3052
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 8208 3000 8260 3052
rect 8668 3000 8720 3052
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 14832 3068 14884 3120
rect 18604 3068 18656 3120
rect 19892 3068 19944 3120
rect 23572 3111 23624 3120
rect 23572 3077 23581 3111
rect 23581 3077 23615 3111
rect 23615 3077 23624 3111
rect 23572 3068 23624 3077
rect 11244 3000 11296 3052
rect 12624 3043 12676 3052
rect 12624 3009 12633 3043
rect 12633 3009 12667 3043
rect 12667 3009 12676 3043
rect 12624 3000 12676 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 16764 3000 16816 3052
rect 16948 3000 17000 3052
rect 3332 2932 3384 2984
rect 9036 2975 9088 2984
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 10508 2932 10560 2984
rect 13360 2975 13412 2984
rect 13360 2941 13369 2975
rect 13369 2941 13403 2975
rect 13403 2941 13412 2975
rect 13360 2932 13412 2941
rect 14188 2932 14240 2984
rect 15660 2932 15712 2984
rect 4896 2864 4948 2916
rect 17132 2864 17184 2916
rect 20628 2864 20680 2916
rect 23388 2864 23440 2916
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 4252 2796 4304 2848
rect 6460 2839 6512 2848
rect 6460 2805 6469 2839
rect 6469 2805 6503 2839
rect 6503 2805 6512 2839
rect 6460 2796 6512 2805
rect 16764 2796 16816 2848
rect 19892 2796 19944 2848
rect 20812 2796 20864 2848
rect 22468 2796 22520 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 1860 2635 1912 2644
rect 1860 2601 1869 2635
rect 1869 2601 1903 2635
rect 1903 2601 1912 2635
rect 1860 2592 1912 2601
rect 2596 2635 2648 2644
rect 2596 2601 2605 2635
rect 2605 2601 2639 2635
rect 2639 2601 2648 2635
rect 2596 2592 2648 2601
rect 4160 2635 4212 2644
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 7104 2635 7156 2644
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 11796 2592 11848 2644
rect 4804 2524 4856 2576
rect 8944 2524 8996 2576
rect 7748 2456 7800 2508
rect 12808 2524 12860 2576
rect 1492 2388 1544 2440
rect 2320 2388 2372 2440
rect 3884 2388 3936 2440
rect 4252 2388 4304 2440
rect 4620 2388 4672 2440
rect 7196 2388 7248 2440
rect 7564 2388 7616 2440
rect 10140 2388 10192 2440
rect 11980 2456 12032 2508
rect 14556 2456 14608 2508
rect 15292 2456 15344 2508
rect 17684 2456 17736 2508
rect 3516 2320 3568 2372
rect 5724 2320 5776 2372
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 14648 2431 14700 2440
rect 14648 2397 14657 2431
rect 14657 2397 14691 2431
rect 14691 2397 14700 2431
rect 14648 2388 14700 2397
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19892 2499 19944 2508
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 12348 2320 12400 2372
rect 13820 2320 13872 2372
rect 18328 2320 18380 2372
rect 25320 2431 25372 2440
rect 25320 2397 25329 2431
rect 25329 2397 25363 2431
rect 25363 2397 25372 2431
rect 25320 2388 25372 2397
rect 15384 2252 15436 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 3148 2048 3200 2100
rect 9036 2048 9088 2100
rect 8300 1980 8352 2032
rect 15936 1980 15988 2032
<< metal2 >>
rect 1490 56200 1546 57000
rect 1858 56200 1914 57000
rect 2226 56200 2282 57000
rect 2594 56200 2650 57000
rect 2962 56200 3018 57000
rect 3330 56200 3386 57000
rect 3698 56200 3754 57000
rect 4066 56200 4122 57000
rect 4434 56200 4490 57000
rect 4802 56200 4858 57000
rect 5170 56200 5226 57000
rect 5538 56200 5594 57000
rect 5906 56200 5962 57000
rect 6274 56200 6330 57000
rect 6642 56200 6698 57000
rect 7010 56200 7066 57000
rect 7378 56200 7434 57000
rect 7746 56200 7802 57000
rect 7852 56222 8064 56250
rect 1306 53000 1362 53009
rect 1306 52935 1362 52944
rect 1320 52630 1348 52935
rect 1308 52624 1360 52630
rect 1308 52566 1360 52572
rect 1306 50552 1362 50561
rect 1306 50487 1362 50496
rect 1320 50386 1348 50487
rect 1308 50380 1360 50386
rect 1308 50322 1360 50328
rect 1504 49298 1532 56200
rect 1872 52902 1900 56200
rect 1860 52896 1912 52902
rect 1860 52838 1912 52844
rect 2240 52698 2268 56200
rect 2608 52986 2636 56200
rect 2778 55448 2834 55457
rect 2778 55383 2834 55392
rect 2792 53242 2820 55383
rect 2976 55214 3004 56200
rect 2884 55186 3004 55214
rect 2780 53236 2832 53242
rect 2780 53178 2832 53184
rect 2608 52958 2820 52986
rect 2228 52692 2280 52698
rect 2228 52634 2280 52640
rect 2792 50862 2820 52958
rect 2884 51474 2912 55186
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 3344 51950 3372 56200
rect 3516 52896 3568 52902
rect 3516 52838 3568 52844
rect 3424 52692 3476 52698
rect 3424 52634 3476 52640
rect 3332 51944 3384 51950
rect 3332 51886 3384 51892
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 2872 51468 2924 51474
rect 2872 51410 2924 51416
rect 2780 50856 2832 50862
rect 2780 50798 2832 50804
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 3436 50318 3464 52634
rect 3424 50312 3476 50318
rect 3424 50254 3476 50260
rect 3528 49910 3556 52838
rect 3712 52562 3740 56200
rect 4080 52986 4108 56200
rect 4448 53174 4476 56200
rect 4528 54188 4580 54194
rect 4528 54130 4580 54136
rect 4620 54188 4672 54194
rect 4620 54130 4672 54136
rect 4436 53168 4488 53174
rect 4436 53110 4488 53116
rect 3976 52964 4028 52970
rect 4080 52958 4292 52986
rect 3976 52906 4028 52912
rect 3792 52624 3844 52630
rect 3792 52566 3844 52572
rect 3700 52556 3752 52562
rect 3700 52498 3752 52504
rect 3804 51610 3832 52566
rect 3792 51604 3844 51610
rect 3792 51546 3844 51552
rect 3516 49904 3568 49910
rect 3516 49846 3568 49852
rect 3332 49836 3384 49842
rect 3332 49778 3384 49784
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 1492 49292 1544 49298
rect 1492 49234 1544 49240
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 1306 48104 1362 48113
rect 1306 48039 1308 48048
rect 1360 48039 1362 48048
rect 1308 48010 1360 48016
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 1308 45960 1360 45966
rect 1308 45902 1360 45908
rect 1320 45665 1348 45902
rect 1306 45656 1362 45665
rect 1306 45591 1308 45600
rect 1360 45591 1362 45600
rect 1308 45562 1360 45568
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 1308 43308 1360 43314
rect 1308 43250 1360 43256
rect 1320 43217 1348 43250
rect 1306 43208 1362 43217
rect 1306 43143 1362 43152
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 3344 41274 3372 49778
rect 3988 49638 4016 52906
rect 4160 50924 4212 50930
rect 4160 50866 4212 50872
rect 3976 49632 4028 49638
rect 3976 49574 4028 49580
rect 3976 43172 4028 43178
rect 3976 43114 4028 43120
rect 3332 41268 3384 41274
rect 3332 41210 3384 41216
rect 1308 41132 1360 41138
rect 1308 41074 1360 41080
rect 1320 40769 1348 41074
rect 1584 40928 1636 40934
rect 1584 40870 1636 40876
rect 1306 40760 1362 40769
rect 1306 40695 1362 40704
rect 1308 38344 1360 38350
rect 1306 38312 1308 38321
rect 1360 38312 1362 38321
rect 1306 38247 1362 38256
rect 1308 33516 1360 33522
rect 1308 33458 1360 33464
rect 1320 33425 1348 33458
rect 1306 33416 1362 33425
rect 1306 33351 1362 33360
rect 1308 31272 1360 31278
rect 1308 31214 1360 31220
rect 1320 30977 1348 31214
rect 1306 30968 1362 30977
rect 1306 30903 1362 30912
rect 1596 30802 1624 40870
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 1768 36168 1820 36174
rect 1768 36110 1820 36116
rect 1780 35873 1808 36110
rect 3424 36032 3476 36038
rect 3424 35974 3476 35980
rect 1766 35864 1822 35873
rect 1766 35799 1822 35808
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 1952 31340 2004 31346
rect 1952 31282 2004 31288
rect 1584 30796 1636 30802
rect 1584 30738 1636 30744
rect 1308 28620 1360 28626
rect 1308 28562 1360 28568
rect 1320 28529 1348 28562
rect 1768 28552 1820 28558
rect 1306 28520 1362 28529
rect 1768 28494 1820 28500
rect 1306 28455 1362 28464
rect 1780 26042 1808 28494
rect 1964 28218 1992 31282
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 3436 28626 3464 35974
rect 3516 33312 3568 33318
rect 3516 33254 3568 33260
rect 3424 28620 3476 28626
rect 3424 28562 3476 28568
rect 1952 28212 2004 28218
rect 1952 28154 2004 28160
rect 3424 28076 3476 28082
rect 3424 28018 3476 28024
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2044 26376 2096 26382
rect 2044 26318 2096 26324
rect 1768 26036 1820 26042
rect 1768 25978 1820 25984
rect 1860 24064 1912 24070
rect 1860 24006 1912 24012
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1308 23656 1360 23662
rect 1306 23624 1308 23633
rect 1360 23624 1362 23633
rect 1306 23559 1362 23568
rect 1780 22778 1808 23666
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 1872 21554 1900 24006
rect 2056 23322 2084 26318
rect 2780 26308 2832 26314
rect 2780 26250 2832 26256
rect 2792 26081 2820 26250
rect 2778 26072 2834 26081
rect 2778 26007 2834 26016
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 2780 25832 2832 25838
rect 2780 25774 2832 25780
rect 2792 24206 2820 25774
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2884 23322 2912 25842
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 3344 24410 3372 26930
rect 3436 25770 3464 28018
rect 3528 26994 3556 33254
rect 3792 30660 3844 30666
rect 3792 30602 3844 30608
rect 3804 28218 3832 30602
rect 3884 29572 3936 29578
rect 3884 29514 3936 29520
rect 3792 28212 3844 28218
rect 3792 28154 3844 28160
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 3516 25968 3568 25974
rect 3516 25910 3568 25916
rect 3424 25764 3476 25770
rect 3424 25706 3476 25712
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2044 23316 2096 23322
rect 2044 23258 2096 23264
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 3344 23186 3372 24346
rect 3528 24206 3556 25910
rect 3620 25838 3648 28018
rect 3896 27130 3924 29514
rect 3988 28642 4016 43114
rect 4172 42294 4200 50866
rect 4264 50862 4292 52958
rect 4540 50998 4568 54130
rect 4344 50992 4396 50998
rect 4344 50934 4396 50940
rect 4528 50992 4580 50998
rect 4528 50934 4580 50940
rect 4252 50856 4304 50862
rect 4252 50798 4304 50804
rect 4356 42362 4384 50934
rect 4632 43382 4660 54130
rect 4712 52012 4764 52018
rect 4712 51954 4764 51960
rect 4724 43994 4752 51954
rect 4816 51950 4844 56200
rect 5184 53258 5212 56200
rect 5552 53718 5580 56200
rect 5920 54126 5948 56200
rect 5908 54120 5960 54126
rect 5908 54062 5960 54068
rect 5540 53712 5592 53718
rect 5540 53654 5592 53660
rect 5184 53230 5580 53258
rect 5172 52488 5224 52494
rect 5172 52430 5224 52436
rect 4896 52080 4948 52086
rect 4896 52022 4948 52028
rect 4804 51944 4856 51950
rect 4804 51886 4856 51892
rect 4712 43988 4764 43994
rect 4712 43930 4764 43936
rect 4620 43376 4672 43382
rect 4620 43318 4672 43324
rect 4908 42770 4936 52022
rect 5080 50176 5132 50182
rect 5080 50118 5132 50124
rect 4896 42764 4948 42770
rect 4896 42706 4948 42712
rect 5092 42362 5120 50118
rect 4344 42356 4396 42362
rect 4344 42298 4396 42304
rect 5080 42356 5132 42362
rect 5080 42298 5132 42304
rect 4160 42288 4212 42294
rect 4160 42230 4212 42236
rect 4252 42220 4304 42226
rect 4252 42162 4304 42168
rect 4068 38208 4120 38214
rect 4068 38150 4120 38156
rect 4080 29714 4108 38150
rect 4264 29850 4292 42162
rect 5184 41818 5212 52430
rect 5552 51474 5580 53230
rect 6288 53174 6316 56200
rect 6276 53168 6328 53174
rect 6276 53110 6328 53116
rect 6368 53100 6420 53106
rect 6368 53042 6420 53048
rect 5632 53032 5684 53038
rect 5632 52974 5684 52980
rect 5644 52154 5672 52974
rect 5724 52488 5776 52494
rect 5724 52430 5776 52436
rect 5632 52148 5684 52154
rect 5632 52090 5684 52096
rect 5540 51468 5592 51474
rect 5540 51410 5592 51416
rect 5540 51332 5592 51338
rect 5540 51274 5592 51280
rect 5552 51066 5580 51274
rect 5540 51060 5592 51066
rect 5540 51002 5592 51008
rect 5736 46170 5764 52430
rect 5816 50312 5868 50318
rect 5816 50254 5868 50260
rect 5724 46164 5776 46170
rect 5724 46106 5776 46112
rect 5828 44538 5856 50254
rect 6380 45082 6408 53042
rect 6656 52494 6684 56200
rect 6828 53576 6880 53582
rect 6828 53518 6880 53524
rect 6644 52488 6696 52494
rect 6644 52430 6696 52436
rect 6736 51400 6788 51406
rect 6736 51342 6788 51348
rect 6368 45076 6420 45082
rect 6368 45018 6420 45024
rect 6460 44736 6512 44742
rect 6460 44678 6512 44684
rect 5816 44532 5868 44538
rect 5816 44474 5868 44480
rect 6472 44402 6500 44678
rect 6748 44538 6776 51342
rect 6840 50522 6868 53518
rect 7024 51474 7052 56200
rect 7392 53650 7420 56200
rect 7380 53644 7432 53650
rect 7380 53586 7432 53592
rect 7380 53508 7432 53514
rect 7380 53450 7432 53456
rect 7288 52488 7340 52494
rect 7288 52430 7340 52436
rect 7012 51468 7064 51474
rect 7012 51410 7064 51416
rect 7104 51400 7156 51406
rect 7104 51342 7156 51348
rect 6828 50516 6880 50522
rect 6828 50458 6880 50464
rect 6736 44532 6788 44538
rect 6736 44474 6788 44480
rect 7116 44470 7144 51342
rect 7300 45014 7328 52430
rect 7392 46594 7420 53450
rect 7760 52562 7788 56200
rect 7852 54262 7880 56222
rect 8036 56114 8064 56222
rect 8114 56200 8170 57000
rect 8482 56200 8538 57000
rect 8850 56200 8906 57000
rect 9218 56200 9274 57000
rect 9586 56200 9642 57000
rect 9954 56200 10010 57000
rect 10322 56200 10378 57000
rect 10690 56200 10746 57000
rect 11058 56200 11114 57000
rect 11426 56200 11482 57000
rect 11794 56200 11850 57000
rect 12162 56200 12218 57000
rect 12530 56200 12586 57000
rect 12898 56200 12954 57000
rect 13266 56200 13322 57000
rect 13634 56200 13690 57000
rect 14002 56200 14058 57000
rect 14370 56200 14426 57000
rect 14738 56200 14794 57000
rect 15106 56200 15162 57000
rect 15474 56200 15530 57000
rect 15842 56200 15898 57000
rect 16210 56200 16266 57000
rect 16578 56200 16634 57000
rect 16946 56200 17002 57000
rect 17314 56200 17370 57000
rect 17682 56200 17738 57000
rect 18050 56200 18106 57000
rect 18156 56222 18368 56250
rect 8128 56114 8156 56200
rect 8036 56086 8156 56114
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 7840 54256 7892 54262
rect 7840 54198 7892 54204
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7748 52556 7800 52562
rect 7748 52498 7800 52504
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 8496 51950 8524 56200
rect 8864 53650 8892 56200
rect 8852 53644 8904 53650
rect 8852 53586 8904 53592
rect 9128 53576 9180 53582
rect 9128 53518 9180 53524
rect 8944 52488 8996 52494
rect 8944 52430 8996 52436
rect 8484 51944 8536 51950
rect 8484 51886 8536 51892
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7656 50924 7708 50930
rect 7656 50866 7708 50872
rect 7840 50924 7892 50930
rect 7840 50866 7892 50872
rect 7472 50856 7524 50862
rect 7472 50798 7524 50804
rect 7484 46714 7512 50798
rect 7564 50244 7616 50250
rect 7564 50186 7616 50192
rect 7472 46708 7524 46714
rect 7472 46650 7524 46656
rect 7392 46566 7512 46594
rect 7380 45892 7432 45898
rect 7380 45834 7432 45840
rect 7288 45008 7340 45014
rect 7288 44950 7340 44956
rect 7392 44826 7420 45834
rect 7300 44798 7420 44826
rect 7104 44464 7156 44470
rect 7104 44406 7156 44412
rect 5356 44396 5408 44402
rect 5356 44338 5408 44344
rect 6460 44396 6512 44402
rect 6460 44338 6512 44344
rect 5264 42560 5316 42566
rect 5264 42502 5316 42508
rect 5172 41812 5224 41818
rect 5172 41754 5224 41760
rect 4620 41132 4672 41138
rect 4620 41074 4672 41080
rect 4632 32570 4660 41074
rect 4988 37868 5040 37874
rect 4988 37810 5040 37816
rect 5000 32570 5028 37810
rect 5276 34474 5304 42502
rect 5368 38010 5396 44338
rect 6276 42016 6328 42022
rect 6276 41958 6328 41964
rect 6184 41676 6236 41682
rect 6184 41618 6236 41624
rect 5724 41472 5776 41478
rect 5724 41414 5776 41420
rect 5356 38004 5408 38010
rect 5356 37946 5408 37952
rect 5540 36916 5592 36922
rect 5540 36858 5592 36864
rect 5448 36712 5500 36718
rect 5448 36654 5500 36660
rect 5264 34468 5316 34474
rect 5264 34410 5316 34416
rect 5356 33448 5408 33454
rect 5356 33390 5408 33396
rect 5368 32570 5396 33390
rect 4620 32564 4672 32570
rect 4620 32506 4672 32512
rect 4988 32564 5040 32570
rect 4988 32506 5040 32512
rect 5356 32564 5408 32570
rect 5356 32506 5408 32512
rect 4896 32496 4948 32502
rect 4896 32438 4948 32444
rect 4252 29844 4304 29850
rect 4252 29786 4304 29792
rect 4068 29708 4120 29714
rect 4068 29650 4120 29656
rect 3988 28614 4108 28642
rect 3976 28484 4028 28490
rect 3976 28426 4028 28432
rect 3884 27124 3936 27130
rect 3884 27066 3936 27072
rect 3884 26784 3936 26790
rect 3884 26726 3936 26732
rect 3608 25832 3660 25838
rect 3608 25774 3660 25780
rect 3516 24200 3568 24206
rect 3516 24142 3568 24148
rect 2872 23180 2924 23186
rect 2872 23122 2924 23128
rect 3332 23180 3384 23186
rect 3332 23122 3384 23128
rect 2884 23066 2912 23122
rect 2792 23038 2912 23066
rect 3792 23044 3844 23050
rect 1860 21548 1912 21554
rect 1860 21490 1912 21496
rect 1308 21480 1360 21486
rect 1308 21422 1360 21428
rect 1320 21185 1348 21422
rect 1306 21176 1362 21185
rect 1306 21111 1362 21120
rect 2792 20806 2820 23038
rect 3792 22986 3844 22992
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2884 21146 2912 22578
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 1768 20800 1820 20806
rect 1768 20742 1820 20748
rect 2780 20800 2832 20806
rect 2780 20742 2832 20748
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 1308 18828 1360 18834
rect 1308 18770 1360 18776
rect 1320 18737 1348 18770
rect 1306 18728 1362 18737
rect 1306 18663 1362 18672
rect 1504 16590 1532 19450
rect 1780 18766 1808 20742
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3620 19378 3648 21422
rect 3804 21418 3832 22986
rect 3792 21412 3844 21418
rect 3792 21354 3844 21360
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 4080 16998 4108 20878
rect 4264 20534 4292 23174
rect 4356 21554 4384 25230
rect 4528 24132 4580 24138
rect 4528 24074 4580 24080
rect 4540 22094 4568 24074
rect 4540 22066 4660 22094
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 4356 20806 4384 21490
rect 4344 20800 4396 20806
rect 4344 20742 4396 20748
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4172 17338 4200 18702
rect 4356 17882 4384 20742
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 1492 16584 1544 16590
rect 1492 16526 1544 16532
rect 2502 16552 2558 16561
rect 1308 16516 1360 16522
rect 2502 16487 2558 16496
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 2516 16182 2544 16487
rect 2504 16176 2556 16182
rect 2504 16118 2556 16124
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 13938 1808 15846
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1308 13864 1360 13870
rect 1306 13832 1308 13841
rect 1360 13832 1362 13841
rect 1306 13767 1362 13776
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1504 2446 1532 2790
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 1688 800 1716 3470
rect 1872 2650 1900 13874
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2056 3058 2084 3334
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 2056 800 2084 2994
rect 2608 2650 2636 5646
rect 2700 3194 2728 15098
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2884 8809 2912 9590
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3068 8945 3096 9114
rect 3054 8936 3110 8945
rect 3054 8871 3110 8880
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2792 4010 2820 7754
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3068 6497 3096 6666
rect 3054 6488 3110 6497
rect 3054 6423 3110 6432
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 3148 4072 3200 4078
rect 3146 4040 3148 4049
rect 3200 4040 3202 4049
rect 2780 4004 2832 4010
rect 3146 3975 3202 3984
rect 2780 3946 2832 3952
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2792 3058 2820 3334
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2320 2440 2372 2446
rect 2372 2400 2452 2428
rect 2320 2382 2372 2388
rect 2424 800 2452 2400
rect 2792 800 2820 2994
rect 2884 1601 2912 3878
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3344 2990 3372 3402
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3436 2938 3464 3334
rect 3528 3058 3556 12038
rect 3896 11665 3924 26726
rect 3988 25158 4016 28426
rect 4080 26586 4108 28614
rect 4344 26920 4396 26926
rect 4344 26862 4396 26868
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 4080 25974 4108 26522
rect 4068 25968 4120 25974
rect 4068 25910 4120 25916
rect 4252 25696 4304 25702
rect 4252 25638 4304 25644
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3988 24206 4016 24550
rect 3976 24200 4028 24206
rect 3976 24142 4028 24148
rect 3988 23662 4016 24142
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 3988 21026 4016 23054
rect 4080 21486 4108 25230
rect 4264 24954 4292 25638
rect 4252 24948 4304 24954
rect 4252 24890 4304 24896
rect 4264 24274 4292 24890
rect 4252 24268 4304 24274
rect 4252 24210 4304 24216
rect 4356 23118 4384 26862
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4436 24404 4488 24410
rect 4436 24346 4488 24352
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 3988 20998 4108 21026
rect 4080 20942 4108 20998
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 4080 16561 4108 20878
rect 4172 19514 4200 21490
rect 4264 20942 4292 22374
rect 4448 22094 4476 24346
rect 4528 24132 4580 24138
rect 4528 24074 4580 24080
rect 4356 22066 4476 22094
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 4356 20534 4384 22066
rect 4540 21894 4568 24074
rect 4528 21888 4580 21894
rect 4528 21830 4580 21836
rect 4540 21554 4568 21830
rect 4528 21548 4580 21554
rect 4528 21490 4580 21496
rect 4344 20528 4396 20534
rect 4344 20470 4396 20476
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4066 16552 4122 16561
rect 4066 16487 4122 16496
rect 3882 11656 3938 11665
rect 3882 11591 3938 11600
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 3344 2632 3372 2926
rect 3436 2910 3556 2938
rect 3160 2604 3372 2632
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 3160 800 3188 2604
rect 3528 2378 3556 2910
rect 3896 2446 3924 3334
rect 4172 2650 4200 18022
rect 4540 17338 4568 21490
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4816 12434 4844 25842
rect 4908 18154 4936 32438
rect 5460 32366 5488 36654
rect 5552 35834 5580 36858
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 5552 35154 5580 35770
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 5552 34066 5580 35090
rect 5632 34468 5684 34474
rect 5632 34410 5684 34416
rect 5540 34060 5592 34066
rect 5540 34002 5592 34008
rect 5552 32978 5580 34002
rect 5540 32972 5592 32978
rect 5540 32914 5592 32920
rect 5552 32502 5580 32914
rect 5540 32496 5592 32502
rect 5540 32438 5592 32444
rect 5448 32360 5500 32366
rect 5448 32302 5500 32308
rect 5644 31278 5672 34410
rect 5736 31686 5764 41414
rect 6196 40526 6224 41618
rect 6288 41414 6316 41958
rect 6472 41414 6500 44338
rect 6920 43308 6972 43314
rect 6920 43250 6972 43256
rect 6736 42220 6788 42226
rect 6736 42162 6788 42168
rect 6748 41682 6776 42162
rect 6736 41676 6788 41682
rect 6736 41618 6788 41624
rect 6288 41386 6408 41414
rect 6472 41386 6684 41414
rect 6184 40520 6236 40526
rect 6184 40462 6236 40468
rect 6196 39506 6224 40462
rect 6184 39500 6236 39506
rect 6184 39442 6236 39448
rect 5816 39296 5868 39302
rect 5816 39238 5868 39244
rect 5828 37806 5856 39238
rect 5816 37800 5868 37806
rect 5816 37742 5868 37748
rect 5828 36718 5856 37742
rect 5816 36712 5868 36718
rect 5816 36654 5868 36660
rect 6000 36712 6052 36718
rect 6000 36654 6052 36660
rect 6012 35834 6040 36654
rect 6000 35828 6052 35834
rect 6000 35770 6052 35776
rect 5816 35624 5868 35630
rect 5816 35566 5868 35572
rect 5828 34066 5856 35566
rect 6012 34678 6040 35770
rect 6092 35148 6144 35154
rect 6092 35090 6144 35096
rect 6000 34672 6052 34678
rect 6000 34614 6052 34620
rect 6104 34610 6132 35090
rect 6092 34604 6144 34610
rect 6092 34546 6144 34552
rect 5816 34060 5868 34066
rect 5816 34002 5868 34008
rect 6184 32428 6236 32434
rect 6184 32370 6236 32376
rect 6196 31890 6224 32370
rect 6184 31884 6236 31890
rect 6184 31826 6236 31832
rect 5724 31680 5776 31686
rect 5724 31622 5776 31628
rect 5632 31272 5684 31278
rect 5632 31214 5684 31220
rect 6276 30660 6328 30666
rect 6276 30602 6328 30608
rect 6092 29572 6144 29578
rect 6092 29514 6144 29520
rect 5908 28620 5960 28626
rect 5908 28562 5960 28568
rect 5920 28218 5948 28562
rect 5908 28212 5960 28218
rect 5908 28154 5960 28160
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 4988 24812 5040 24818
rect 4988 24754 5040 24760
rect 5000 24274 5028 24754
rect 4988 24268 5040 24274
rect 4988 24210 5040 24216
rect 5000 24138 5028 24210
rect 4988 24132 5040 24138
rect 4988 24074 5040 24080
rect 5080 23044 5132 23050
rect 5080 22986 5132 22992
rect 5092 20058 5120 22986
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5080 20052 5132 20058
rect 5080 19994 5132 20000
rect 4896 18148 4948 18154
rect 4896 18090 4948 18096
rect 4724 12406 4844 12434
rect 4724 6914 4752 12406
rect 4724 6886 4844 6914
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4264 2446 4292 2790
rect 4816 2582 4844 6886
rect 4908 2922 4936 18090
rect 5460 13938 5488 20742
rect 5552 18086 5580 25094
rect 5724 23520 5776 23526
rect 5724 23462 5776 23468
rect 5736 23186 5764 23462
rect 5724 23180 5776 23186
rect 5724 23122 5776 23128
rect 5736 20398 5764 23122
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5736 20058 5764 20334
rect 5828 20262 5856 21286
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5828 13530 5856 20198
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 3516 2372 3568 2378
rect 3516 2314 3568 2320
rect 3528 800 3556 2314
rect 3896 800 3924 2382
rect 4264 800 4292 2382
rect 4632 800 4660 2382
rect 5000 800 5028 3334
rect 5184 3194 5212 11766
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5276 3738 5304 10406
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5552 3670 5580 9454
rect 5920 9178 5948 28154
rect 6000 24744 6052 24750
rect 6000 24686 6052 24692
rect 6012 23866 6040 24686
rect 6104 24342 6132 29514
rect 6184 25832 6236 25838
rect 6184 25774 6236 25780
rect 6196 24410 6224 25774
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6092 24336 6144 24342
rect 6092 24278 6144 24284
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 6012 22574 6040 23802
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 6104 22094 6132 24278
rect 6288 22438 6316 30602
rect 6380 29782 6408 41386
rect 6552 40588 6604 40594
rect 6552 40530 6604 40536
rect 6564 39642 6592 40530
rect 6552 39636 6604 39642
rect 6552 39578 6604 39584
rect 6460 38412 6512 38418
rect 6512 38372 6592 38400
rect 6460 38354 6512 38360
rect 6564 37806 6592 38372
rect 6552 37800 6604 37806
rect 6552 37742 6604 37748
rect 6564 37262 6592 37742
rect 6656 37670 6684 41386
rect 6932 40610 6960 43250
rect 7196 42016 7248 42022
rect 7196 41958 7248 41964
rect 7012 41472 7064 41478
rect 7012 41414 7064 41420
rect 7024 41386 7144 41414
rect 6932 40582 7052 40610
rect 6736 39568 6788 39574
rect 6736 39510 6788 39516
rect 6644 37664 6696 37670
rect 6644 37606 6696 37612
rect 6552 37256 6604 37262
rect 6552 37198 6604 37204
rect 6564 36922 6592 37198
rect 6552 36916 6604 36922
rect 6552 36858 6604 36864
rect 6368 29776 6420 29782
rect 6368 29718 6420 29724
rect 6552 29096 6604 29102
rect 6552 29038 6604 29044
rect 6564 28626 6592 29038
rect 6552 28620 6604 28626
rect 6552 28562 6604 28568
rect 6564 27538 6592 28562
rect 6552 27532 6604 27538
rect 6552 27474 6604 27480
rect 6564 26994 6592 27474
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 6564 26466 6592 26930
rect 6472 26450 6592 26466
rect 6460 26444 6592 26450
rect 6512 26438 6592 26444
rect 6460 26386 6512 26392
rect 6472 23186 6500 26386
rect 6460 23180 6512 23186
rect 6460 23122 6512 23128
rect 6276 22432 6328 22438
rect 6276 22374 6328 22380
rect 6288 22094 6316 22374
rect 6012 22066 6132 22094
rect 6196 22066 6316 22094
rect 6012 12434 6040 22066
rect 6012 12406 6132 12434
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 6104 6914 6132 12406
rect 6012 6886 6132 6914
rect 6012 6730 6040 6886
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 5906 6352 5962 6361
rect 5906 6287 5962 6296
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5920 3194 5948 6287
rect 6196 4078 6224 22066
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6564 20466 6592 20538
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6564 20058 6592 20402
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6288 17882 6316 19314
rect 6564 18766 6592 19314
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6564 17202 6592 18702
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6368 16652 6420 16658
rect 6564 16640 6592 17138
rect 6420 16612 6592 16640
rect 6368 16594 6420 16600
rect 6564 16114 6592 16612
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6564 13394 6592 16050
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6472 8090 6500 13126
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6564 9450 6592 12786
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6472 7886 6500 8026
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6104 3534 6132 3878
rect 6748 3738 6776 39510
rect 6920 38412 6972 38418
rect 6920 38354 6972 38360
rect 6932 37942 6960 38354
rect 6920 37936 6972 37942
rect 6920 37878 6972 37884
rect 6920 36848 6972 36854
rect 6920 36790 6972 36796
rect 6932 35834 6960 36790
rect 7024 36378 7052 40582
rect 7116 40390 7144 41386
rect 7104 40384 7156 40390
rect 7104 40326 7156 40332
rect 7012 36372 7064 36378
rect 7012 36314 7064 36320
rect 6920 35828 6972 35834
rect 6920 35770 6972 35776
rect 6932 35018 6960 35770
rect 7102 35728 7158 35737
rect 7102 35663 7158 35672
rect 6920 35012 6972 35018
rect 6920 34954 6972 34960
rect 6932 34678 6960 34954
rect 6920 34672 6972 34678
rect 6920 34614 6972 34620
rect 6920 34536 6972 34542
rect 6920 34478 6972 34484
rect 6932 31890 6960 34478
rect 6920 31884 6972 31890
rect 6920 31826 6972 31832
rect 6932 29714 6960 31826
rect 6920 29708 6972 29714
rect 6920 29650 6972 29656
rect 7116 29578 7144 35663
rect 7208 33318 7236 41958
rect 7300 38321 7328 44798
rect 7380 44736 7432 44742
rect 7380 44678 7432 44684
rect 7392 44402 7420 44678
rect 7484 44538 7512 46566
rect 7472 44532 7524 44538
rect 7472 44474 7524 44480
rect 7380 44396 7432 44402
rect 7380 44338 7432 44344
rect 7472 44396 7524 44402
rect 7472 44338 7524 44344
rect 7380 39296 7432 39302
rect 7380 39238 7432 39244
rect 7392 39098 7420 39238
rect 7380 39092 7432 39098
rect 7380 39034 7432 39040
rect 7392 38350 7420 39034
rect 7380 38344 7432 38350
rect 7286 38312 7342 38321
rect 7380 38286 7432 38292
rect 7286 38247 7342 38256
rect 7392 37942 7420 38286
rect 7380 37936 7432 37942
rect 7380 37878 7432 37884
rect 7392 37194 7420 37878
rect 7380 37188 7432 37194
rect 7380 37130 7432 37136
rect 7392 36854 7420 37130
rect 7484 36922 7512 44338
rect 7576 42106 7604 50186
rect 7668 46102 7696 50866
rect 7748 49836 7800 49842
rect 7748 49778 7800 49784
rect 7656 46096 7708 46102
rect 7656 46038 7708 46044
rect 7760 43450 7788 49778
rect 7852 44538 7880 50866
rect 8392 50312 8444 50318
rect 8392 50254 8444 50260
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 8300 48068 8352 48074
rect 8300 48010 8352 48016
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 7840 44532 7892 44538
rect 7840 44474 7892 44480
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 7748 43444 7800 43450
rect 7748 43386 7800 43392
rect 8312 42566 8340 48010
rect 8404 43994 8432 50254
rect 8852 49768 8904 49774
rect 8852 49710 8904 49716
rect 8668 45960 8720 45966
rect 8668 45902 8720 45908
rect 8576 44804 8628 44810
rect 8576 44746 8628 44752
rect 8392 43988 8444 43994
rect 8392 43930 8444 43936
rect 8484 43308 8536 43314
rect 8484 43250 8536 43256
rect 8496 42906 8524 43250
rect 8484 42900 8536 42906
rect 8484 42842 8536 42848
rect 8300 42560 8352 42566
rect 8496 42537 8524 42842
rect 8300 42502 8352 42508
rect 8482 42528 8538 42537
rect 7950 42460 8258 42469
rect 8482 42463 8538 42472
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 8484 42356 8536 42362
rect 8484 42298 8536 42304
rect 7748 42152 7800 42158
rect 7576 42078 7696 42106
rect 7748 42094 7800 42100
rect 7564 42016 7616 42022
rect 7564 41958 7616 41964
rect 7576 38554 7604 41958
rect 7668 40497 7696 42078
rect 7760 41818 7788 42094
rect 7748 41812 7800 41818
rect 7748 41754 7800 41760
rect 8300 41812 8352 41818
rect 8300 41754 8352 41760
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 8312 40730 8340 41754
rect 8300 40724 8352 40730
rect 8300 40666 8352 40672
rect 7654 40488 7710 40497
rect 8312 40458 8340 40666
rect 7654 40423 7710 40432
rect 8300 40452 8352 40458
rect 8300 40394 8352 40400
rect 7748 40384 7800 40390
rect 7668 40332 7748 40338
rect 7668 40326 7800 40332
rect 7668 40310 7788 40326
rect 7564 38548 7616 38554
rect 7564 38490 7616 38496
rect 7668 38486 7696 40310
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 8496 40050 8524 42298
rect 8484 40044 8536 40050
rect 8484 39986 8536 39992
rect 7748 39976 7800 39982
rect 7748 39918 7800 39924
rect 7840 39976 7892 39982
rect 7840 39918 7892 39924
rect 7760 39642 7788 39918
rect 7748 39636 7800 39642
rect 7748 39578 7800 39584
rect 7656 38480 7708 38486
rect 7656 38422 7708 38428
rect 7852 38418 7880 39918
rect 8588 39574 8616 44746
rect 8680 40186 8708 45902
rect 8760 45552 8812 45558
rect 8760 45494 8812 45500
rect 8772 45286 8800 45494
rect 8760 45280 8812 45286
rect 8760 45222 8812 45228
rect 8772 43314 8800 45222
rect 8760 43308 8812 43314
rect 8760 43250 8812 43256
rect 8864 42634 8892 49710
rect 8956 43450 8984 52430
rect 9036 52080 9088 52086
rect 9036 52022 9088 52028
rect 9048 47802 9076 52022
rect 9140 50522 9168 53518
rect 9232 53174 9260 56200
rect 9600 53564 9628 56200
rect 9968 54330 9996 56200
rect 9956 54324 10008 54330
rect 9956 54266 10008 54272
rect 9956 54188 10008 54194
rect 9956 54130 10008 54136
rect 9600 53536 9904 53564
rect 9220 53168 9272 53174
rect 9220 53110 9272 53116
rect 9680 53100 9732 53106
rect 9680 53042 9732 53048
rect 9220 51400 9272 51406
rect 9220 51342 9272 51348
rect 9128 50516 9180 50522
rect 9128 50458 9180 50464
rect 9036 47796 9088 47802
rect 9036 47738 9088 47744
rect 9232 46170 9260 51342
rect 9692 49910 9720 53042
rect 9772 52012 9824 52018
rect 9772 51954 9824 51960
rect 9680 49904 9732 49910
rect 9680 49846 9732 49852
rect 9496 49836 9548 49842
rect 9496 49778 9548 49784
rect 9312 46572 9364 46578
rect 9312 46514 9364 46520
rect 9220 46164 9272 46170
rect 9220 46106 9272 46112
rect 9220 46028 9272 46034
rect 9220 45970 9272 45976
rect 9036 43784 9088 43790
rect 9036 43726 9088 43732
rect 9128 43784 9180 43790
rect 9128 43726 9180 43732
rect 8944 43444 8996 43450
rect 8944 43386 8996 43392
rect 8944 43308 8996 43314
rect 8944 43250 8996 43256
rect 8956 42906 8984 43250
rect 8944 42900 8996 42906
rect 8944 42842 8996 42848
rect 8852 42628 8904 42634
rect 8852 42570 8904 42576
rect 8760 42560 8812 42566
rect 8760 42502 8812 42508
rect 8772 41414 8800 42502
rect 8864 42226 8892 42570
rect 8956 42566 8984 42842
rect 8944 42560 8996 42566
rect 8944 42502 8996 42508
rect 8852 42220 8904 42226
rect 8852 42162 8904 42168
rect 8864 41818 8892 42162
rect 8852 41812 8904 41818
rect 8852 41754 8904 41760
rect 8772 41386 8892 41414
rect 8668 40180 8720 40186
rect 8668 40122 8720 40128
rect 8760 40112 8812 40118
rect 8760 40054 8812 40060
rect 8576 39568 8628 39574
rect 8628 39528 8708 39556
rect 8576 39510 8628 39516
rect 8576 39432 8628 39438
rect 8576 39374 8628 39380
rect 8300 39296 8352 39302
rect 8300 39238 8352 39244
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7840 38412 7892 38418
rect 7840 38354 7892 38360
rect 8312 38350 8340 39238
rect 8484 38820 8536 38826
rect 8484 38762 8536 38768
rect 8300 38344 8352 38350
rect 8206 38312 8262 38321
rect 8300 38286 8352 38292
rect 8206 38247 8262 38256
rect 8220 38214 8248 38247
rect 8208 38208 8260 38214
rect 8208 38150 8260 38156
rect 8392 38208 8444 38214
rect 8392 38150 8444 38156
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 7840 38004 7892 38010
rect 7840 37946 7892 37952
rect 7472 36916 7524 36922
rect 7472 36858 7524 36864
rect 7380 36848 7432 36854
rect 7380 36790 7432 36796
rect 7656 36644 7708 36650
rect 7656 36586 7708 36592
rect 7472 36236 7524 36242
rect 7472 36178 7524 36184
rect 7288 34672 7340 34678
rect 7288 34614 7340 34620
rect 7300 34202 7328 34614
rect 7288 34196 7340 34202
rect 7288 34138 7340 34144
rect 7300 33930 7328 34138
rect 7288 33924 7340 33930
rect 7288 33866 7340 33872
rect 7300 33658 7328 33866
rect 7380 33856 7432 33862
rect 7380 33798 7432 33804
rect 7288 33652 7340 33658
rect 7288 33594 7340 33600
rect 7196 33312 7248 33318
rect 7196 33254 7248 33260
rect 7300 32910 7328 33594
rect 7288 32904 7340 32910
rect 7288 32846 7340 32852
rect 7300 32502 7328 32846
rect 7288 32496 7340 32502
rect 7288 32438 7340 32444
rect 7392 31210 7420 33798
rect 7484 32978 7512 36178
rect 7668 36174 7696 36586
rect 7852 36378 7880 37946
rect 8300 37324 8352 37330
rect 8300 37266 8352 37272
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 8312 36802 8340 37266
rect 8404 36922 8432 38150
rect 8496 37806 8524 38762
rect 8588 38282 8616 39374
rect 8680 39030 8708 39528
rect 8668 39024 8720 39030
rect 8668 38966 8720 38972
rect 8576 38276 8628 38282
rect 8576 38218 8628 38224
rect 8484 37800 8536 37806
rect 8484 37742 8536 37748
rect 8496 37398 8524 37742
rect 8588 37466 8616 38218
rect 8576 37460 8628 37466
rect 8576 37402 8628 37408
rect 8484 37392 8536 37398
rect 8484 37334 8536 37340
rect 8392 36916 8444 36922
rect 8392 36858 8444 36864
rect 8312 36774 8432 36802
rect 7840 36372 7892 36378
rect 7840 36314 7892 36320
rect 7656 36168 7708 36174
rect 7656 36110 7708 36116
rect 7668 35290 7696 36110
rect 7748 36032 7800 36038
rect 7748 35974 7800 35980
rect 7656 35284 7708 35290
rect 7656 35226 7708 35232
rect 7656 33924 7708 33930
rect 7656 33866 7708 33872
rect 7472 32972 7524 32978
rect 7472 32914 7524 32920
rect 7484 32366 7512 32914
rect 7472 32360 7524 32366
rect 7472 32302 7524 32308
rect 7668 31482 7696 33866
rect 7760 33114 7788 35974
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 8300 33380 8352 33386
rect 8300 33322 8352 33328
rect 7748 33108 7800 33114
rect 7748 33050 7800 33056
rect 8312 32978 8340 33322
rect 8300 32972 8352 32978
rect 8300 32914 8352 32920
rect 7748 32836 7800 32842
rect 7748 32778 7800 32784
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 7380 31204 7432 31210
rect 7380 31146 7432 31152
rect 7760 29850 7788 32778
rect 7840 32768 7892 32774
rect 7840 32710 7892 32716
rect 7852 32570 7880 32710
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 7840 32564 7892 32570
rect 7840 32506 7892 32512
rect 8312 32026 8340 32914
rect 8300 32020 8352 32026
rect 8300 31962 8352 31968
rect 8404 31958 8432 36774
rect 8496 33862 8524 37334
rect 8588 35222 8616 37402
rect 8668 36848 8720 36854
rect 8668 36790 8720 36796
rect 8680 35766 8708 36790
rect 8668 35760 8720 35766
rect 8668 35702 8720 35708
rect 8680 35290 8708 35702
rect 8772 35290 8800 40054
rect 8864 38894 8892 41386
rect 8852 38888 8904 38894
rect 8852 38830 8904 38836
rect 8956 38010 8984 42502
rect 8944 38004 8996 38010
rect 8944 37946 8996 37952
rect 9048 36922 9076 43726
rect 9140 42770 9168 43726
rect 9232 43246 9260 45970
rect 9220 43240 9272 43246
rect 9220 43182 9272 43188
rect 9128 42764 9180 42770
rect 9128 42706 9180 42712
rect 9140 41206 9168 42706
rect 9324 42022 9352 46514
rect 9508 45558 9536 49778
rect 9496 45552 9548 45558
rect 9496 45494 9548 45500
rect 9680 44736 9732 44742
rect 9680 44678 9732 44684
rect 9404 44396 9456 44402
rect 9404 44338 9456 44344
rect 9416 44305 9444 44338
rect 9402 44296 9458 44305
rect 9402 44231 9458 44240
rect 9496 43444 9548 43450
rect 9496 43386 9548 43392
rect 9220 42016 9272 42022
rect 9220 41958 9272 41964
rect 9312 42016 9364 42022
rect 9312 41958 9364 41964
rect 9232 41750 9260 41958
rect 9220 41744 9272 41750
rect 9220 41686 9272 41692
rect 9128 41200 9180 41206
rect 9128 41142 9180 41148
rect 9508 40730 9536 43386
rect 9588 43240 9640 43246
rect 9588 43182 9640 43188
rect 9496 40724 9548 40730
rect 9496 40666 9548 40672
rect 9404 40588 9456 40594
rect 9404 40530 9456 40536
rect 9220 40452 9272 40458
rect 9220 40394 9272 40400
rect 9232 40118 9260 40394
rect 9416 40390 9444 40530
rect 9404 40384 9456 40390
rect 9404 40326 9456 40332
rect 9220 40112 9272 40118
rect 9220 40054 9272 40060
rect 9232 39098 9260 40054
rect 9220 39092 9272 39098
rect 9220 39034 9272 39040
rect 9128 38752 9180 38758
rect 9128 38694 9180 38700
rect 9140 38418 9168 38694
rect 9128 38412 9180 38418
rect 9128 38354 9180 38360
rect 9220 38344 9272 38350
rect 9220 38286 9272 38292
rect 9036 36916 9088 36922
rect 9036 36858 9088 36864
rect 9128 36780 9180 36786
rect 9128 36722 9180 36728
rect 8852 35488 8904 35494
rect 8852 35430 8904 35436
rect 8668 35284 8720 35290
rect 8668 35226 8720 35232
rect 8760 35284 8812 35290
rect 8760 35226 8812 35232
rect 8576 35216 8628 35222
rect 8576 35158 8628 35164
rect 8680 35170 8708 35226
rect 8680 35142 8800 35170
rect 8668 35012 8720 35018
rect 8668 34954 8720 34960
rect 8484 33856 8536 33862
rect 8484 33798 8536 33804
rect 8484 32564 8536 32570
rect 8484 32506 8536 32512
rect 8392 31952 8444 31958
rect 8392 31894 8444 31900
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 8404 31414 8432 31894
rect 8496 31890 8524 32506
rect 8484 31884 8536 31890
rect 8484 31826 8536 31832
rect 8484 31680 8536 31686
rect 8484 31622 8536 31628
rect 8392 31408 8444 31414
rect 8392 31350 8444 31356
rect 7840 31340 7892 31346
rect 7840 31282 7892 31288
rect 7852 30802 7880 31282
rect 8496 31278 8524 31622
rect 8680 31482 8708 34954
rect 8772 34746 8800 35142
rect 8760 34740 8812 34746
rect 8760 34682 8812 34688
rect 8864 34610 8892 35430
rect 8852 34604 8904 34610
rect 8852 34546 8904 34552
rect 8864 33969 8892 34546
rect 9140 34202 9168 36722
rect 9128 34196 9180 34202
rect 9128 34138 9180 34144
rect 9232 34066 9260 38286
rect 9416 36922 9444 40326
rect 9508 39098 9536 40666
rect 9600 40594 9628 43182
rect 9692 42242 9720 44678
rect 9784 44538 9812 51954
rect 9876 51950 9904 53536
rect 9864 51944 9916 51950
rect 9864 51886 9916 51892
rect 9968 51610 9996 54130
rect 10336 53038 10364 56200
rect 10416 53576 10468 53582
rect 10416 53518 10468 53524
rect 10232 53032 10284 53038
rect 10232 52974 10284 52980
rect 10324 53032 10376 53038
rect 10324 52974 10376 52980
rect 10244 52850 10272 52974
rect 10244 52822 10364 52850
rect 10140 52080 10192 52086
rect 10140 52022 10192 52028
rect 9956 51604 10008 51610
rect 9956 51546 10008 51552
rect 9772 44532 9824 44538
rect 9772 44474 9824 44480
rect 10152 43450 10180 52022
rect 10232 49972 10284 49978
rect 10232 49914 10284 49920
rect 10244 47122 10272 49914
rect 10232 47116 10284 47122
rect 10232 47058 10284 47064
rect 10244 45286 10272 47058
rect 10232 45280 10284 45286
rect 10232 45222 10284 45228
rect 10140 43444 10192 43450
rect 10140 43386 10192 43392
rect 10244 42362 10272 45222
rect 10336 44470 10364 52822
rect 10428 44946 10456 53518
rect 10704 52562 10732 56200
rect 11072 53650 11100 56200
rect 11440 54262 11468 56200
rect 11428 54256 11480 54262
rect 11428 54198 11480 54204
rect 11244 54120 11296 54126
rect 11244 54062 11296 54068
rect 11060 53644 11112 53650
rect 11060 53586 11112 53592
rect 10692 52556 10744 52562
rect 10692 52498 10744 52504
rect 10784 52488 10836 52494
rect 10784 52430 10836 52436
rect 10796 50998 10824 52430
rect 10876 52012 10928 52018
rect 10876 51954 10928 51960
rect 10784 50992 10836 50998
rect 10784 50934 10836 50940
rect 10600 49224 10652 49230
rect 10600 49166 10652 49172
rect 10692 49224 10744 49230
rect 10692 49166 10744 49172
rect 10612 45554 10640 49166
rect 10704 46170 10732 49166
rect 10784 46980 10836 46986
rect 10784 46922 10836 46928
rect 10692 46164 10744 46170
rect 10692 46106 10744 46112
rect 10612 45526 10732 45554
rect 10416 44940 10468 44946
rect 10416 44882 10468 44888
rect 10324 44464 10376 44470
rect 10324 44406 10376 44412
rect 10600 44328 10652 44334
rect 10600 44270 10652 44276
rect 10324 43648 10376 43654
rect 10324 43590 10376 43596
rect 10232 42356 10284 42362
rect 10232 42298 10284 42304
rect 9692 42214 9812 42242
rect 9588 40588 9640 40594
rect 9588 40530 9640 40536
rect 9680 40588 9732 40594
rect 9680 40530 9732 40536
rect 9586 40488 9642 40497
rect 9586 40423 9588 40432
rect 9640 40423 9642 40432
rect 9588 40394 9640 40400
rect 9692 40338 9720 40530
rect 9600 40310 9720 40338
rect 9600 40186 9628 40310
rect 9588 40180 9640 40186
rect 9588 40122 9640 40128
rect 9496 39092 9548 39098
rect 9496 39034 9548 39040
rect 9600 38978 9628 40122
rect 9508 38950 9628 38978
rect 9508 37330 9536 38950
rect 9588 38888 9640 38894
rect 9586 38856 9588 38865
rect 9640 38856 9642 38865
rect 9586 38791 9642 38800
rect 9496 37324 9548 37330
rect 9496 37266 9548 37272
rect 9404 36916 9456 36922
rect 9404 36858 9456 36864
rect 9784 36825 9812 42214
rect 10140 42152 10192 42158
rect 10140 42094 10192 42100
rect 9956 40928 10008 40934
rect 9956 40870 10008 40876
rect 9968 39982 9996 40870
rect 9956 39976 10008 39982
rect 9956 39918 10008 39924
rect 10152 38486 10180 42094
rect 10244 41682 10272 42298
rect 10232 41676 10284 41682
rect 10232 41618 10284 41624
rect 10336 41614 10364 43590
rect 10416 43308 10468 43314
rect 10416 43250 10468 43256
rect 10428 42566 10456 43250
rect 10416 42560 10468 42566
rect 10414 42528 10416 42537
rect 10468 42528 10470 42537
rect 10414 42463 10470 42472
rect 10324 41608 10376 41614
rect 10324 41550 10376 41556
rect 10416 41540 10468 41546
rect 10416 41482 10468 41488
rect 10232 40656 10284 40662
rect 10232 40598 10284 40604
rect 10244 39506 10272 40598
rect 10232 39500 10284 39506
rect 10232 39442 10284 39448
rect 10140 38480 10192 38486
rect 10140 38422 10192 38428
rect 9956 37800 10008 37806
rect 9956 37742 10008 37748
rect 9968 37108 9996 37742
rect 10140 37664 10192 37670
rect 10140 37606 10192 37612
rect 9968 37080 10088 37108
rect 9770 36816 9826 36825
rect 9312 36780 9364 36786
rect 9770 36751 9826 36760
rect 9954 36816 10010 36825
rect 9954 36751 10010 36760
rect 9312 36722 9364 36728
rect 9220 34060 9272 34066
rect 9220 34002 9272 34008
rect 8850 33960 8906 33969
rect 8850 33895 8906 33904
rect 9324 33114 9352 36722
rect 9588 36712 9640 36718
rect 9588 36654 9640 36660
rect 9600 35630 9628 36654
rect 9588 35624 9640 35630
rect 9588 35566 9640 35572
rect 9600 34728 9628 35566
rect 9772 35488 9824 35494
rect 9772 35430 9824 35436
rect 9784 35154 9812 35430
rect 9772 35148 9824 35154
rect 9772 35090 9824 35096
rect 9772 34740 9824 34746
rect 9600 34700 9772 34728
rect 9772 34682 9824 34688
rect 9864 34400 9916 34406
rect 9864 34342 9916 34348
rect 9402 33960 9458 33969
rect 9402 33895 9458 33904
rect 9632 33930 9688 33935
rect 9632 33926 9732 33930
rect 9688 33924 9732 33926
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9416 31822 9444 33895
rect 9688 33870 9732 33872
rect 9632 33866 9732 33870
rect 9632 33861 9688 33866
rect 9772 33448 9824 33454
rect 9772 33390 9824 33396
rect 9680 33040 9732 33046
rect 9680 32982 9732 32988
rect 9496 32768 9548 32774
rect 9496 32710 9548 32716
rect 9404 31816 9456 31822
rect 9404 31758 9456 31764
rect 8668 31476 8720 31482
rect 8668 31418 8720 31424
rect 8944 31340 8996 31346
rect 8944 31282 8996 31288
rect 8116 31272 8168 31278
rect 8116 31214 8168 31220
rect 8484 31272 8536 31278
rect 8484 31214 8536 31220
rect 8128 30938 8156 31214
rect 8116 30932 8168 30938
rect 8116 30874 8168 30880
rect 7840 30796 7892 30802
rect 7840 30738 7892 30744
rect 8496 30598 8524 31214
rect 8484 30592 8536 30598
rect 8484 30534 8536 30540
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 8392 30320 8444 30326
rect 8392 30262 8444 30268
rect 7656 29844 7708 29850
rect 7656 29786 7708 29792
rect 7748 29844 7800 29850
rect 7748 29786 7800 29792
rect 7104 29572 7156 29578
rect 7104 29514 7156 29520
rect 7668 29510 7696 29786
rect 7840 29640 7892 29646
rect 7840 29582 7892 29588
rect 7380 29504 7432 29510
rect 7656 29504 7708 29510
rect 7380 29446 7432 29452
rect 7484 29452 7656 29458
rect 7484 29446 7708 29452
rect 7012 27532 7064 27538
rect 7012 27474 7064 27480
rect 7024 27402 7052 27474
rect 7012 27396 7064 27402
rect 7012 27338 7064 27344
rect 7024 27282 7052 27338
rect 7024 27254 7144 27282
rect 7116 27062 7144 27254
rect 7104 27056 7156 27062
rect 7104 26998 7156 27004
rect 7116 26246 7144 26998
rect 7104 26240 7156 26246
rect 7392 26194 7420 29446
rect 7104 26182 7156 26188
rect 7116 26042 7144 26182
rect 7208 26166 7420 26194
rect 7484 29430 7696 29446
rect 7104 26036 7156 26042
rect 7104 25978 7156 25984
rect 7116 25226 7144 25978
rect 7104 25220 7156 25226
rect 7104 25162 7156 25168
rect 7116 24886 7144 25162
rect 7104 24880 7156 24886
rect 7104 24822 7156 24828
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 6840 19310 6868 23802
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6932 21418 6960 22578
rect 7024 21690 7052 24142
rect 7104 23792 7156 23798
rect 7104 23734 7156 23740
rect 7116 23186 7144 23734
rect 7104 23180 7156 23186
rect 7104 23122 7156 23128
rect 7012 21684 7064 21690
rect 7012 21626 7064 21632
rect 6920 21412 6972 21418
rect 6920 21354 6972 21360
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7116 19854 7144 20470
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7116 19446 7144 19790
rect 7104 19440 7156 19446
rect 7104 19382 7156 19388
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6932 17134 6960 17682
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6932 16794 6960 17070
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 6840 7954 6868 13330
rect 7116 9518 7144 13330
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 7010 5672 7066 5681
rect 7010 5607 7066 5616
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5368 800 5396 2994
rect 5736 2378 5764 2994
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5736 800 5764 2314
rect 6104 800 6132 3470
rect 6472 2854 6500 3470
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 3058 6868 3334
rect 7024 3194 7052 5607
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6472 800 6500 2790
rect 6840 800 6868 2994
rect 7116 2650 7144 9318
rect 7208 3194 7236 26166
rect 7484 26058 7512 29430
rect 7656 29300 7708 29306
rect 7656 29242 7708 29248
rect 7668 26246 7696 29242
rect 7852 27606 7880 29582
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 7840 27600 7892 27606
rect 7840 27542 7892 27548
rect 7852 26926 7880 27542
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 7840 26920 7892 26926
rect 7760 26880 7840 26908
rect 7656 26240 7708 26246
rect 7656 26182 7708 26188
rect 7392 26030 7512 26058
rect 7392 24818 7420 26030
rect 7668 25498 7696 26182
rect 7472 25492 7524 25498
rect 7472 25434 7524 25440
rect 7656 25492 7708 25498
rect 7656 25434 7708 25440
rect 7484 24886 7512 25434
rect 7656 25356 7708 25362
rect 7656 25298 7708 25304
rect 7472 24880 7524 24886
rect 7472 24822 7524 24828
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7472 24608 7524 24614
rect 7472 24550 7524 24556
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7300 21146 7328 22510
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 17882 7328 19654
rect 7484 18426 7512 24550
rect 7668 23662 7696 25298
rect 7760 24818 7788 26880
rect 7840 26862 7892 26868
rect 8300 26852 8352 26858
rect 8300 26794 8352 26800
rect 8312 26450 8340 26794
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 7840 25832 7892 25838
rect 7840 25774 7892 25780
rect 8404 25786 8432 30262
rect 8496 25906 8524 30534
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 8680 28014 8708 28902
rect 8576 28008 8628 28014
rect 8576 27950 8628 27956
rect 8668 28008 8720 28014
rect 8668 27950 8720 27956
rect 8588 26586 8616 27950
rect 8956 26926 8984 31282
rect 9416 31278 9444 31758
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9416 30802 9444 31214
rect 9404 30796 9456 30802
rect 9404 30738 9456 30744
rect 9508 29850 9536 32710
rect 9692 32570 9720 32982
rect 9784 32910 9812 33390
rect 9876 32978 9904 34342
rect 9864 32972 9916 32978
rect 9864 32914 9916 32920
rect 9772 32904 9824 32910
rect 9772 32846 9824 32852
rect 9680 32564 9732 32570
rect 9680 32506 9732 32512
rect 9692 32026 9720 32506
rect 9864 32360 9916 32366
rect 9864 32302 9916 32308
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 9496 29844 9548 29850
rect 9496 29786 9548 29792
rect 9312 29776 9364 29782
rect 9312 29718 9364 29724
rect 9588 29776 9640 29782
rect 9588 29718 9640 29724
rect 9036 29232 9088 29238
rect 9036 29174 9088 29180
rect 9048 29034 9076 29174
rect 9036 29028 9088 29034
rect 9036 28970 9088 28976
rect 9048 28422 9076 28970
rect 9036 28416 9088 28422
rect 9036 28358 9088 28364
rect 9048 28150 9076 28358
rect 9036 28144 9088 28150
rect 9036 28086 9088 28092
rect 9048 27538 9076 28086
rect 9036 27532 9088 27538
rect 9036 27474 9088 27480
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 8944 26920 8996 26926
rect 8944 26862 8996 26868
rect 8576 26580 8628 26586
rect 8576 26522 8628 26528
rect 8484 25900 8536 25906
rect 8484 25842 8536 25848
rect 7852 24954 7880 25774
rect 8404 25758 8524 25786
rect 8588 25770 8616 26522
rect 8956 26314 8984 26862
rect 9140 26450 9168 26930
rect 9128 26444 9180 26450
rect 9128 26386 9180 26392
rect 8944 26308 8996 26314
rect 8944 26250 8996 26256
rect 8852 26036 8904 26042
rect 8852 25978 8904 25984
rect 8392 25220 8444 25226
rect 8392 25162 8444 25168
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7840 24948 7892 24954
rect 7840 24890 7892 24896
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 8116 24744 8168 24750
rect 8116 24686 8168 24692
rect 8128 24426 8156 24686
rect 8404 24682 8432 25162
rect 8392 24676 8444 24682
rect 8392 24618 8444 24624
rect 8128 24398 8432 24426
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8208 23792 8260 23798
rect 8312 23746 8340 24210
rect 8260 23740 8340 23746
rect 8208 23734 8340 23740
rect 8220 23718 8340 23734
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7576 23322 7604 23598
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7576 22574 7604 23258
rect 7656 23112 7708 23118
rect 7656 23054 7708 23060
rect 7564 22568 7616 22574
rect 7564 22510 7616 22516
rect 7576 22094 7604 22510
rect 7668 22420 7696 23054
rect 7748 23044 7800 23050
rect 7748 22986 7800 22992
rect 7760 22522 7788 22986
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7760 22494 7880 22522
rect 7668 22392 7788 22420
rect 7576 22066 7696 22094
rect 7668 21622 7696 22066
rect 7656 21616 7708 21622
rect 7656 21558 7708 21564
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7668 19786 7696 21422
rect 7760 19854 7788 22392
rect 7852 21010 7880 22494
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7840 21004 7892 21010
rect 7840 20946 7892 20952
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8312 19922 8340 20198
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 8208 19848 8260 19854
rect 8260 19796 8340 19802
rect 8208 19790 8340 19796
rect 7656 19780 7708 19786
rect 8220 19774 8340 19790
rect 7656 19722 7708 19728
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7576 18222 7604 19110
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7300 16250 7328 17478
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7484 16522 7512 16730
rect 7472 16516 7524 16522
rect 7472 16458 7524 16464
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7484 16182 7512 16458
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 7484 15706 7512 16118
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7576 13394 7604 18158
rect 7852 17746 7880 19450
rect 8312 18970 8340 19774
rect 8404 19378 8432 24398
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8312 17814 8340 18906
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7852 16522 7880 17478
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8312 17270 8340 17750
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 8312 16794 8340 17206
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8404 16726 8432 17682
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 7840 16516 7892 16522
rect 7840 16458 7892 16464
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8312 16046 8340 16594
rect 8404 16046 8432 16662
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8312 12986 8340 17478
rect 8496 16046 8524 19468
rect 8680 18834 8708 22510
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8588 18222 8616 18702
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8772 17320 8800 19178
rect 8680 17292 8800 17320
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8496 13530 8524 14010
rect 8588 13870 8616 14350
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8496 13258 8524 13466
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8496 12918 8524 13194
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8588 12782 8616 13126
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8680 12434 8708 17292
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8772 15910 8800 17138
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8864 15910 8892 16526
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8864 14822 8892 15846
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8864 14482 8892 14758
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8588 12406 8708 12434
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7760 2514 7788 8910
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8588 6914 8616 12406
rect 8864 12170 8892 12718
rect 8852 12164 8904 12170
rect 8852 12106 8904 12112
rect 8588 6886 8892 6914
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8220 3738 8248 4150
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7208 800 7236 2382
rect 7576 800 7604 2382
rect 7852 1986 7880 3334
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8208 3052 8260 3058
rect 8312 3040 8340 3538
rect 8496 3194 8524 25758
rect 8576 25764 8628 25770
rect 8576 25706 8628 25712
rect 8864 25498 8892 25978
rect 8852 25492 8904 25498
rect 8852 25434 8904 25440
rect 8576 25356 8628 25362
rect 8576 25298 8628 25304
rect 8588 24206 8616 25298
rect 8668 24404 8720 24410
rect 8668 24346 8720 24352
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8588 23662 8616 24142
rect 8576 23656 8628 23662
rect 8576 23598 8628 23604
rect 8680 20874 8708 24346
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8772 22778 8800 24006
rect 8760 22772 8812 22778
rect 8760 22714 8812 22720
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 8772 20330 8800 21422
rect 8864 20602 8892 22510
rect 8956 22094 8984 26250
rect 9324 24750 9352 29718
rect 9600 29578 9628 29718
rect 9692 29714 9720 31962
rect 9772 31680 9824 31686
rect 9772 31622 9824 31628
rect 9680 29708 9732 29714
rect 9680 29650 9732 29656
rect 9588 29572 9640 29578
rect 9588 29514 9640 29520
rect 9784 29306 9812 31622
rect 9876 31482 9904 32302
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 9968 29578 9996 36751
rect 10060 30190 10088 37080
rect 10152 36174 10180 37606
rect 10428 37466 10456 41482
rect 10612 41313 10640 44270
rect 10704 43654 10732 45526
rect 10796 45354 10824 46922
rect 10888 46714 10916 51954
rect 10876 46708 10928 46714
rect 10876 46650 10928 46656
rect 11060 46572 11112 46578
rect 11060 46514 11112 46520
rect 10968 45960 11020 45966
rect 10968 45902 11020 45908
rect 10876 45552 10928 45558
rect 10876 45494 10928 45500
rect 10784 45348 10836 45354
rect 10784 45290 10836 45296
rect 10888 45286 10916 45494
rect 10876 45280 10928 45286
rect 10876 45222 10928 45228
rect 10784 43716 10836 43722
rect 10888 43704 10916 45222
rect 10836 43676 10916 43704
rect 10784 43658 10836 43664
rect 10692 43648 10744 43654
rect 10692 43590 10744 43596
rect 10796 43110 10824 43658
rect 10784 43104 10836 43110
rect 10784 43046 10836 43052
rect 10876 42560 10928 42566
rect 10876 42502 10928 42508
rect 10784 42016 10836 42022
rect 10784 41958 10836 41964
rect 10692 41676 10744 41682
rect 10692 41618 10744 41624
rect 10598 41304 10654 41313
rect 10598 41239 10654 41248
rect 10704 40934 10732 41618
rect 10796 41546 10824 41958
rect 10888 41750 10916 42502
rect 10876 41744 10928 41750
rect 10876 41686 10928 41692
rect 10784 41540 10836 41546
rect 10784 41482 10836 41488
rect 10888 41426 10916 41686
rect 10796 41398 10916 41426
rect 10692 40928 10744 40934
rect 10692 40870 10744 40876
rect 10796 39846 10824 41398
rect 10876 41064 10928 41070
rect 10876 41006 10928 41012
rect 10784 39840 10836 39846
rect 10784 39782 10836 39788
rect 10796 38962 10824 39782
rect 10888 39642 10916 41006
rect 10980 40118 11008 45902
rect 11072 41818 11100 46514
rect 11152 45824 11204 45830
rect 11152 45766 11204 45772
rect 11164 44538 11192 45766
rect 11256 45082 11284 54062
rect 11704 53984 11756 53990
rect 11704 53926 11756 53932
rect 11716 49774 11744 53926
rect 11808 53038 11836 56200
rect 12176 53650 12204 56200
rect 12348 54188 12400 54194
rect 12348 54130 12400 54136
rect 12164 53644 12216 53650
rect 12164 53586 12216 53592
rect 11888 53100 11940 53106
rect 11888 53042 11940 53048
rect 11796 53032 11848 53038
rect 11796 52974 11848 52980
rect 11900 52154 11928 53042
rect 12360 52154 12388 54130
rect 12544 54126 12572 56200
rect 12912 54262 12940 56200
rect 13280 55214 13308 56200
rect 13280 55186 13400 55214
rect 12900 54256 12952 54262
rect 12900 54198 12952 54204
rect 12532 54120 12584 54126
rect 12532 54062 12584 54068
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12624 53576 12676 53582
rect 12624 53518 12676 53524
rect 12636 52698 12664 53518
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12624 52692 12676 52698
rect 12624 52634 12676 52640
rect 12808 52488 12860 52494
rect 12808 52430 12860 52436
rect 11888 52148 11940 52154
rect 11888 52090 11940 52096
rect 12348 52148 12400 52154
rect 12348 52090 12400 52096
rect 11980 52012 12032 52018
rect 11980 51954 12032 51960
rect 11704 49768 11756 49774
rect 11704 49710 11756 49716
rect 11992 49434 12020 51954
rect 12716 49768 12768 49774
rect 12716 49710 12768 49716
rect 11980 49428 12032 49434
rect 11980 49370 12032 49376
rect 12532 48748 12584 48754
rect 12532 48690 12584 48696
rect 11796 47660 11848 47666
rect 11796 47602 11848 47608
rect 11704 45892 11756 45898
rect 11704 45834 11756 45840
rect 11244 45076 11296 45082
rect 11244 45018 11296 45024
rect 11520 44804 11572 44810
rect 11520 44746 11572 44752
rect 11532 44577 11560 44746
rect 11518 44568 11574 44577
rect 11152 44532 11204 44538
rect 11518 44503 11574 44512
rect 11152 44474 11204 44480
rect 11612 44464 11664 44470
rect 11612 44406 11664 44412
rect 11520 44396 11572 44402
rect 11520 44338 11572 44344
rect 11152 44328 11204 44334
rect 11152 44270 11204 44276
rect 11164 43178 11192 44270
rect 11532 44198 11560 44338
rect 11520 44192 11572 44198
rect 11520 44134 11572 44140
rect 11244 43648 11296 43654
rect 11244 43590 11296 43596
rect 11152 43172 11204 43178
rect 11152 43114 11204 43120
rect 11152 42220 11204 42226
rect 11152 42162 11204 42168
rect 11060 41812 11112 41818
rect 11060 41754 11112 41760
rect 11060 41472 11112 41478
rect 11060 41414 11112 41420
rect 10968 40112 11020 40118
rect 10968 40054 11020 40060
rect 10968 39976 11020 39982
rect 10968 39918 11020 39924
rect 10876 39636 10928 39642
rect 10876 39578 10928 39584
rect 10784 38956 10836 38962
rect 10784 38898 10836 38904
rect 10888 38418 10916 39578
rect 10980 39098 11008 39918
rect 10968 39092 11020 39098
rect 10968 39034 11020 39040
rect 11072 38554 11100 41414
rect 11164 38826 11192 42162
rect 11152 38820 11204 38826
rect 11152 38762 11204 38768
rect 11060 38548 11112 38554
rect 11060 38490 11112 38496
rect 10876 38412 10928 38418
rect 10876 38354 10928 38360
rect 10784 38208 10836 38214
rect 10784 38150 10836 38156
rect 10876 38208 10928 38214
rect 10876 38150 10928 38156
rect 10796 38010 10824 38150
rect 10784 38004 10836 38010
rect 10784 37946 10836 37952
rect 10416 37460 10468 37466
rect 10416 37402 10468 37408
rect 10428 37262 10456 37402
rect 10416 37256 10468 37262
rect 10416 37198 10468 37204
rect 10428 36854 10456 37198
rect 10508 37120 10560 37126
rect 10508 37062 10560 37068
rect 10416 36848 10468 36854
rect 10416 36790 10468 36796
rect 10140 36168 10192 36174
rect 10140 36110 10192 36116
rect 10324 36032 10376 36038
rect 10324 35974 10376 35980
rect 10232 35488 10284 35494
rect 10232 35430 10284 35436
rect 10140 34944 10192 34950
rect 10140 34886 10192 34892
rect 10152 32026 10180 34886
rect 10244 34474 10272 35430
rect 10232 34468 10284 34474
rect 10232 34410 10284 34416
rect 10336 33658 10364 35974
rect 10416 34536 10468 34542
rect 10416 34478 10468 34484
rect 10428 33998 10456 34478
rect 10416 33992 10468 33998
rect 10416 33934 10468 33940
rect 10324 33652 10376 33658
rect 10324 33594 10376 33600
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 10048 30184 10100 30190
rect 10048 30126 10100 30132
rect 10416 30048 10468 30054
rect 10416 29990 10468 29996
rect 10428 29850 10456 29990
rect 10416 29844 10468 29850
rect 10416 29786 10468 29792
rect 9956 29572 10008 29578
rect 9956 29514 10008 29520
rect 9772 29300 9824 29306
rect 9772 29242 9824 29248
rect 9784 29102 9812 29242
rect 9404 29096 9456 29102
rect 9404 29038 9456 29044
rect 9772 29096 9824 29102
rect 9772 29038 9824 29044
rect 9416 28558 9444 29038
rect 9864 28620 9916 28626
rect 9864 28562 9916 28568
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9416 26926 9444 28494
rect 9588 28416 9640 28422
rect 9588 28358 9640 28364
rect 9600 28082 9628 28358
rect 9588 28076 9640 28082
rect 9588 28018 9640 28024
rect 9876 27674 9904 28562
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 9968 27878 9996 28494
rect 9956 27872 10008 27878
rect 9956 27814 10008 27820
rect 9864 27668 9916 27674
rect 9864 27610 9916 27616
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9680 26852 9732 26858
rect 9680 26794 9732 26800
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9416 25362 9444 25842
rect 9692 25362 9720 26794
rect 9876 25838 9904 27610
rect 9968 27470 9996 27814
rect 9956 27464 10008 27470
rect 9956 27406 10008 27412
rect 9968 26382 9996 27406
rect 10520 27062 10548 37062
rect 10600 36780 10652 36786
rect 10600 36722 10652 36728
rect 10612 35290 10640 36722
rect 10784 36576 10836 36582
rect 10784 36518 10836 36524
rect 10600 35284 10652 35290
rect 10600 35226 10652 35232
rect 10692 34196 10744 34202
rect 10692 34138 10744 34144
rect 10600 33312 10652 33318
rect 10600 33254 10652 33260
rect 10612 33114 10640 33254
rect 10600 33108 10652 33114
rect 10600 33050 10652 33056
rect 10612 32774 10640 33050
rect 10600 32768 10652 32774
rect 10600 32710 10652 32716
rect 10704 30818 10732 34138
rect 10796 33658 10824 36518
rect 10784 33652 10836 33658
rect 10784 33594 10836 33600
rect 10888 33114 10916 38150
rect 11256 37330 11284 43590
rect 11532 41426 11560 44134
rect 11624 43994 11652 44406
rect 11612 43988 11664 43994
rect 11612 43930 11664 43936
rect 11532 41398 11652 41426
rect 11336 40928 11388 40934
rect 11336 40870 11388 40876
rect 11348 40662 11376 40870
rect 11336 40656 11388 40662
rect 11336 40598 11388 40604
rect 11428 40384 11480 40390
rect 11428 40326 11480 40332
rect 11440 38418 11468 40326
rect 11520 39364 11572 39370
rect 11520 39306 11572 39312
rect 11428 38412 11480 38418
rect 11428 38354 11480 38360
rect 11334 38312 11390 38321
rect 11334 38247 11390 38256
rect 11244 37324 11296 37330
rect 11244 37266 11296 37272
rect 10968 36712 11020 36718
rect 10968 36654 11020 36660
rect 10980 35630 11008 36654
rect 10968 35624 11020 35630
rect 10968 35566 11020 35572
rect 10980 34542 11008 35566
rect 11060 35148 11112 35154
rect 11060 35090 11112 35096
rect 10968 34536 11020 34542
rect 10968 34478 11020 34484
rect 10968 34400 11020 34406
rect 11072 34354 11100 35090
rect 11020 34348 11100 34354
rect 10968 34342 11100 34348
rect 10980 34326 11100 34342
rect 10876 33108 10928 33114
rect 10876 33050 10928 33056
rect 11152 32972 11204 32978
rect 11152 32914 11204 32920
rect 11060 32360 11112 32366
rect 11060 32302 11112 32308
rect 10968 32224 11020 32230
rect 10968 32166 11020 32172
rect 10980 31754 11008 32166
rect 11072 31906 11100 32302
rect 11164 32026 11192 32914
rect 11152 32020 11204 32026
rect 11152 31962 11204 31968
rect 11072 31878 11192 31906
rect 11060 31816 11112 31822
rect 11060 31758 11112 31764
rect 10968 31748 11020 31754
rect 10968 31690 11020 31696
rect 10612 30802 10732 30818
rect 10600 30796 10732 30802
rect 10652 30790 10732 30796
rect 10600 30738 10652 30744
rect 10600 30184 10652 30190
rect 10600 30126 10652 30132
rect 10508 27056 10560 27062
rect 10508 26998 10560 27004
rect 10232 26852 10284 26858
rect 10232 26794 10284 26800
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9864 25832 9916 25838
rect 9864 25774 9916 25780
rect 9404 25356 9456 25362
rect 9404 25298 9456 25304
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 9312 24744 9364 24750
rect 9312 24686 9364 24692
rect 9680 24744 9732 24750
rect 9680 24686 9732 24692
rect 9324 24410 9352 24686
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9692 23866 9720 24686
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 9784 23866 9812 24006
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9968 23594 9996 26318
rect 10048 24268 10100 24274
rect 10048 24210 10100 24216
rect 9956 23588 10008 23594
rect 9956 23530 10008 23536
rect 9680 23248 9732 23254
rect 9680 23190 9732 23196
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9324 22778 9352 23054
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9404 22500 9456 22506
rect 9404 22442 9456 22448
rect 8956 22066 9076 22094
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8956 20602 8984 21490
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8864 19922 8892 20538
rect 9048 20482 9076 22066
rect 9128 21480 9180 21486
rect 9128 21422 9180 21428
rect 8956 20466 9076 20482
rect 8944 20460 9076 20466
rect 8996 20454 9076 20460
rect 8944 20402 8996 20408
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 8956 19802 8984 20402
rect 9140 20262 9168 21422
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 8864 19774 8984 19802
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 8864 19718 8892 19774
rect 9048 19718 9076 19790
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8588 18630 8616 19314
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8588 15162 8616 18566
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8680 12986 8708 18022
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8772 12782 8800 13126
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8864 12434 8892 19654
rect 9416 19514 9444 22442
rect 9692 21690 9720 23190
rect 9968 22982 9996 23530
rect 9956 22976 10008 22982
rect 9956 22918 10008 22924
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9588 20392 9640 20398
rect 9588 20334 9640 20340
rect 9600 20262 9628 20334
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9876 19938 9904 22714
rect 9968 20874 9996 22918
rect 10060 21010 10088 24210
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9876 19910 10088 19938
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 9048 16794 9076 17138
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 8772 12406 8892 12434
rect 8944 12436 8996 12442
rect 8772 5710 8800 12406
rect 8944 12378 8996 12384
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8680 3058 8708 3334
rect 8260 3012 8340 3040
rect 8208 2994 8260 3000
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 7852 1958 7972 1986
rect 7944 800 7972 1958
rect 8312 800 8340 3012
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8680 800 8708 2994
rect 8956 2582 8984 12378
rect 9140 7818 9168 18566
rect 9232 16658 9260 19246
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9324 18358 9352 18702
rect 9312 18352 9364 18358
rect 9312 18294 9364 18300
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9784 18086 9812 18226
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9784 17746 9812 18022
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9324 16590 9352 17546
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9324 15162 9352 15642
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9416 15094 9444 17682
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9508 17338 9536 17478
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 16561 9536 16934
rect 9600 16590 9628 17478
rect 9588 16584 9640 16590
rect 9494 16552 9550 16561
rect 9588 16526 9640 16532
rect 9494 16487 9550 16496
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9404 15088 9456 15094
rect 9456 15048 9536 15076
rect 9404 15030 9456 15036
rect 9508 13870 9536 15048
rect 9784 14006 9812 15098
rect 9876 14618 9904 18022
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9968 14482 9996 14758
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9600 12102 9628 13874
rect 9784 13462 9812 13942
rect 9876 13734 9904 14214
rect 9968 14074 9996 14418
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9864 13388 9916 13394
rect 9968 13376 9996 14010
rect 9916 13348 9996 13376
rect 9864 13330 9916 13336
rect 9968 12918 9996 13348
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 9692 12238 9720 12854
rect 10060 12434 10088 19910
rect 10244 16454 10272 26794
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 10520 26042 10548 26726
rect 10508 26036 10560 26042
rect 10508 25978 10560 25984
rect 10508 24064 10560 24070
rect 10508 24006 10560 24012
rect 10520 23866 10548 24006
rect 10508 23860 10560 23866
rect 10508 23802 10560 23808
rect 10612 22094 10640 30126
rect 10704 30122 10732 30790
rect 10692 30116 10744 30122
rect 10692 30058 10744 30064
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10704 25140 10732 29446
rect 10796 25294 10824 29446
rect 10876 29028 10928 29034
rect 10876 28970 10928 28976
rect 10888 26042 10916 28970
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 10980 26994 11008 27406
rect 11072 27130 11100 31758
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 11164 26908 11192 31878
rect 11348 31822 11376 38247
rect 11426 38176 11482 38185
rect 11426 38111 11482 38120
rect 11440 33454 11468 38111
rect 11532 36310 11560 39306
rect 11520 36304 11572 36310
rect 11520 36246 11572 36252
rect 11428 33448 11480 33454
rect 11428 33390 11480 33396
rect 11532 32978 11560 36246
rect 11624 33674 11652 41398
rect 11716 41274 11744 45834
rect 11808 42362 11836 47602
rect 12164 46912 12216 46918
rect 12164 46854 12216 46860
rect 11888 46368 11940 46374
rect 11888 46310 11940 46316
rect 11900 46034 11928 46310
rect 12176 46034 12204 46854
rect 11888 46028 11940 46034
rect 11888 45970 11940 45976
rect 12164 46028 12216 46034
rect 12164 45970 12216 45976
rect 12256 45348 12308 45354
rect 12256 45290 12308 45296
rect 12268 44266 12296 45290
rect 12440 45280 12492 45286
rect 12440 45222 12492 45228
rect 12452 44878 12480 45222
rect 12544 45082 12572 48690
rect 12532 45076 12584 45082
rect 12532 45018 12584 45024
rect 12624 44940 12676 44946
rect 12624 44882 12676 44888
rect 12440 44872 12492 44878
rect 12440 44814 12492 44820
rect 12348 44464 12400 44470
rect 12348 44406 12400 44412
rect 12256 44260 12308 44266
rect 12256 44202 12308 44208
rect 11888 43716 11940 43722
rect 11888 43658 11940 43664
rect 11796 42356 11848 42362
rect 11796 42298 11848 42304
rect 11900 42242 11928 43658
rect 12164 43104 12216 43110
rect 12164 43046 12216 43052
rect 12176 42702 12204 43046
rect 12164 42696 12216 42702
rect 12164 42638 12216 42644
rect 11808 42214 11928 42242
rect 11704 41268 11756 41274
rect 11704 41210 11756 41216
rect 11704 38752 11756 38758
rect 11704 38694 11756 38700
rect 11716 37262 11744 38694
rect 11704 37256 11756 37262
rect 11704 37198 11756 37204
rect 11624 33646 11744 33674
rect 11612 33516 11664 33522
rect 11612 33458 11664 33464
rect 11520 32972 11572 32978
rect 11520 32914 11572 32920
rect 11624 32026 11652 33458
rect 11716 32842 11744 33646
rect 11808 33590 11836 42214
rect 11888 41608 11940 41614
rect 11888 41550 11940 41556
rect 11900 36378 11928 41550
rect 12072 41132 12124 41138
rect 12072 41074 12124 41080
rect 11980 39024 12032 39030
rect 11980 38966 12032 38972
rect 11992 37330 12020 38966
rect 12084 37738 12112 41074
rect 12268 41070 12296 44202
rect 12360 43314 12388 44406
rect 12348 43308 12400 43314
rect 12348 43250 12400 43256
rect 12360 42770 12388 43250
rect 12452 42838 12480 44814
rect 12636 43382 12664 44882
rect 12624 43376 12676 43382
rect 12624 43318 12676 43324
rect 12440 42832 12492 42838
rect 12440 42774 12492 42780
rect 12348 42764 12400 42770
rect 12348 42706 12400 42712
rect 12360 41682 12388 42706
rect 12624 42696 12676 42702
rect 12624 42638 12676 42644
rect 12636 42566 12664 42638
rect 12440 42560 12492 42566
rect 12440 42502 12492 42508
rect 12624 42560 12676 42566
rect 12624 42502 12676 42508
rect 12452 42158 12480 42502
rect 12440 42152 12492 42158
rect 12440 42094 12492 42100
rect 12532 42152 12584 42158
rect 12532 42094 12584 42100
rect 12348 41676 12400 41682
rect 12348 41618 12400 41624
rect 12256 41064 12308 41070
rect 12256 41006 12308 41012
rect 12256 40928 12308 40934
rect 12256 40870 12308 40876
rect 12268 39438 12296 40870
rect 12438 40488 12494 40497
rect 12438 40423 12440 40432
rect 12492 40423 12494 40432
rect 12440 40394 12492 40400
rect 12452 40202 12480 40394
rect 12360 40174 12480 40202
rect 12256 39432 12308 39438
rect 12256 39374 12308 39380
rect 12360 39386 12388 40174
rect 12360 39358 12480 39386
rect 12256 39296 12308 39302
rect 12256 39238 12308 39244
rect 12268 39098 12296 39238
rect 12256 39092 12308 39098
rect 12256 39034 12308 39040
rect 12256 38208 12308 38214
rect 12256 38150 12308 38156
rect 12072 37732 12124 37738
rect 12072 37674 12124 37680
rect 12164 37732 12216 37738
rect 12164 37674 12216 37680
rect 12176 37398 12204 37674
rect 12164 37392 12216 37398
rect 12164 37334 12216 37340
rect 11980 37324 12032 37330
rect 11980 37266 12032 37272
rect 11980 36644 12032 36650
rect 11980 36586 12032 36592
rect 11888 36372 11940 36378
rect 11888 36314 11940 36320
rect 11992 34406 12020 36586
rect 12162 36272 12218 36281
rect 12162 36207 12218 36216
rect 11980 34400 12032 34406
rect 11980 34342 12032 34348
rect 11796 33584 11848 33590
rect 11796 33526 11848 33532
rect 11704 32836 11756 32842
rect 11704 32778 11756 32784
rect 11888 32768 11940 32774
rect 11888 32710 11940 32716
rect 11612 32020 11664 32026
rect 11612 31962 11664 31968
rect 11336 31816 11388 31822
rect 11336 31758 11388 31764
rect 11612 31816 11664 31822
rect 11612 31758 11664 31764
rect 11624 30870 11652 31758
rect 11900 31754 11928 32710
rect 11992 32298 12020 34342
rect 12072 33992 12124 33998
rect 12072 33934 12124 33940
rect 12084 33862 12112 33934
rect 12072 33856 12124 33862
rect 12072 33798 12124 33804
rect 11980 32292 12032 32298
rect 11980 32234 12032 32240
rect 12084 31822 12112 33798
rect 12176 32366 12204 36207
rect 12268 32502 12296 38150
rect 12452 38010 12480 39358
rect 12440 38004 12492 38010
rect 12440 37946 12492 37952
rect 12438 37768 12494 37777
rect 12438 37703 12494 37712
rect 12452 36530 12480 37703
rect 12360 36502 12480 36530
rect 12360 35222 12388 36502
rect 12544 36378 12572 42094
rect 12636 40934 12664 42502
rect 12624 40928 12676 40934
rect 12624 40870 12676 40876
rect 12728 40526 12756 49710
rect 12820 48890 12848 52430
rect 13372 52426 13400 55186
rect 13648 53174 13676 56200
rect 14016 53582 14044 56200
rect 14096 53984 14148 53990
rect 14096 53926 14148 53932
rect 14004 53576 14056 53582
rect 14004 53518 14056 53524
rect 13636 53168 13688 53174
rect 13636 53110 13688 53116
rect 13648 52698 13676 53110
rect 14004 52964 14056 52970
rect 14004 52906 14056 52912
rect 13636 52692 13688 52698
rect 13636 52634 13688 52640
rect 14016 52601 14044 52906
rect 14002 52592 14058 52601
rect 14002 52527 14058 52536
rect 13544 52488 13596 52494
rect 13544 52430 13596 52436
rect 13360 52420 13412 52426
rect 13360 52362 13412 52368
rect 13372 52154 13400 52362
rect 13360 52148 13412 52154
rect 13360 52090 13412 52096
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12808 48884 12860 48890
rect 12808 48826 12860 48832
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 13360 46368 13412 46374
rect 13360 46310 13412 46316
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 13372 44470 13400 46310
rect 13452 44872 13504 44878
rect 13452 44814 13504 44820
rect 13360 44464 13412 44470
rect 13360 44406 13412 44412
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 13464 42362 13492 44814
rect 13452 42356 13504 42362
rect 13452 42298 13504 42304
rect 13452 42016 13504 42022
rect 13452 41958 13504 41964
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 12808 41676 12860 41682
rect 12808 41618 12860 41624
rect 12716 40520 12768 40526
rect 12716 40462 12768 40468
rect 12820 40050 12848 41618
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 13360 40656 13412 40662
rect 13360 40598 13412 40604
rect 12716 40044 12768 40050
rect 12716 39986 12768 39992
rect 12808 40044 12860 40050
rect 12808 39986 12860 39992
rect 12728 39574 12756 39986
rect 12716 39568 12768 39574
rect 12716 39510 12768 39516
rect 12820 39506 12848 39986
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12900 39636 12952 39642
rect 12900 39578 12952 39584
rect 13084 39636 13136 39642
rect 13084 39578 13136 39584
rect 12624 39500 12676 39506
rect 12624 39442 12676 39448
rect 12808 39500 12860 39506
rect 12808 39442 12860 39448
rect 12636 39030 12664 39442
rect 12912 39386 12940 39578
rect 13096 39438 13124 39578
rect 12728 39358 12940 39386
rect 13084 39432 13136 39438
rect 13084 39374 13136 39380
rect 12728 39302 12756 39358
rect 12716 39296 12768 39302
rect 12716 39238 12768 39244
rect 12624 39024 12676 39030
rect 12624 38966 12676 38972
rect 12622 38448 12678 38457
rect 12728 38418 12756 39238
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12622 38383 12678 38392
rect 12716 38412 12768 38418
rect 12440 36372 12492 36378
rect 12440 36314 12492 36320
rect 12532 36372 12584 36378
rect 12636 36360 12664 38383
rect 12716 38354 12768 38360
rect 12808 37664 12860 37670
rect 12808 37606 12860 37612
rect 12820 37194 12848 37606
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12808 37188 12860 37194
rect 12808 37130 12860 37136
rect 12716 37120 12768 37126
rect 12716 37062 12768 37068
rect 12728 36786 12756 37062
rect 12716 36780 12768 36786
rect 12716 36722 12768 36728
rect 12728 36689 12756 36722
rect 12808 36712 12860 36718
rect 12714 36680 12770 36689
rect 12808 36654 12860 36660
rect 12714 36615 12770 36624
rect 12636 36332 12756 36360
rect 12532 36314 12584 36320
rect 12452 36258 12480 36314
rect 12452 36230 12664 36258
rect 12728 36242 12756 36332
rect 12440 36168 12492 36174
rect 12440 36110 12492 36116
rect 12452 36038 12480 36110
rect 12636 36038 12664 36230
rect 12716 36236 12768 36242
rect 12716 36178 12768 36184
rect 12716 36100 12768 36106
rect 12716 36042 12768 36048
rect 12440 36032 12492 36038
rect 12440 35974 12492 35980
rect 12624 36032 12676 36038
rect 12624 35974 12676 35980
rect 12452 35873 12480 35974
rect 12438 35864 12494 35873
rect 12438 35799 12494 35808
rect 12348 35216 12400 35222
rect 12348 35158 12400 35164
rect 12532 33924 12584 33930
rect 12532 33866 12584 33872
rect 12440 33516 12492 33522
rect 12440 33458 12492 33464
rect 12256 32496 12308 32502
rect 12256 32438 12308 32444
rect 12164 32360 12216 32366
rect 12164 32302 12216 32308
rect 12072 31816 12124 31822
rect 12072 31758 12124 31764
rect 11900 31726 12020 31754
rect 11612 30864 11664 30870
rect 11612 30806 11664 30812
rect 11244 30728 11296 30734
rect 11244 30670 11296 30676
rect 11256 30326 11284 30670
rect 11336 30592 11388 30598
rect 11336 30534 11388 30540
rect 11244 30320 11296 30326
rect 11244 30262 11296 30268
rect 11348 29782 11376 30534
rect 11796 30388 11848 30394
rect 11796 30330 11848 30336
rect 11336 29776 11388 29782
rect 11336 29718 11388 29724
rect 11244 29300 11296 29306
rect 11244 29242 11296 29248
rect 11072 26880 11192 26908
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 10704 25112 10824 25140
rect 10796 23050 10824 25112
rect 10968 24132 11020 24138
rect 10968 24074 11020 24080
rect 10876 23316 10928 23322
rect 10876 23258 10928 23264
rect 10784 23044 10836 23050
rect 10784 22986 10836 22992
rect 10692 22094 10744 22098
rect 10612 22092 10744 22094
rect 10612 22066 10692 22092
rect 10692 22034 10744 22040
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10336 20874 10364 21286
rect 10324 20868 10376 20874
rect 10324 20810 10376 20816
rect 10336 18290 10364 20810
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10428 18426 10456 20742
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10336 17134 10364 18226
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10244 16130 10272 16390
rect 10152 16102 10272 16130
rect 10152 14226 10180 16102
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10244 15366 10272 15982
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10244 14346 10272 15302
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 10152 14198 10272 14226
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10152 12442 10180 14010
rect 9876 12406 10088 12434
rect 10140 12436 10192 12442
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9876 10470 9904 12406
rect 10140 12378 10192 12384
rect 10244 12170 10272 14198
rect 10232 12164 10284 12170
rect 10232 12106 10284 12112
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 9048 2990 9076 3946
rect 9324 3058 9352 5510
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9416 3534 9444 3878
rect 9508 3738 9536 9590
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9784 3534 9812 3878
rect 10060 3738 10088 5578
rect 10336 4214 10364 16934
rect 10520 16250 10548 17070
rect 10612 16250 10640 21898
rect 10704 21894 10732 22034
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10704 16130 10732 21830
rect 10796 16998 10824 22986
rect 10888 22778 10916 23258
rect 10876 22772 10928 22778
rect 10876 22714 10928 22720
rect 10980 22658 11008 24074
rect 10888 22630 11008 22658
rect 10888 21350 10916 22630
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 10980 20806 11008 22510
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 10876 19168 10928 19174
rect 10874 19136 10876 19145
rect 10928 19136 10930 19145
rect 10874 19071 10930 19080
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10888 16726 10916 17070
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10612 16102 10732 16130
rect 10428 13938 10456 16050
rect 10612 14226 10640 16102
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10612 14198 10732 14226
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10704 11830 10732 14198
rect 10796 14074 10824 14554
rect 10888 14278 10916 16662
rect 10980 16250 11008 20470
rect 11072 19310 11100 26880
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 11164 24206 11192 24550
rect 11256 24274 11284 29242
rect 11348 28626 11376 29718
rect 11808 29646 11836 30330
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11796 29640 11848 29646
rect 11796 29582 11848 29588
rect 11900 29510 11928 29990
rect 11888 29504 11940 29510
rect 11888 29446 11940 29452
rect 11336 28620 11388 28626
rect 11336 28562 11388 28568
rect 11796 27940 11848 27946
rect 11796 27882 11848 27888
rect 11428 27396 11480 27402
rect 11428 27338 11480 27344
rect 11336 27056 11388 27062
rect 11336 26998 11388 27004
rect 11348 26790 11376 26998
rect 11336 26784 11388 26790
rect 11336 26726 11388 26732
rect 11348 26382 11376 26726
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 11164 20398 11192 24006
rect 11244 23860 11296 23866
rect 11244 23802 11296 23808
rect 11152 20392 11204 20398
rect 11152 20334 11204 20340
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11072 18630 11100 19110
rect 11164 18970 11192 19110
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11060 18216 11112 18222
rect 11058 18184 11060 18193
rect 11112 18184 11114 18193
rect 11058 18119 11114 18128
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10968 15972 11020 15978
rect 10968 15914 11020 15920
rect 10980 15434 11008 15914
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10980 15094 11008 15370
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 11256 14006 11284 23802
rect 11348 23526 11376 26318
rect 11440 25702 11468 27338
rect 11704 27328 11756 27334
rect 11704 27270 11756 27276
rect 11520 27124 11572 27130
rect 11520 27066 11572 27072
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11428 25696 11480 25702
rect 11428 25638 11480 25644
rect 11440 25362 11468 25638
rect 11428 25356 11480 25362
rect 11428 25298 11480 25304
rect 11532 24138 11560 27066
rect 11624 26926 11652 27066
rect 11612 26920 11664 26926
rect 11612 26862 11664 26868
rect 11716 26450 11744 27270
rect 11808 26450 11836 27882
rect 11704 26444 11756 26450
rect 11704 26386 11756 26392
rect 11796 26444 11848 26450
rect 11796 26386 11848 26392
rect 11796 25832 11848 25838
rect 11796 25774 11848 25780
rect 11808 25294 11836 25774
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11520 24132 11572 24138
rect 11520 24074 11572 24080
rect 11532 23866 11560 24074
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11900 23798 11928 29446
rect 11992 25158 12020 31726
rect 12452 26466 12480 33458
rect 12544 30938 12572 33866
rect 12636 33522 12664 35974
rect 12728 33658 12756 36042
rect 12820 34746 12848 36654
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 13372 35465 13400 40598
rect 13464 38457 13492 41958
rect 13556 40712 13584 52430
rect 13912 46912 13964 46918
rect 13912 46854 13964 46860
rect 13924 46646 13952 46854
rect 13912 46640 13964 46646
rect 13912 46582 13964 46588
rect 13728 46368 13780 46374
rect 13728 46310 13780 46316
rect 13636 45824 13688 45830
rect 13636 45766 13688 45772
rect 13648 44198 13676 45766
rect 13740 44946 13768 46310
rect 13924 45898 13952 46582
rect 13912 45892 13964 45898
rect 13912 45834 13964 45840
rect 13728 44940 13780 44946
rect 13728 44882 13780 44888
rect 13636 44192 13688 44198
rect 13636 44134 13688 44140
rect 13648 42022 13676 44134
rect 13728 43308 13780 43314
rect 13728 43250 13780 43256
rect 13740 42566 13768 43250
rect 13728 42560 13780 42566
rect 13728 42502 13780 42508
rect 13636 42016 13688 42022
rect 13636 41958 13688 41964
rect 13636 41676 13688 41682
rect 13636 41618 13688 41624
rect 13648 41138 13676 41618
rect 13636 41132 13688 41138
rect 13636 41074 13688 41080
rect 14004 41064 14056 41070
rect 14004 41006 14056 41012
rect 13556 40684 13768 40712
rect 13636 40588 13688 40594
rect 13636 40530 13688 40536
rect 13450 38448 13506 38457
rect 13450 38383 13506 38392
rect 13452 37800 13504 37806
rect 13452 37742 13504 37748
rect 13544 37800 13596 37806
rect 13544 37742 13596 37748
rect 13464 37074 13492 37742
rect 13556 37262 13584 37742
rect 13544 37256 13596 37262
rect 13544 37198 13596 37204
rect 13464 37046 13584 37074
rect 13452 36780 13504 36786
rect 13452 36722 13504 36728
rect 13464 35873 13492 36722
rect 13450 35864 13506 35873
rect 13556 35834 13584 37046
rect 13450 35799 13506 35808
rect 13544 35828 13596 35834
rect 13544 35770 13596 35776
rect 13358 35456 13414 35465
rect 12950 35388 13258 35397
rect 13358 35391 13414 35400
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 13452 35216 13504 35222
rect 13358 35184 13414 35193
rect 13452 35158 13504 35164
rect 13358 35119 13414 35128
rect 12808 34740 12860 34746
rect 12808 34682 12860 34688
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 13372 34066 13400 35119
rect 13360 34060 13412 34066
rect 13360 34002 13412 34008
rect 13464 33946 13492 35158
rect 13372 33918 13492 33946
rect 12808 33856 12860 33862
rect 12808 33798 12860 33804
rect 13176 33856 13228 33862
rect 13176 33798 13228 33804
rect 12716 33652 12768 33658
rect 12716 33594 12768 33600
rect 12624 33516 12676 33522
rect 12624 33458 12676 33464
rect 12716 33516 12768 33522
rect 12716 33458 12768 33464
rect 12624 33380 12676 33386
rect 12624 33322 12676 33328
rect 12636 30977 12664 33322
rect 12622 30968 12678 30977
rect 12532 30932 12584 30938
rect 12622 30903 12678 30912
rect 12532 30874 12584 30880
rect 12532 28484 12584 28490
rect 12532 28426 12584 28432
rect 12544 28082 12572 28426
rect 12532 28076 12584 28082
rect 12532 28018 12584 28024
rect 12624 27872 12676 27878
rect 12624 27814 12676 27820
rect 12636 27146 12664 27814
rect 12544 27130 12664 27146
rect 12532 27124 12664 27130
rect 12584 27118 12664 27124
rect 12532 27066 12584 27072
rect 12360 26438 12480 26466
rect 12360 25838 12388 26438
rect 12544 26364 12572 27066
rect 12452 26336 12572 26364
rect 12348 25832 12400 25838
rect 12348 25774 12400 25780
rect 12256 25764 12308 25770
rect 12256 25706 12308 25712
rect 12268 25514 12296 25706
rect 12268 25486 12388 25514
rect 12256 25424 12308 25430
rect 12256 25366 12308 25372
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 11980 24064 12032 24070
rect 12176 24041 12204 24074
rect 11980 24006 12032 24012
rect 12162 24032 12218 24041
rect 11888 23792 11940 23798
rect 11888 23734 11940 23740
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11612 23588 11664 23594
rect 11612 23530 11664 23536
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11348 20942 11376 23462
rect 11624 23118 11652 23530
rect 11716 23118 11744 23598
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11612 22704 11664 22710
rect 11612 22646 11664 22652
rect 11624 22438 11652 22646
rect 11612 22432 11664 22438
rect 11612 22374 11664 22380
rect 11900 21570 11928 23122
rect 11992 21690 12020 24006
rect 12162 23967 12218 23976
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 12084 23526 12112 23598
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 12084 22982 12112 23462
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11900 21542 12020 21570
rect 11888 21480 11940 21486
rect 11888 21422 11940 21428
rect 11520 21412 11572 21418
rect 11520 21354 11572 21360
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11348 19174 11376 20878
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11348 17134 11376 17546
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11348 15570 11376 17070
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11348 14550 11376 15506
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10980 10742 11008 12582
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 8944 2576 8996 2582
rect 8944 2518 8996 2524
rect 9048 800 9076 2926
rect 9416 800 9444 3470
rect 9784 800 9812 3470
rect 10520 2990 10548 3878
rect 11256 3602 11284 6326
rect 11440 5574 11468 19722
rect 11532 18154 11560 21354
rect 11900 21010 11928 21422
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11612 20324 11664 20330
rect 11612 20266 11664 20272
rect 11624 19514 11652 20266
rect 11716 20058 11744 20402
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11716 18358 11744 19110
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11808 18170 11836 18566
rect 11900 18290 11928 20946
rect 11992 20602 12020 21542
rect 12084 21146 12112 22918
rect 12162 22808 12218 22817
rect 12162 22743 12218 22752
rect 12176 22710 12204 22743
rect 12164 22704 12216 22710
rect 12164 22646 12216 22652
rect 12164 22092 12216 22098
rect 12164 22034 12216 22040
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11992 20058 12020 20538
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11520 18148 11572 18154
rect 11808 18142 11928 18170
rect 11520 18090 11572 18096
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11532 13530 11560 17002
rect 11624 15042 11652 17546
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11716 15706 11744 16390
rect 11808 16182 11836 16390
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11900 16046 11928 18142
rect 11992 16590 12020 18566
rect 12084 17338 12112 20198
rect 12176 19990 12204 22034
rect 12268 20534 12296 25366
rect 12360 21418 12388 25486
rect 12452 24698 12480 26336
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12544 25974 12572 26182
rect 12532 25968 12584 25974
rect 12532 25910 12584 25916
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 12544 25226 12572 25774
rect 12532 25220 12584 25226
rect 12532 25162 12584 25168
rect 12544 24834 12572 25162
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12636 24954 12664 25094
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12544 24806 12664 24834
rect 12452 24682 12572 24698
rect 12452 24676 12584 24682
rect 12452 24670 12532 24676
rect 12532 24618 12584 24624
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12452 23866 12480 24550
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12440 23520 12492 23526
rect 12544 23508 12572 24618
rect 12636 24614 12664 24806
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 12492 23480 12572 23508
rect 12440 23462 12492 23468
rect 12440 23248 12492 23254
rect 12440 23190 12492 23196
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12256 20528 12308 20534
rect 12256 20470 12308 20476
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12164 19984 12216 19990
rect 12164 19926 12216 19932
rect 12268 19922 12296 19994
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12162 19408 12218 19417
rect 12162 19343 12218 19352
rect 12176 18970 12204 19343
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12176 18426 12204 18906
rect 12268 18698 12296 19858
rect 12452 19854 12480 23190
rect 12544 22778 12572 23480
rect 12636 23322 12664 24550
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12346 19272 12402 19281
rect 12346 19207 12402 19216
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 12176 15162 12204 18158
rect 12360 18154 12388 19207
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 18222 12480 19110
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 12360 18034 12388 18090
rect 12268 18006 12388 18034
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 11980 15088 12032 15094
rect 11624 15014 11744 15042
rect 11980 15030 12032 15036
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11532 12434 11560 13466
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11624 12918 11652 13194
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11532 12406 11652 12434
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11532 11762 11560 12174
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11624 8362 11652 12406
rect 11716 9382 11744 15014
rect 11992 14550 12020 15030
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11808 12986 11836 13738
rect 11992 13530 12020 14486
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11992 13258 12020 13466
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11808 12306 11836 12922
rect 12176 12442 12204 14010
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12268 12322 12296 18006
rect 12452 16130 12480 18158
rect 12544 16250 12572 22374
rect 12728 22094 12756 33458
rect 12820 29646 12848 33798
rect 13188 33522 13216 33798
rect 13176 33516 13228 33522
rect 13176 33458 13228 33464
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 13372 31482 13400 33918
rect 13556 33454 13584 35770
rect 13648 35562 13676 40530
rect 13740 35714 13768 40684
rect 13820 39296 13872 39302
rect 13820 39238 13872 39244
rect 13832 38321 13860 39238
rect 13912 38752 13964 38758
rect 13912 38694 13964 38700
rect 13818 38312 13874 38321
rect 13818 38247 13874 38256
rect 13924 36718 13952 38694
rect 14016 37466 14044 41006
rect 14004 37460 14056 37466
rect 14004 37402 14056 37408
rect 13912 36712 13964 36718
rect 13912 36654 13964 36660
rect 14108 36394 14136 53926
rect 14384 53106 14412 56200
rect 14752 54330 14780 56200
rect 14740 54324 14792 54330
rect 14740 54266 14792 54272
rect 15120 54176 15148 56200
rect 15200 54188 15252 54194
rect 15120 54148 15200 54176
rect 15200 54130 15252 54136
rect 15384 54052 15436 54058
rect 15384 53994 15436 54000
rect 15292 53984 15344 53990
rect 15292 53926 15344 53932
rect 14464 53440 14516 53446
rect 14464 53382 14516 53388
rect 14372 53100 14424 53106
rect 14372 53042 14424 53048
rect 14476 53009 14504 53382
rect 14462 53000 14518 53009
rect 14462 52935 14518 52944
rect 14464 52896 14516 52902
rect 14464 52838 14516 52844
rect 14188 46708 14240 46714
rect 14188 46650 14240 46656
rect 14200 44334 14228 46650
rect 14188 44328 14240 44334
rect 14188 44270 14240 44276
rect 14200 42090 14228 44270
rect 14476 43450 14504 52838
rect 15016 45824 15068 45830
rect 15016 45766 15068 45772
rect 14832 45280 14884 45286
rect 14832 45222 14884 45228
rect 14844 44878 14872 45222
rect 14832 44872 14884 44878
rect 14832 44814 14884 44820
rect 14464 43444 14516 43450
rect 14464 43386 14516 43392
rect 14740 43172 14792 43178
rect 14740 43114 14792 43120
rect 14648 43104 14700 43110
rect 14648 43046 14700 43052
rect 14556 42832 14608 42838
rect 14556 42774 14608 42780
rect 14188 42084 14240 42090
rect 14188 42026 14240 42032
rect 14464 41812 14516 41818
rect 14464 41754 14516 41760
rect 14188 41472 14240 41478
rect 14188 41414 14240 41420
rect 14476 41414 14504 41754
rect 14200 38554 14228 41414
rect 14384 41386 14504 41414
rect 14280 40044 14332 40050
rect 14280 39986 14332 39992
rect 14292 39642 14320 39986
rect 14280 39636 14332 39642
rect 14280 39578 14332 39584
rect 14292 38962 14320 39578
rect 14280 38956 14332 38962
rect 14280 38898 14332 38904
rect 14188 38548 14240 38554
rect 14188 38490 14240 38496
rect 14292 38350 14320 38898
rect 14384 38865 14412 41386
rect 14568 39930 14596 42774
rect 14476 39902 14596 39930
rect 14370 38856 14426 38865
rect 14370 38791 14426 38800
rect 14280 38344 14332 38350
rect 14280 38286 14332 38292
rect 14188 37188 14240 37194
rect 14188 37130 14240 37136
rect 14200 36786 14228 37130
rect 14188 36780 14240 36786
rect 14188 36722 14240 36728
rect 14292 36530 14320 38286
rect 14384 37466 14412 38791
rect 14372 37460 14424 37466
rect 14372 37402 14424 37408
rect 14384 36718 14412 37402
rect 14476 37398 14504 39902
rect 14556 39840 14608 39846
rect 14556 39782 14608 39788
rect 14568 38894 14596 39782
rect 14556 38888 14608 38894
rect 14556 38830 14608 38836
rect 14464 37392 14516 37398
rect 14464 37334 14516 37340
rect 14660 36854 14688 43046
rect 14752 39846 14780 43114
rect 14844 42770 14872 44814
rect 15028 44470 15056 45766
rect 15200 44736 15252 44742
rect 15200 44678 15252 44684
rect 15108 44532 15160 44538
rect 15108 44474 15160 44480
rect 15016 44464 15068 44470
rect 15016 44406 15068 44412
rect 15028 44198 15056 44406
rect 15016 44192 15068 44198
rect 15016 44134 15068 44140
rect 14832 42764 14884 42770
rect 14832 42706 14884 42712
rect 15028 42566 15056 44134
rect 15120 42770 15148 44474
rect 15108 42764 15160 42770
rect 15108 42706 15160 42712
rect 15016 42560 15068 42566
rect 15016 42502 15068 42508
rect 15212 42362 15240 44678
rect 15200 42356 15252 42362
rect 15200 42298 15252 42304
rect 15108 42288 15160 42294
rect 15108 42230 15160 42236
rect 14924 41268 14976 41274
rect 14924 41210 14976 41216
rect 14832 40724 14884 40730
rect 14832 40666 14884 40672
rect 14844 40390 14872 40666
rect 14832 40384 14884 40390
rect 14832 40326 14884 40332
rect 14740 39840 14792 39846
rect 14740 39782 14792 39788
rect 14740 39296 14792 39302
rect 14740 39238 14792 39244
rect 14752 39098 14780 39238
rect 14740 39092 14792 39098
rect 14740 39034 14792 39040
rect 14832 38548 14884 38554
rect 14832 38490 14884 38496
rect 14740 37256 14792 37262
rect 14740 37198 14792 37204
rect 14752 37126 14780 37198
rect 14740 37120 14792 37126
rect 14740 37062 14792 37068
rect 14648 36848 14700 36854
rect 14648 36790 14700 36796
rect 14372 36712 14424 36718
rect 14372 36654 14424 36660
rect 14464 36576 14516 36582
rect 14292 36502 14412 36530
rect 14464 36518 14516 36524
rect 14556 36576 14608 36582
rect 14556 36518 14608 36524
rect 14108 36366 14320 36394
rect 13818 36272 13874 36281
rect 13818 36207 13820 36216
rect 13872 36207 13874 36216
rect 13820 36178 13872 36184
rect 14004 35828 14056 35834
rect 14004 35770 14056 35776
rect 13740 35686 13952 35714
rect 13820 35624 13872 35630
rect 13820 35566 13872 35572
rect 13636 35556 13688 35562
rect 13636 35498 13688 35504
rect 13648 33998 13676 35498
rect 13728 34740 13780 34746
rect 13728 34682 13780 34688
rect 13636 33992 13688 33998
rect 13636 33934 13688 33940
rect 13636 33856 13688 33862
rect 13636 33798 13688 33804
rect 13544 33448 13596 33454
rect 13544 33390 13596 33396
rect 13452 33312 13504 33318
rect 13452 33254 13504 33260
rect 13360 31476 13412 31482
rect 13360 31418 13412 31424
rect 13268 31272 13320 31278
rect 13464 31260 13492 33254
rect 13648 33046 13676 33798
rect 13636 33040 13688 33046
rect 13636 32982 13688 32988
rect 13544 31476 13596 31482
rect 13544 31418 13596 31424
rect 13320 31232 13492 31260
rect 13268 31214 13320 31220
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 12992 29844 13044 29850
rect 12992 29786 13044 29792
rect 12808 29640 12860 29646
rect 12808 29582 12860 29588
rect 13004 29578 13032 29786
rect 12992 29572 13044 29578
rect 12992 29514 13044 29520
rect 13084 29096 13136 29102
rect 13268 29096 13320 29102
rect 13136 29044 13268 29050
rect 13084 29038 13320 29044
rect 13096 29022 13308 29038
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 13372 28626 13400 31232
rect 13556 30734 13584 31418
rect 13544 30728 13596 30734
rect 13544 30670 13596 30676
rect 13542 30560 13598 30569
rect 13542 30495 13598 30504
rect 13452 29028 13504 29034
rect 13452 28970 13504 28976
rect 13360 28620 13412 28626
rect 13360 28562 13412 28568
rect 13084 28484 13136 28490
rect 13084 28426 13136 28432
rect 12808 28416 12860 28422
rect 12808 28358 12860 28364
rect 12820 27538 12848 28358
rect 13096 27878 13124 28426
rect 13176 28416 13228 28422
rect 13176 28358 13228 28364
rect 13188 28218 13216 28358
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 13360 28076 13412 28082
rect 13360 28018 13412 28024
rect 13372 27878 13400 28018
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 13360 27872 13412 27878
rect 13360 27814 13412 27820
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12820 26926 12848 27474
rect 13372 27470 13400 27814
rect 13360 27464 13412 27470
rect 13360 27406 13412 27412
rect 13084 27396 13136 27402
rect 13084 27338 13136 27344
rect 12900 27328 12952 27334
rect 12900 27270 12952 27276
rect 12912 27130 12940 27270
rect 12900 27124 12952 27130
rect 12900 27066 12952 27072
rect 13096 27062 13124 27338
rect 13360 27328 13412 27334
rect 13360 27270 13412 27276
rect 13084 27056 13136 27062
rect 13084 26998 13136 27004
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12820 25362 12848 26862
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12820 24274 12848 25094
rect 13372 24886 13400 27270
rect 13360 24880 13412 24886
rect 13360 24822 13412 24828
rect 13372 24614 13400 24822
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 12808 23860 12860 23866
rect 12808 23802 12860 23808
rect 12820 22438 12848 23802
rect 13372 23526 13400 24550
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13464 22094 13492 28970
rect 13556 27334 13584 30495
rect 13648 28778 13676 32982
rect 13740 31890 13768 34682
rect 13832 34542 13860 35566
rect 13820 34536 13872 34542
rect 13820 34478 13872 34484
rect 13820 34196 13872 34202
rect 13820 34138 13872 34144
rect 13832 33658 13860 34138
rect 13924 33862 13952 35686
rect 14016 34746 14044 35770
rect 14096 35760 14148 35766
rect 14096 35702 14148 35708
rect 14004 34740 14056 34746
rect 14004 34682 14056 34688
rect 14108 33998 14136 35702
rect 14188 34740 14240 34746
rect 14188 34682 14240 34688
rect 14096 33992 14148 33998
rect 14096 33934 14148 33940
rect 13912 33856 13964 33862
rect 13912 33798 13964 33804
rect 14004 33856 14056 33862
rect 14004 33798 14056 33804
rect 13820 33652 13872 33658
rect 13820 33594 13872 33600
rect 14016 33590 14044 33798
rect 14004 33584 14056 33590
rect 14004 33526 14056 33532
rect 14016 33130 14044 33526
rect 13924 33102 14044 33130
rect 13728 31884 13780 31890
rect 13728 31826 13780 31832
rect 13924 31686 13952 33102
rect 14004 32768 14056 32774
rect 14004 32710 14056 32716
rect 13912 31680 13964 31686
rect 13912 31622 13964 31628
rect 13728 29640 13780 29646
rect 13728 29582 13780 29588
rect 13740 29170 13768 29582
rect 13728 29164 13780 29170
rect 13728 29106 13780 29112
rect 13912 29096 13964 29102
rect 13912 29038 13964 29044
rect 13648 28750 13768 28778
rect 13636 28620 13688 28626
rect 13636 28562 13688 28568
rect 13544 27328 13596 27334
rect 13544 27270 13596 27276
rect 13544 26920 13596 26926
rect 13544 26862 13596 26868
rect 13556 25498 13584 26862
rect 13648 26586 13676 28562
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 13740 26466 13768 28750
rect 13924 28370 13952 29038
rect 14016 28506 14044 32710
rect 14200 29170 14228 34682
rect 14292 31260 14320 36366
rect 14384 35834 14412 36502
rect 14372 35828 14424 35834
rect 14372 35770 14424 35776
rect 14476 32978 14504 36518
rect 14568 35086 14596 36518
rect 14844 36242 14872 38490
rect 14936 37126 14964 41210
rect 15016 41132 15068 41138
rect 15016 41074 15068 41080
rect 15028 40186 15056 41074
rect 15120 40186 15148 42230
rect 15200 41676 15252 41682
rect 15200 41618 15252 41624
rect 15212 41070 15240 41618
rect 15200 41064 15252 41070
rect 15200 41006 15252 41012
rect 15200 40384 15252 40390
rect 15200 40326 15252 40332
rect 15016 40180 15068 40186
rect 15016 40122 15068 40128
rect 15108 40180 15160 40186
rect 15108 40122 15160 40128
rect 15016 39364 15068 39370
rect 15016 39306 15068 39312
rect 15028 37330 15056 39306
rect 15212 38350 15240 40326
rect 15200 38344 15252 38350
rect 15200 38286 15252 38292
rect 15200 37800 15252 37806
rect 15200 37742 15252 37748
rect 15212 37330 15240 37742
rect 15016 37324 15068 37330
rect 15016 37266 15068 37272
rect 15108 37324 15160 37330
rect 15108 37266 15160 37272
rect 15200 37324 15252 37330
rect 15200 37266 15252 37272
rect 15120 37126 15148 37266
rect 14924 37120 14976 37126
rect 14924 37062 14976 37068
rect 15108 37120 15160 37126
rect 15108 37062 15160 37068
rect 15212 36854 15240 37266
rect 15200 36848 15252 36854
rect 15200 36790 15252 36796
rect 15108 36712 15160 36718
rect 15108 36654 15160 36660
rect 14832 36236 14884 36242
rect 14832 36178 14884 36184
rect 14648 36032 14700 36038
rect 14648 35974 14700 35980
rect 14660 35834 14688 35974
rect 14648 35828 14700 35834
rect 14648 35770 14700 35776
rect 14556 35080 14608 35086
rect 14556 35022 14608 35028
rect 14832 34536 14884 34542
rect 14832 34478 14884 34484
rect 14740 33924 14792 33930
rect 14740 33866 14792 33872
rect 14556 33652 14608 33658
rect 14556 33594 14608 33600
rect 14464 32972 14516 32978
rect 14464 32914 14516 32920
rect 14464 32768 14516 32774
rect 14464 32710 14516 32716
rect 14476 31754 14504 32710
rect 14568 32434 14596 33594
rect 14648 32768 14700 32774
rect 14648 32710 14700 32716
rect 14660 32570 14688 32710
rect 14648 32564 14700 32570
rect 14648 32506 14700 32512
rect 14556 32428 14608 32434
rect 14556 32370 14608 32376
rect 14568 32230 14596 32370
rect 14556 32224 14608 32230
rect 14556 32166 14608 32172
rect 14752 31754 14780 33866
rect 14844 32978 14872 34478
rect 15120 33114 15148 36654
rect 15108 33108 15160 33114
rect 15108 33050 15160 33056
rect 14832 32972 14884 32978
rect 14832 32914 14884 32920
rect 14476 31726 14596 31754
rect 14372 31272 14424 31278
rect 14292 31232 14372 31260
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14188 29164 14240 29170
rect 14188 29106 14240 29112
rect 14108 28762 14136 29106
rect 14292 29102 14320 31232
rect 14372 31214 14424 31220
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14370 30288 14426 30297
rect 14476 30258 14504 31078
rect 14370 30223 14372 30232
rect 14424 30223 14426 30232
rect 14464 30252 14516 30258
rect 14372 30194 14424 30200
rect 14464 30194 14516 30200
rect 14384 30054 14412 30194
rect 14372 30048 14424 30054
rect 14372 29990 14424 29996
rect 14280 29096 14332 29102
rect 14280 29038 14332 29044
rect 14096 28756 14148 28762
rect 14096 28698 14148 28704
rect 14016 28478 14504 28506
rect 14004 28416 14056 28422
rect 13924 28364 14004 28370
rect 13924 28358 14056 28364
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 13924 28342 14044 28358
rect 13912 27396 13964 27402
rect 13912 27338 13964 27344
rect 13924 26994 13952 27338
rect 13912 26988 13964 26994
rect 13912 26930 13964 26936
rect 13648 26438 13768 26466
rect 13544 25492 13596 25498
rect 13544 25434 13596 25440
rect 13648 24818 13676 26438
rect 13728 26308 13780 26314
rect 13728 26250 13780 26256
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13636 24404 13688 24410
rect 13636 24346 13688 24352
rect 13648 24070 13676 24346
rect 13636 24064 13688 24070
rect 13636 24006 13688 24012
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 12728 22066 12848 22094
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12624 19984 12676 19990
rect 12624 19926 12676 19932
rect 12636 18086 12664 19926
rect 12728 18902 12756 20334
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12820 18850 12848 22066
rect 13372 22066 13492 22094
rect 13372 22030 13400 22066
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 19378 13400 21830
rect 13452 21344 13504 21350
rect 13452 21286 13504 21292
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 12992 19304 13044 19310
rect 12990 19272 12992 19281
rect 13044 19272 13046 19281
rect 12990 19207 13046 19216
rect 13084 19236 13136 19242
rect 13268 19236 13320 19242
rect 13136 19196 13268 19224
rect 13084 19178 13136 19184
rect 13268 19178 13320 19184
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12820 18822 13308 18850
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12714 17912 12770 17921
rect 12714 17847 12770 17856
rect 12728 17814 12756 17847
rect 12716 17808 12768 17814
rect 12716 17750 12768 17756
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12636 16658 12664 16730
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12636 16402 12664 16594
rect 12728 16590 12756 17478
rect 12820 17270 12848 18634
rect 13280 18204 13308 18822
rect 13372 18714 13400 19314
rect 13464 18834 13492 21286
rect 13556 19378 13584 23122
rect 13636 22500 13688 22506
rect 13636 22442 13688 22448
rect 13648 21622 13676 22442
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13740 21486 13768 26250
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13832 24274 13860 24754
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13912 23792 13964 23798
rect 13912 23734 13964 23740
rect 13924 23118 13952 23734
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13832 21690 13860 22578
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13924 21690 13952 22510
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13648 20262 13676 20538
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13372 18686 13492 18714
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13372 18426 13400 18566
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13464 18204 13492 18686
rect 13280 18176 13400 18204
rect 13464 18176 13584 18204
rect 13372 18136 13400 18176
rect 13372 18108 13492 18136
rect 13268 18080 13320 18086
rect 13320 18040 13400 18068
rect 13268 18022 13320 18028
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12806 17912 12862 17921
rect 12950 17915 13258 17924
rect 13372 17354 13400 18040
rect 13280 17326 13400 17354
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 13280 17134 13308 17326
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 13372 17134 13400 17206
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 13464 16402 13492 18108
rect 12636 16374 12756 16402
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12452 16102 12572 16130
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12360 13530 12388 15846
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11900 12294 12296 12322
rect 11900 11778 11928 12294
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 11808 11750 11928 11778
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10152 800 10180 2382
rect 10520 800 10548 2926
rect 10888 800 10916 3470
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11256 3058 11284 3334
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11256 800 11284 2994
rect 11624 800 11652 4014
rect 11808 2650 11836 11750
rect 12084 10674 12112 12106
rect 12360 11898 12388 12378
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11900 3194 11928 8026
rect 12452 3534 12480 15574
rect 12544 12986 12572 16102
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12636 15502 12664 15846
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12636 15094 12664 15438
rect 12728 15366 12756 16374
rect 13372 16374 13492 16402
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11992 800 12020 2450
rect 12544 2446 12572 10474
rect 12636 6914 12664 14418
rect 12728 13394 12756 15302
rect 12820 14618 12848 16050
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13372 15144 13400 16374
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13464 15502 13492 16186
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13280 15116 13400 15144
rect 13280 14822 13308 15116
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 13372 14346 13400 14962
rect 13464 14482 13492 15030
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13360 14340 13412 14346
rect 13360 14282 13412 14288
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12728 8090 12756 12922
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11694 13216 12038
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13556 9654 13584 12702
rect 13832 12458 13860 17088
rect 13740 12430 13860 12458
rect 13740 9674 13768 12430
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13832 10810 13860 11834
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13648 9646 13768 9674
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12636 6886 12848 6914
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12636 3058 12664 4150
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12348 2372 12400 2378
rect 12348 2314 12400 2320
rect 12360 800 12388 2314
rect 12728 800 12756 3538
rect 12820 2582 12848 6886
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 13464 4146 13492 13806
rect 13556 12434 13584 18176
rect 13648 12850 13676 20198
rect 13832 20058 13860 21490
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13740 18970 13768 19654
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13740 18358 13768 18634
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13832 18193 13860 18838
rect 13818 18184 13874 18193
rect 13818 18119 13874 18128
rect 13832 14958 13860 18119
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13740 14074 13768 14758
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13740 13530 13768 14010
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 12442 13860 12786
rect 13820 12436 13872 12442
rect 13556 12406 13676 12434
rect 13648 10062 13676 12406
rect 13820 12378 13872 12384
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13924 9654 13952 20742
rect 14016 20602 14044 28342
rect 14188 27600 14240 27606
rect 14188 27542 14240 27548
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 14108 24138 14136 24686
rect 14096 24132 14148 24138
rect 14096 24074 14148 24080
rect 14200 22094 14228 27542
rect 14292 26382 14320 28358
rect 14372 26784 14424 26790
rect 14372 26726 14424 26732
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14384 25838 14412 26726
rect 14372 25832 14424 25838
rect 14372 25774 14424 25780
rect 14384 24750 14412 25774
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 14292 22098 14320 23122
rect 14108 22066 14228 22094
rect 14280 22092 14332 22098
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 14108 19378 14136 22066
rect 14280 22034 14332 22040
rect 14188 21956 14240 21962
rect 14188 21898 14240 21904
rect 14200 21486 14228 21898
rect 14476 21486 14504 28478
rect 14568 27470 14596 31726
rect 14660 31726 14780 31754
rect 14660 31142 14688 31726
rect 14832 31680 14884 31686
rect 14832 31622 14884 31628
rect 14648 31136 14700 31142
rect 14648 31078 14700 31084
rect 14660 29102 14688 31078
rect 14740 29572 14792 29578
rect 14740 29514 14792 29520
rect 14648 29096 14700 29102
rect 14648 29038 14700 29044
rect 14752 28762 14780 29514
rect 14740 28756 14792 28762
rect 14740 28698 14792 28704
rect 14740 28416 14792 28422
rect 14740 28358 14792 28364
rect 14752 27878 14780 28358
rect 14740 27872 14792 27878
rect 14740 27814 14792 27820
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14556 26988 14608 26994
rect 14556 26930 14608 26936
rect 14568 26246 14596 26930
rect 14556 26240 14608 26246
rect 14556 26182 14608 26188
rect 14568 25974 14596 26182
rect 14556 25968 14608 25974
rect 14556 25910 14608 25916
rect 14568 25770 14596 25910
rect 14556 25764 14608 25770
rect 14556 25706 14608 25712
rect 14752 23662 14780 27814
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14568 21962 14596 23258
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14200 19310 14228 19858
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14004 19236 14056 19242
rect 14004 19178 14056 19184
rect 14016 18902 14044 19178
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 14016 15978 14044 17682
rect 14200 17338 14228 18770
rect 14292 17746 14320 20878
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14188 17332 14240 17338
rect 14108 17292 14188 17320
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 14016 12306 14044 15914
rect 14108 15570 14136 17292
rect 14188 17274 14240 17280
rect 14292 16182 14320 17478
rect 14384 16726 14412 20742
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14280 16176 14332 16182
rect 14186 16144 14242 16153
rect 14280 16118 14332 16124
rect 14186 16079 14188 16088
rect 14240 16079 14242 16088
rect 14188 16050 14240 16056
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14108 15434 14136 15506
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14200 11762 14228 12106
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14292 11370 14320 15846
rect 14476 13410 14504 21082
rect 14844 20874 14872 31622
rect 15120 31414 15148 33050
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15108 31408 15160 31414
rect 15108 31350 15160 31356
rect 15212 30802 15240 32166
rect 15200 30796 15252 30802
rect 15200 30738 15252 30744
rect 15198 30424 15254 30433
rect 15198 30359 15254 30368
rect 14924 29708 14976 29714
rect 14924 29650 14976 29656
rect 14936 25838 14964 29650
rect 15108 29504 15160 29510
rect 15108 29446 15160 29452
rect 15016 27328 15068 27334
rect 15016 27270 15068 27276
rect 14924 25832 14976 25838
rect 14924 25774 14976 25780
rect 14924 25696 14976 25702
rect 14924 25638 14976 25644
rect 14936 22778 14964 25638
rect 15028 24818 15056 27270
rect 15120 27130 15148 29446
rect 15212 29102 15240 30359
rect 15200 29096 15252 29102
rect 15200 29038 15252 29044
rect 15212 28422 15240 29038
rect 15200 28416 15252 28422
rect 15198 28384 15200 28393
rect 15252 28384 15254 28393
rect 15198 28319 15254 28328
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 15212 27402 15240 28018
rect 15304 27946 15332 53926
rect 15396 43314 15424 53994
rect 15488 53582 15516 56200
rect 15476 53576 15528 53582
rect 15476 53518 15528 53524
rect 15856 53106 15884 56200
rect 16224 54330 16252 56200
rect 16212 54324 16264 54330
rect 16212 54266 16264 54272
rect 16592 53786 16620 56200
rect 16960 54194 16988 56200
rect 16948 54188 17000 54194
rect 16948 54130 17000 54136
rect 17040 53984 17092 53990
rect 17038 53952 17040 53961
rect 17092 53952 17094 53961
rect 17038 53887 17094 53896
rect 16580 53780 16632 53786
rect 16580 53722 16632 53728
rect 16592 53582 16620 53722
rect 17328 53582 17356 56200
rect 17696 54262 17724 56200
rect 18064 56114 18092 56200
rect 18156 56114 18184 56222
rect 18064 56086 18184 56114
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 17684 54256 17736 54262
rect 17684 54198 17736 54204
rect 18340 53582 18368 56222
rect 18418 56200 18474 57000
rect 18786 56200 18842 57000
rect 19154 56200 19210 57000
rect 19522 56200 19578 57000
rect 19890 56200 19946 57000
rect 20258 56200 20314 57000
rect 20626 56200 20682 57000
rect 20994 56200 21050 57000
rect 21362 56200 21418 57000
rect 21730 56200 21786 57000
rect 22098 56200 22154 57000
rect 22466 56200 22522 57000
rect 22834 56200 22890 57000
rect 23202 56200 23258 57000
rect 23570 56200 23626 57000
rect 18432 54126 18460 56200
rect 18420 54120 18472 54126
rect 18420 54062 18472 54068
rect 18512 53984 18564 53990
rect 18512 53926 18564 53932
rect 16580 53576 16632 53582
rect 16580 53518 16632 53524
rect 17316 53576 17368 53582
rect 17316 53518 17368 53524
rect 18328 53576 18380 53582
rect 18328 53518 18380 53524
rect 16396 53508 16448 53514
rect 16396 53450 16448 53456
rect 15844 53100 15896 53106
rect 15844 53042 15896 53048
rect 15936 52896 15988 52902
rect 15936 52838 15988 52844
rect 15844 50856 15896 50862
rect 15844 50798 15896 50804
rect 15660 44804 15712 44810
rect 15660 44746 15712 44752
rect 15476 43376 15528 43382
rect 15476 43318 15528 43324
rect 15384 43308 15436 43314
rect 15384 43250 15436 43256
rect 15396 43110 15424 43250
rect 15384 43104 15436 43110
rect 15384 43046 15436 43052
rect 15396 39386 15424 43046
rect 15488 40594 15516 43318
rect 15672 43246 15700 44746
rect 15660 43240 15712 43246
rect 15660 43182 15712 43188
rect 15568 40928 15620 40934
rect 15568 40870 15620 40876
rect 15476 40588 15528 40594
rect 15476 40530 15528 40536
rect 15580 39982 15608 40870
rect 15568 39976 15620 39982
rect 15568 39918 15620 39924
rect 15396 39358 15516 39386
rect 15384 39296 15436 39302
rect 15384 39238 15436 39244
rect 15396 36378 15424 39238
rect 15488 38758 15516 39358
rect 15476 38752 15528 38758
rect 15476 38694 15528 38700
rect 15476 38004 15528 38010
rect 15476 37946 15528 37952
rect 15488 37670 15516 37946
rect 15476 37664 15528 37670
rect 15476 37606 15528 37612
rect 15580 37466 15608 39918
rect 15672 39506 15700 43182
rect 15752 42220 15804 42226
rect 15752 42162 15804 42168
rect 15764 41750 15792 42162
rect 15752 41744 15804 41750
rect 15752 41686 15804 41692
rect 15856 40662 15884 50798
rect 15948 47802 15976 52838
rect 16408 52601 16436 53450
rect 16856 53440 16908 53446
rect 16856 53382 16908 53388
rect 16394 52592 16450 52601
rect 16394 52527 16450 52536
rect 16868 50862 16896 53382
rect 17328 53242 17356 53518
rect 17408 53440 17460 53446
rect 17408 53382 17460 53388
rect 18328 53440 18380 53446
rect 18328 53382 18380 53388
rect 17316 53236 17368 53242
rect 17316 53178 17368 53184
rect 16856 50856 16908 50862
rect 16856 50798 16908 50804
rect 17316 48272 17368 48278
rect 17316 48214 17368 48220
rect 17328 47802 17356 48214
rect 17420 47802 17448 53382
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 18340 53242 18368 53518
rect 17868 53236 17920 53242
rect 17868 53178 17920 53184
rect 18328 53236 18380 53242
rect 18328 53178 18380 53184
rect 18432 53174 18460 54198
rect 18616 54194 18644 56200
rect 18604 54188 18656 54194
rect 18604 54130 18656 54136
rect 18604 54052 18656 54058
rect 18604 53994 18656 54000
rect 18512 53440 18564 53446
rect 18512 53382 18564 53388
rect 18420 53168 18472 53174
rect 18420 53110 18472 53116
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17684 48272 17736 48278
rect 17684 48214 17736 48220
rect 15936 47796 15988 47802
rect 15936 47738 15988 47744
rect 17316 47796 17368 47802
rect 17316 47738 17368 47744
rect 17408 47796 17460 47802
rect 17408 47738 17460 47744
rect 16304 47524 16356 47530
rect 16304 47466 16356 47472
rect 16316 46374 16344 47466
rect 16580 47456 16632 47462
rect 16580 47398 16632 47404
rect 17500 47456 17552 47462
rect 17500 47398 17552 47404
rect 16396 46980 16448 46986
rect 16396 46922 16448 46928
rect 16304 46368 16356 46374
rect 16304 46310 16356 46316
rect 15936 45552 15988 45558
rect 15936 45494 15988 45500
rect 15948 45082 15976 45494
rect 16316 45422 16344 46310
rect 16408 45830 16436 46922
rect 16396 45824 16448 45830
rect 16396 45766 16448 45772
rect 16304 45416 16356 45422
rect 16304 45358 16356 45364
rect 16120 45280 16172 45286
rect 16120 45222 16172 45228
rect 15936 45076 15988 45082
rect 15936 45018 15988 45024
rect 15948 44810 15976 45018
rect 15936 44804 15988 44810
rect 15936 44746 15988 44752
rect 16028 43852 16080 43858
rect 16028 43794 16080 43800
rect 16040 41414 16068 43794
rect 16132 41682 16160 45222
rect 16396 42016 16448 42022
rect 16396 41958 16448 41964
rect 16408 41818 16436 41958
rect 16396 41812 16448 41818
rect 16396 41754 16448 41760
rect 16120 41676 16172 41682
rect 16120 41618 16172 41624
rect 16592 41596 16620 47398
rect 16672 47116 16724 47122
rect 16672 47058 16724 47064
rect 17224 47116 17276 47122
rect 17224 47058 17276 47064
rect 16684 47002 16712 47058
rect 16684 46974 16896 47002
rect 16868 46510 16896 46974
rect 16672 46504 16724 46510
rect 16672 46446 16724 46452
rect 16856 46504 16908 46510
rect 16856 46446 16908 46452
rect 16684 44742 16712 46446
rect 16764 45076 16816 45082
rect 16764 45018 16816 45024
rect 16672 44736 16724 44742
rect 16672 44678 16724 44684
rect 16776 43450 16804 45018
rect 16868 44946 16896 46446
rect 16856 44940 16908 44946
rect 16856 44882 16908 44888
rect 16868 44334 16896 44882
rect 16948 44736 17000 44742
rect 16948 44678 17000 44684
rect 16856 44328 16908 44334
rect 16856 44270 16908 44276
rect 16764 43444 16816 43450
rect 16764 43386 16816 43392
rect 16764 42560 16816 42566
rect 16764 42502 16816 42508
rect 16672 41608 16724 41614
rect 16592 41568 16672 41596
rect 16672 41550 16724 41556
rect 16488 41472 16540 41478
rect 16488 41414 16540 41420
rect 16040 41386 16160 41414
rect 15844 40656 15896 40662
rect 15844 40598 15896 40604
rect 15752 40588 15804 40594
rect 15752 40530 15804 40536
rect 15660 39500 15712 39506
rect 15660 39442 15712 39448
rect 15660 38888 15712 38894
rect 15660 38830 15712 38836
rect 15672 37806 15700 38830
rect 15660 37800 15712 37806
rect 15660 37742 15712 37748
rect 15568 37460 15620 37466
rect 15568 37402 15620 37408
rect 15568 37324 15620 37330
rect 15568 37266 15620 37272
rect 15384 36372 15436 36378
rect 15384 36314 15436 36320
rect 15580 35034 15608 37266
rect 15672 35290 15700 37742
rect 15764 36310 15792 40530
rect 15856 40497 15884 40598
rect 15842 40488 15898 40497
rect 15842 40423 15898 40432
rect 15844 40112 15896 40118
rect 15844 40054 15896 40060
rect 15856 37874 15884 40054
rect 16028 39976 16080 39982
rect 16028 39918 16080 39924
rect 16040 39574 16068 39918
rect 16028 39568 16080 39574
rect 16028 39510 16080 39516
rect 16040 39386 16068 39510
rect 15948 39358 16068 39386
rect 15948 39098 15976 39358
rect 16028 39296 16080 39302
rect 16028 39238 16080 39244
rect 16040 39098 16068 39238
rect 15936 39092 15988 39098
rect 15936 39034 15988 39040
rect 16028 39092 16080 39098
rect 16028 39034 16080 39040
rect 16132 38894 16160 41386
rect 16120 38888 16172 38894
rect 16120 38830 16172 38836
rect 16028 38752 16080 38758
rect 16026 38720 16028 38729
rect 16212 38752 16264 38758
rect 16080 38720 16082 38729
rect 16212 38694 16264 38700
rect 16026 38655 16082 38664
rect 15936 38344 15988 38350
rect 15936 38286 15988 38292
rect 15844 37868 15896 37874
rect 15844 37810 15896 37816
rect 15844 37120 15896 37126
rect 15844 37062 15896 37068
rect 15856 36854 15884 37062
rect 15844 36848 15896 36854
rect 15844 36790 15896 36796
rect 15844 36712 15896 36718
rect 15844 36654 15896 36660
rect 15856 36582 15884 36654
rect 15844 36576 15896 36582
rect 15844 36518 15896 36524
rect 15856 36378 15884 36518
rect 15844 36372 15896 36378
rect 15844 36314 15896 36320
rect 15752 36304 15804 36310
rect 15804 36252 15884 36258
rect 15752 36246 15884 36252
rect 15764 36230 15884 36246
rect 15856 36038 15884 36230
rect 15752 36032 15804 36038
rect 15750 36000 15752 36009
rect 15844 36032 15896 36038
rect 15804 36000 15806 36009
rect 15844 35974 15896 35980
rect 15750 35935 15806 35944
rect 15948 35494 15976 38286
rect 16120 37868 16172 37874
rect 16120 37810 16172 37816
rect 16028 37800 16080 37806
rect 16028 37742 16080 37748
rect 16040 36922 16068 37742
rect 16028 36916 16080 36922
rect 16028 36858 16080 36864
rect 15936 35488 15988 35494
rect 15936 35430 15988 35436
rect 15660 35284 15712 35290
rect 15660 35226 15712 35232
rect 15948 35170 15976 35430
rect 15764 35154 15976 35170
rect 15752 35148 15976 35154
rect 15804 35142 15976 35148
rect 15752 35090 15804 35096
rect 15580 35006 15792 35034
rect 15568 34944 15620 34950
rect 15568 34886 15620 34892
rect 15580 34610 15608 34886
rect 15568 34604 15620 34610
rect 15568 34546 15620 34552
rect 15476 32972 15528 32978
rect 15476 32914 15528 32920
rect 15382 29064 15438 29073
rect 15382 28999 15438 29008
rect 15292 27940 15344 27946
rect 15292 27882 15344 27888
rect 15396 27606 15424 28999
rect 15384 27600 15436 27606
rect 15384 27542 15436 27548
rect 15200 27396 15252 27402
rect 15200 27338 15252 27344
rect 15384 27396 15436 27402
rect 15384 27338 15436 27344
rect 15396 27305 15424 27338
rect 15382 27296 15438 27305
rect 15382 27231 15438 27240
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 15384 26376 15436 26382
rect 15384 26318 15436 26324
rect 15396 26042 15424 26318
rect 15384 26036 15436 26042
rect 15384 25978 15436 25984
rect 15396 25362 15424 25978
rect 15384 25356 15436 25362
rect 15384 25298 15436 25304
rect 15108 25152 15160 25158
rect 15108 25094 15160 25100
rect 15016 24812 15068 24818
rect 15016 24754 15068 24760
rect 15120 24682 15148 25094
rect 15396 24970 15424 25298
rect 15304 24942 15424 24970
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 15304 23186 15332 24942
rect 15488 24410 15516 32914
rect 15658 32872 15714 32881
rect 15658 32807 15714 32816
rect 15672 29306 15700 32807
rect 15660 29300 15712 29306
rect 15660 29242 15712 29248
rect 15568 29232 15620 29238
rect 15568 29174 15620 29180
rect 15580 28558 15608 29174
rect 15764 29073 15792 35006
rect 15844 34468 15896 34474
rect 15844 34410 15896 34416
rect 15856 33318 15884 34410
rect 15948 34066 15976 35142
rect 15936 34060 15988 34066
rect 15936 34002 15988 34008
rect 15948 33658 15976 34002
rect 15936 33652 15988 33658
rect 15936 33594 15988 33600
rect 15936 33516 15988 33522
rect 15936 33458 15988 33464
rect 15844 33312 15896 33318
rect 15844 33254 15896 33260
rect 15948 32434 15976 33458
rect 15936 32428 15988 32434
rect 15936 32370 15988 32376
rect 15948 31482 15976 32370
rect 15936 31476 15988 31482
rect 15936 31418 15988 31424
rect 15948 30938 15976 31418
rect 15936 30932 15988 30938
rect 15856 30892 15936 30920
rect 15856 30258 15884 30892
rect 15936 30874 15988 30880
rect 15844 30252 15896 30258
rect 15844 30194 15896 30200
rect 15750 29064 15806 29073
rect 15750 28999 15806 29008
rect 15568 28552 15620 28558
rect 15568 28494 15620 28500
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15660 28212 15712 28218
rect 15660 28154 15712 28160
rect 15568 27872 15620 27878
rect 15568 27814 15620 27820
rect 15580 26042 15608 27814
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 14924 22772 14976 22778
rect 14924 22714 14976 22720
rect 15488 22094 15516 24346
rect 15672 22710 15700 28154
rect 15660 22704 15712 22710
rect 15660 22646 15712 22652
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15396 22066 15516 22094
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 15120 20262 15148 21422
rect 15212 21078 15240 21490
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 15200 21072 15252 21078
rect 15200 21014 15252 21020
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14556 19304 14608 19310
rect 14554 19272 14556 19281
rect 14608 19272 14610 19281
rect 14554 19207 14610 19216
rect 14568 18834 14596 19207
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14752 17746 14780 19314
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14844 17746 14872 18770
rect 14936 18086 14964 19382
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 14844 17338 14872 17682
rect 14936 17678 14964 18022
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 14832 17332 14884 17338
rect 14752 17292 14832 17320
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14660 15502 14688 16390
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14568 14550 14596 14962
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14752 14482 14780 17292
rect 14832 17274 14884 17280
rect 15028 16998 15056 18226
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14384 13382 14504 13410
rect 14384 12918 14412 13382
rect 14844 13258 14872 14894
rect 14464 13252 14516 13258
rect 14832 13252 14884 13258
rect 14464 13194 14516 13200
rect 14568 13212 14832 13240
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14200 11342 14320 11370
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 14200 4214 14228 11342
rect 14384 6914 14412 12650
rect 14476 12442 14504 13194
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14568 11898 14596 13212
rect 14832 13194 14884 13200
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14292 6886 14412 6914
rect 14188 4208 14240 4214
rect 14188 4150 14240 4156
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 13096 870 13216 898
rect 13096 800 13124 870
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13188 762 13216 870
rect 13372 762 13400 2926
rect 13464 800 13492 3946
rect 14292 3058 14320 6886
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13832 800 13860 2314
rect 14200 800 14228 2926
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14568 800 14596 2450
rect 14660 2446 14688 12650
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14752 11218 14780 11698
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14936 6914 14964 12038
rect 15028 8974 15056 16934
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14844 6886 14964 6914
rect 14844 3126 14872 6886
rect 15120 5642 15148 20198
rect 15304 18222 15332 21286
rect 15396 20874 15424 22066
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15488 21350 15516 21422
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15476 20800 15528 20806
rect 15396 20748 15476 20754
rect 15396 20742 15528 20748
rect 15396 20726 15516 20742
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15396 17610 15424 20726
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15200 15904 15252 15910
rect 15396 15892 15424 17546
rect 15488 16046 15516 20198
rect 15580 17678 15608 22374
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15396 15864 15516 15892
rect 15200 15846 15252 15852
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15212 5250 15240 15846
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15304 12102 15332 14554
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15396 13394 15424 14418
rect 15488 14090 15516 15864
rect 15580 14278 15608 17478
rect 15672 15450 15700 22646
rect 15764 20942 15792 28358
rect 15856 28082 15884 30194
rect 16040 29850 16068 36858
rect 16132 34490 16160 37810
rect 16224 34678 16252 38694
rect 16304 38276 16356 38282
rect 16304 38218 16356 38224
rect 16316 37466 16344 38218
rect 16394 38176 16450 38185
rect 16394 38111 16450 38120
rect 16408 38010 16436 38111
rect 16396 38004 16448 38010
rect 16396 37946 16448 37952
rect 16304 37460 16356 37466
rect 16304 37402 16356 37408
rect 16500 37346 16528 41414
rect 16776 41070 16804 42502
rect 16764 41064 16816 41070
rect 16764 41006 16816 41012
rect 16960 40662 16988 44678
rect 17236 43246 17264 47058
rect 17408 43716 17460 43722
rect 17408 43658 17460 43664
rect 17224 43240 17276 43246
rect 17224 43182 17276 43188
rect 17040 43104 17092 43110
rect 17040 43046 17092 43052
rect 16948 40656 17000 40662
rect 16948 40598 17000 40604
rect 17052 40594 17080 43046
rect 17316 41812 17368 41818
rect 17316 41754 17368 41760
rect 17328 41478 17356 41754
rect 17316 41472 17368 41478
rect 17316 41414 17368 41420
rect 17040 40588 17092 40594
rect 17040 40530 17092 40536
rect 17040 40384 17092 40390
rect 17040 40326 17092 40332
rect 17316 40384 17368 40390
rect 17316 40326 17368 40332
rect 16948 40112 17000 40118
rect 16948 40054 17000 40060
rect 16856 38888 16908 38894
rect 16856 38830 16908 38836
rect 16580 38548 16632 38554
rect 16580 38490 16632 38496
rect 16408 37330 16528 37346
rect 16396 37324 16528 37330
rect 16448 37318 16528 37324
rect 16396 37266 16448 37272
rect 16304 37120 16356 37126
rect 16304 37062 16356 37068
rect 16212 34672 16264 34678
rect 16212 34614 16264 34620
rect 16132 34462 16252 34490
rect 16224 32774 16252 34462
rect 16316 34456 16344 37062
rect 16316 34428 16436 34456
rect 16304 33448 16356 33454
rect 16304 33390 16356 33396
rect 16120 32768 16172 32774
rect 16120 32710 16172 32716
rect 16212 32768 16264 32774
rect 16212 32710 16264 32716
rect 16132 32586 16160 32710
rect 16132 32570 16252 32586
rect 16132 32564 16264 32570
rect 16132 32558 16212 32564
rect 16212 32506 16264 32512
rect 16212 32360 16264 32366
rect 16212 32302 16264 32308
rect 16224 30190 16252 32302
rect 16316 32298 16344 33390
rect 16304 32292 16356 32298
rect 16304 32234 16356 32240
rect 16408 30326 16436 34428
rect 16592 31890 16620 38490
rect 16868 38010 16896 38830
rect 16856 38004 16908 38010
rect 16856 37946 16908 37952
rect 16960 37738 16988 40054
rect 17052 39642 17080 40326
rect 17132 40044 17184 40050
rect 17132 39986 17184 39992
rect 17040 39636 17092 39642
rect 17040 39578 17092 39584
rect 16764 37732 16816 37738
rect 16764 37674 16816 37680
rect 16948 37732 17000 37738
rect 16948 37674 17000 37680
rect 16776 37330 16804 37674
rect 17040 37392 17092 37398
rect 17040 37334 17092 37340
rect 16764 37324 16816 37330
rect 16764 37266 16816 37272
rect 17052 36922 17080 37334
rect 17040 36916 17092 36922
rect 17040 36858 17092 36864
rect 16762 36816 16818 36825
rect 16762 36751 16764 36760
rect 16816 36751 16818 36760
rect 16764 36722 16816 36728
rect 17144 35766 17172 39986
rect 17222 38312 17278 38321
rect 17222 38247 17278 38256
rect 17236 38214 17264 38247
rect 17224 38208 17276 38214
rect 17224 38150 17276 38156
rect 17224 36576 17276 36582
rect 17224 36518 17276 36524
rect 17132 35760 17184 35766
rect 17132 35702 17184 35708
rect 16948 32972 17000 32978
rect 16948 32914 17000 32920
rect 16856 32224 16908 32230
rect 16856 32166 16908 32172
rect 16580 31884 16632 31890
rect 16580 31826 16632 31832
rect 16764 31680 16816 31686
rect 16764 31622 16816 31628
rect 16488 31204 16540 31210
rect 16488 31146 16540 31152
rect 16500 30433 16528 31146
rect 16580 30660 16632 30666
rect 16580 30602 16632 30608
rect 16486 30424 16542 30433
rect 16486 30359 16542 30368
rect 16396 30320 16448 30326
rect 16396 30262 16448 30268
rect 16212 30184 16264 30190
rect 16212 30126 16264 30132
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 16028 29028 16080 29034
rect 16028 28970 16080 28976
rect 16040 28558 16068 28970
rect 16120 28960 16172 28966
rect 16120 28902 16172 28908
rect 16028 28552 16080 28558
rect 16028 28494 16080 28500
rect 15934 28248 15990 28257
rect 15934 28183 15936 28192
rect 15988 28183 15990 28192
rect 15936 28154 15988 28160
rect 16132 28150 16160 28902
rect 16224 28626 16252 30126
rect 16592 29850 16620 30602
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16580 29844 16632 29850
rect 16580 29786 16632 29792
rect 16396 29572 16448 29578
rect 16396 29514 16448 29520
rect 16304 29232 16356 29238
rect 16304 29174 16356 29180
rect 16212 28620 16264 28626
rect 16212 28562 16264 28568
rect 16120 28144 16172 28150
rect 16120 28086 16172 28092
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 15844 27600 15896 27606
rect 15844 27542 15896 27548
rect 15856 27334 15884 27542
rect 15844 27328 15896 27334
rect 15844 27270 15896 27276
rect 15948 25480 15976 28018
rect 16028 28008 16080 28014
rect 16028 27950 16080 27956
rect 16040 27878 16068 27950
rect 16028 27872 16080 27878
rect 16028 27814 16080 27820
rect 16212 27600 16264 27606
rect 16212 27542 16264 27548
rect 16028 25832 16080 25838
rect 16028 25774 16080 25780
rect 15856 25452 15976 25480
rect 15856 22982 15884 25452
rect 16040 23322 16068 25774
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 15936 23044 15988 23050
rect 15936 22986 15988 22992
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15856 22506 15884 22918
rect 15948 22574 15976 22986
rect 15936 22568 15988 22574
rect 15988 22516 16160 22522
rect 15936 22510 16160 22516
rect 15844 22500 15896 22506
rect 15948 22494 16160 22510
rect 15844 22442 15896 22448
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15856 18834 15884 22442
rect 16028 22228 16080 22234
rect 16028 22170 16080 22176
rect 16040 21962 16068 22170
rect 16132 22098 16160 22494
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16028 21956 16080 21962
rect 16028 21898 16080 21904
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15948 20754 15976 21830
rect 16026 20768 16082 20777
rect 15948 20726 16026 20754
rect 16026 20703 16082 20712
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15948 16658 15976 18158
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15764 16114 15792 16594
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15672 15422 15792 15450
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15488 14062 15608 14090
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15120 5222 15240 5250
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14832 3120 14884 3126
rect 14832 3062 14884 3068
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14936 800 14964 3538
rect 15120 3534 15148 5222
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15304 800 15332 2450
rect 15396 2310 15424 12038
rect 15488 11354 15516 13126
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15580 9654 15608 14062
rect 15672 12442 15700 15302
rect 15764 12986 15792 15422
rect 15948 14906 15976 16594
rect 16040 15026 16068 20703
rect 16224 18850 16252 27542
rect 16316 22094 16344 29174
rect 16408 29170 16436 29514
rect 16396 29164 16448 29170
rect 16396 29106 16448 29112
rect 16408 29073 16436 29106
rect 16394 29064 16450 29073
rect 16394 28999 16450 29008
rect 16396 27872 16448 27878
rect 16396 27814 16448 27820
rect 16408 23338 16436 27814
rect 16500 23594 16528 29786
rect 16592 24750 16620 29786
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16684 25362 16712 26522
rect 16776 26518 16804 31622
rect 16868 28558 16896 32166
rect 16960 31686 16988 32914
rect 17236 32434 17264 36518
rect 17224 32428 17276 32434
rect 17224 32370 17276 32376
rect 17328 31754 17356 40326
rect 17420 33114 17448 43658
rect 17512 43450 17540 47398
rect 17592 46912 17644 46918
rect 17592 46854 17644 46860
rect 17604 46646 17632 46854
rect 17592 46640 17644 46646
rect 17592 46582 17644 46588
rect 17604 45830 17632 46582
rect 17592 45824 17644 45830
rect 17592 45766 17644 45772
rect 17604 45082 17632 45766
rect 17592 45076 17644 45082
rect 17592 45018 17644 45024
rect 17604 44470 17632 45018
rect 17592 44464 17644 44470
rect 17592 44406 17644 44412
rect 17592 43648 17644 43654
rect 17592 43590 17644 43596
rect 17500 43444 17552 43450
rect 17500 43386 17552 43392
rect 17604 43382 17632 43590
rect 17592 43376 17644 43382
rect 17592 43318 17644 43324
rect 17500 41608 17552 41614
rect 17500 41550 17552 41556
rect 17512 36242 17540 41550
rect 17696 41414 17724 48214
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 18340 47734 18368 53382
rect 18524 48278 18552 53926
rect 18800 53106 18828 56200
rect 18880 54256 18932 54262
rect 18880 54198 18932 54204
rect 18892 53786 18920 54198
rect 18880 53780 18932 53786
rect 18880 53722 18932 53728
rect 19168 53582 19196 56200
rect 19536 54194 19564 56200
rect 19524 54188 19576 54194
rect 19524 54130 19576 54136
rect 19708 54120 19760 54126
rect 19708 54062 19760 54068
rect 19340 53984 19392 53990
rect 19340 53926 19392 53932
rect 19156 53576 19208 53582
rect 19156 53518 19208 53524
rect 19168 53242 19196 53518
rect 19156 53236 19208 53242
rect 19156 53178 19208 53184
rect 18788 53100 18840 53106
rect 18788 53042 18840 53048
rect 18604 52896 18656 52902
rect 18604 52838 18656 52844
rect 18512 48272 18564 48278
rect 18512 48214 18564 48220
rect 18328 47728 18380 47734
rect 18328 47670 18380 47676
rect 18512 47184 18564 47190
rect 18512 47126 18564 47132
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 18328 45416 18380 45422
rect 18328 45358 18380 45364
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 18340 44198 18368 45358
rect 18328 44192 18380 44198
rect 18328 44134 18380 44140
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 18340 43246 18368 44134
rect 18328 43240 18380 43246
rect 18328 43182 18380 43188
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 18328 42016 18380 42022
rect 18328 41958 18380 41964
rect 18340 41546 18368 41958
rect 18524 41682 18552 47126
rect 18616 47122 18644 52838
rect 18788 47728 18840 47734
rect 18786 47696 18788 47705
rect 18840 47696 18842 47705
rect 18786 47631 18842 47640
rect 18696 47592 18748 47598
rect 18696 47534 18748 47540
rect 18708 47258 18736 47534
rect 19352 47258 19380 53926
rect 19616 53440 19668 53446
rect 19616 53382 19668 53388
rect 18696 47252 18748 47258
rect 18696 47194 18748 47200
rect 19340 47252 19392 47258
rect 19340 47194 19392 47200
rect 18604 47116 18656 47122
rect 18604 47058 18656 47064
rect 18604 46980 18656 46986
rect 18604 46922 18656 46928
rect 18616 43722 18644 46922
rect 18708 46714 18736 47194
rect 19340 47116 19392 47122
rect 19340 47058 19392 47064
rect 18696 46708 18748 46714
rect 18696 46650 18748 46656
rect 18972 46708 19024 46714
rect 18972 46650 19024 46656
rect 18788 46504 18840 46510
rect 18788 46446 18840 46452
rect 18800 44198 18828 46446
rect 18984 44334 19012 46650
rect 19352 46510 19380 47058
rect 19340 46504 19392 46510
rect 19340 46446 19392 46452
rect 19064 45824 19116 45830
rect 19064 45766 19116 45772
rect 18972 44328 19024 44334
rect 18972 44270 19024 44276
rect 18788 44192 18840 44198
rect 18788 44134 18840 44140
rect 18604 43716 18656 43722
rect 18604 43658 18656 43664
rect 18512 41676 18564 41682
rect 18512 41618 18564 41624
rect 18328 41540 18380 41546
rect 18328 41482 18380 41488
rect 17604 41386 17724 41414
rect 17604 39409 17632 41386
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17684 40452 17736 40458
rect 17684 40394 17736 40400
rect 17590 39400 17646 39409
rect 17590 39335 17646 39344
rect 17604 38729 17632 39335
rect 17590 38720 17646 38729
rect 17590 38655 17646 38664
rect 17590 38584 17646 38593
rect 17590 38519 17646 38528
rect 17604 37806 17632 38519
rect 17592 37800 17644 37806
rect 17592 37742 17644 37748
rect 17500 36236 17552 36242
rect 17500 36178 17552 36184
rect 17408 33108 17460 33114
rect 17408 33050 17460 33056
rect 17696 32570 17724 40394
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17868 39500 17920 39506
rect 17868 39442 17920 39448
rect 17776 39024 17828 39030
rect 17776 38966 17828 38972
rect 17788 38554 17816 38966
rect 17776 38548 17828 38554
rect 17776 38490 17828 38496
rect 17776 38344 17828 38350
rect 17776 38286 17828 38292
rect 17788 37398 17816 38286
rect 17880 38214 17908 39442
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 18236 38752 18288 38758
rect 18236 38694 18288 38700
rect 18248 38418 18276 38694
rect 18236 38412 18288 38418
rect 18236 38354 18288 38360
rect 17868 38208 17920 38214
rect 17868 38150 17920 38156
rect 17776 37392 17828 37398
rect 17776 37334 17828 37340
rect 17776 37256 17828 37262
rect 17774 37224 17776 37233
rect 17828 37224 17830 37233
rect 17774 37159 17830 37168
rect 17776 36848 17828 36854
rect 17776 36790 17828 36796
rect 17788 35834 17816 36790
rect 17776 35828 17828 35834
rect 17776 35770 17828 35776
rect 17880 35766 17908 38150
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 18340 37738 18368 41482
rect 18420 41472 18472 41478
rect 18472 41432 18552 41460
rect 18420 41414 18472 41420
rect 18420 41200 18472 41206
rect 18420 41142 18472 41148
rect 18432 40934 18460 41142
rect 18420 40928 18472 40934
rect 18420 40870 18472 40876
rect 18432 39828 18460 40870
rect 18524 39982 18552 41432
rect 18604 41132 18656 41138
rect 18604 41074 18656 41080
rect 18616 40730 18644 41074
rect 18696 40928 18748 40934
rect 18696 40870 18748 40876
rect 18604 40724 18656 40730
rect 18604 40666 18656 40672
rect 18512 39976 18564 39982
rect 18512 39918 18564 39924
rect 18432 39800 18552 39828
rect 18420 39296 18472 39302
rect 18420 39238 18472 39244
rect 18432 38894 18460 39238
rect 18420 38888 18472 38894
rect 18418 38856 18420 38865
rect 18472 38856 18474 38865
rect 18418 38791 18474 38800
rect 18524 38654 18552 39800
rect 18616 39506 18644 40666
rect 18604 39500 18656 39506
rect 18604 39442 18656 39448
rect 18604 39364 18656 39370
rect 18604 39306 18656 39312
rect 18432 38626 18552 38654
rect 18432 38282 18460 38626
rect 18616 38486 18644 39306
rect 18708 38758 18736 40870
rect 18800 39982 18828 44134
rect 18984 41682 19012 44270
rect 18972 41676 19024 41682
rect 18972 41618 19024 41624
rect 18880 41472 18932 41478
rect 18880 41414 18932 41420
rect 18892 40934 18920 41414
rect 18880 40928 18932 40934
rect 18880 40870 18932 40876
rect 18892 40594 18920 40870
rect 18880 40588 18932 40594
rect 18880 40530 18932 40536
rect 18892 40390 18920 40530
rect 18880 40384 18932 40390
rect 18880 40326 18932 40332
rect 18788 39976 18840 39982
rect 18788 39918 18840 39924
rect 18788 39500 18840 39506
rect 18788 39442 18840 39448
rect 18696 38752 18748 38758
rect 18696 38694 18748 38700
rect 18604 38480 18656 38486
rect 18604 38422 18656 38428
rect 18420 38276 18472 38282
rect 18420 38218 18472 38224
rect 18432 38010 18460 38218
rect 18512 38208 18564 38214
rect 18512 38150 18564 38156
rect 18420 38004 18472 38010
rect 18420 37946 18472 37952
rect 18328 37732 18380 37738
rect 18328 37674 18380 37680
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 18432 35766 18460 37946
rect 18524 37466 18552 38150
rect 18604 37936 18656 37942
rect 18604 37878 18656 37884
rect 18512 37460 18564 37466
rect 18512 37402 18564 37408
rect 18512 37120 18564 37126
rect 18512 37062 18564 37068
rect 18524 36922 18552 37062
rect 18512 36916 18564 36922
rect 18512 36858 18564 36864
rect 17868 35760 17920 35766
rect 18420 35760 18472 35766
rect 17868 35702 17920 35708
rect 18340 35720 18420 35748
rect 17960 35488 18012 35494
rect 17960 35430 18012 35436
rect 17868 35284 17920 35290
rect 17868 35226 17920 35232
rect 17776 34060 17828 34066
rect 17776 34002 17828 34008
rect 17684 32564 17736 32570
rect 17684 32506 17736 32512
rect 17684 32224 17736 32230
rect 17684 32166 17736 32172
rect 17052 31726 17356 31754
rect 17592 31748 17644 31754
rect 16948 31680 17000 31686
rect 16948 31622 17000 31628
rect 16960 30802 16988 31622
rect 16948 30796 17000 30802
rect 16948 30738 17000 30744
rect 16948 30388 17000 30394
rect 16948 30330 17000 30336
rect 16960 29034 16988 30330
rect 17052 29646 17080 31726
rect 17592 31690 17644 31696
rect 17604 31482 17632 31690
rect 17592 31476 17644 31482
rect 17592 31418 17644 31424
rect 17132 31136 17184 31142
rect 17132 31078 17184 31084
rect 17040 29640 17092 29646
rect 17040 29582 17092 29588
rect 16948 29028 17000 29034
rect 16948 28970 17000 28976
rect 16856 28552 16908 28558
rect 16856 28494 16908 28500
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16764 26512 16816 26518
rect 16764 26454 16816 26460
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16776 24206 16804 25434
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 16868 24954 16896 25094
rect 16856 24948 16908 24954
rect 16856 24890 16908 24896
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16868 24410 16896 24754
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16488 23588 16540 23594
rect 16488 23530 16540 23536
rect 16500 23474 16528 23530
rect 16500 23446 16620 23474
rect 16408 23310 16528 23338
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16408 22982 16436 23054
rect 16396 22976 16448 22982
rect 16396 22918 16448 22924
rect 16408 22778 16436 22918
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16408 22234 16436 22714
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16316 22066 16436 22094
rect 16132 18822 16252 18850
rect 16132 15502 16160 18822
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16224 18222 16252 18702
rect 16304 18352 16356 18358
rect 16304 18294 16356 18300
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16316 16454 16344 18294
rect 16408 17746 16436 22066
rect 16500 18358 16528 23310
rect 16592 22778 16620 23446
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16592 21146 16620 22578
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16592 20806 16620 21082
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16488 18352 16540 18358
rect 16488 18294 16540 18300
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16394 16280 16450 16289
rect 16394 16215 16396 16224
rect 16448 16215 16450 16224
rect 16396 16186 16448 16192
rect 16304 16108 16356 16114
rect 16500 16096 16528 18158
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 16998 16620 17478
rect 16684 17202 16712 24006
rect 16868 22642 16896 24346
rect 16960 24274 16988 28358
rect 17052 28098 17080 29582
rect 17144 28626 17172 31078
rect 17408 30252 17460 30258
rect 17408 30194 17460 30200
rect 17224 30184 17276 30190
rect 17224 30126 17276 30132
rect 17236 29306 17264 30126
rect 17316 29776 17368 29782
rect 17316 29718 17368 29724
rect 17224 29300 17276 29306
rect 17224 29242 17276 29248
rect 17132 28620 17184 28626
rect 17132 28562 17184 28568
rect 17052 28070 17172 28098
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 17052 24274 17080 25094
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 17040 24268 17092 24274
rect 17040 24210 17092 24216
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 17052 22030 17080 23598
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 16764 20868 16816 20874
rect 16764 20810 16816 20816
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16580 16108 16632 16114
rect 16500 16068 16580 16096
rect 16304 16050 16356 16056
rect 16580 16050 16632 16056
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 16132 14958 16160 15438
rect 16120 14952 16172 14958
rect 15948 14878 16068 14906
rect 16120 14894 16172 14900
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15948 13530 15976 14282
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15948 12850 15976 13466
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15660 12436 15712 12442
rect 16040 12434 16068 14878
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 16040 12406 16160 12434
rect 15660 12378 15712 12384
rect 16132 12306 16160 12406
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 15672 11218 15700 12242
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15764 10674 15792 11494
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15948 3942 15976 11086
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 16132 3670 16160 4082
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 15672 800 15700 2926
rect 16040 800 16068 3538
rect 16224 3534 16252 12650
rect 16316 6914 16344 16050
rect 16592 14498 16620 16050
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16684 15094 16712 15302
rect 16776 15094 16804 20810
rect 17040 20324 17092 20330
rect 17040 20266 17092 20272
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16868 16402 16896 20198
rect 17052 19378 17080 20266
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 17144 19174 17172 28070
rect 17222 27432 17278 27441
rect 17222 27367 17224 27376
rect 17276 27367 17278 27376
rect 17224 27338 17276 27344
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17236 26790 17264 26930
rect 17224 26784 17276 26790
rect 17224 26726 17276 26732
rect 17236 26353 17264 26726
rect 17222 26344 17278 26353
rect 17222 26279 17278 26288
rect 17224 26240 17276 26246
rect 17224 26182 17276 26188
rect 17236 25770 17264 26182
rect 17224 25764 17276 25770
rect 17224 25706 17276 25712
rect 17236 25294 17264 25706
rect 17224 25288 17276 25294
rect 17224 25230 17276 25236
rect 17328 24206 17356 29718
rect 17420 29102 17448 30194
rect 17592 30048 17644 30054
rect 17592 29990 17644 29996
rect 17604 29782 17632 29990
rect 17592 29776 17644 29782
rect 17592 29718 17644 29724
rect 17592 29572 17644 29578
rect 17592 29514 17644 29520
rect 17500 29504 17552 29510
rect 17500 29446 17552 29452
rect 17512 29306 17540 29446
rect 17604 29306 17632 29514
rect 17500 29300 17552 29306
rect 17500 29242 17552 29248
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17696 29186 17724 32166
rect 17788 31278 17816 34002
rect 17880 33998 17908 35226
rect 17972 35154 18000 35430
rect 18340 35290 18368 35720
rect 18420 35702 18472 35708
rect 18616 35630 18644 37878
rect 18696 37868 18748 37874
rect 18696 37810 18748 37816
rect 18708 37777 18736 37810
rect 18694 37768 18750 37777
rect 18694 37703 18750 37712
rect 18800 37448 18828 39442
rect 18878 38584 18934 38593
rect 18984 38570 19012 41618
rect 18934 38542 19012 38570
rect 18878 38519 18934 38528
rect 18880 38480 18932 38486
rect 18880 38422 18932 38428
rect 18892 37942 18920 38422
rect 18880 37936 18932 37942
rect 18880 37878 18932 37884
rect 18880 37732 18932 37738
rect 18880 37674 18932 37680
rect 18708 37420 18828 37448
rect 18604 35624 18656 35630
rect 18604 35566 18656 35572
rect 18328 35284 18380 35290
rect 18328 35226 18380 35232
rect 18420 35284 18472 35290
rect 18420 35226 18472 35232
rect 17960 35148 18012 35154
rect 17960 35090 18012 35096
rect 18328 35148 18380 35154
rect 18328 35090 18380 35096
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17868 33992 17920 33998
rect 17868 33934 17920 33940
rect 17880 33658 17908 33934
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 17868 33652 17920 33658
rect 17868 33594 17920 33600
rect 17880 33046 17908 33594
rect 18340 33590 18368 35090
rect 18432 34202 18460 35226
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 18420 34196 18472 34202
rect 18420 34138 18472 34144
rect 18328 33584 18380 33590
rect 18328 33526 18380 33532
rect 17868 33040 17920 33046
rect 17868 32982 17920 32988
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 17868 32360 17920 32366
rect 17868 32302 17920 32308
rect 17776 31272 17828 31278
rect 17776 31214 17828 31220
rect 17512 29158 17724 29186
rect 17408 29096 17460 29102
rect 17408 29038 17460 29044
rect 17408 26852 17460 26858
rect 17408 26794 17460 26800
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 17420 21554 17448 26794
rect 17512 25906 17540 29158
rect 17788 29102 17816 31214
rect 17880 30598 17908 32302
rect 18420 31884 18472 31890
rect 18420 31826 18472 31832
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 18328 31340 18380 31346
rect 18328 31282 18380 31288
rect 17868 30592 17920 30598
rect 17868 30534 17920 30540
rect 17880 30258 17908 30534
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18340 30394 18368 31282
rect 18328 30388 18380 30394
rect 18328 30330 18380 30336
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 18328 30116 18380 30122
rect 18328 30058 18380 30064
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 18340 29238 18368 30058
rect 18328 29232 18380 29238
rect 18328 29174 18380 29180
rect 17592 29096 17644 29102
rect 17592 29038 17644 29044
rect 17776 29096 17828 29102
rect 17776 29038 17828 29044
rect 17604 26450 17632 29038
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 17788 26586 17816 28562
rect 18326 28520 18382 28529
rect 18326 28455 18382 28464
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 18340 28218 18368 28455
rect 18432 28422 18460 31826
rect 18524 31482 18552 34546
rect 18616 32230 18644 35566
rect 18708 32502 18736 37420
rect 18892 37398 18920 37674
rect 18880 37392 18932 37398
rect 18786 37360 18842 37369
rect 18880 37334 18932 37340
rect 18786 37295 18842 37304
rect 18800 34082 18828 37295
rect 18880 36712 18932 36718
rect 18880 36654 18932 36660
rect 18970 36680 19026 36689
rect 18892 34218 18920 36654
rect 18970 36615 18972 36624
rect 19024 36615 19026 36624
rect 18972 36586 19024 36592
rect 18892 34190 19012 34218
rect 18800 34054 18920 34082
rect 18696 32496 18748 32502
rect 18696 32438 18748 32444
rect 18696 32360 18748 32366
rect 18696 32302 18748 32308
rect 18604 32224 18656 32230
rect 18604 32166 18656 32172
rect 18512 31476 18564 31482
rect 18512 31418 18564 31424
rect 18604 30932 18656 30938
rect 18604 30874 18656 30880
rect 18512 30660 18564 30666
rect 18512 30602 18564 30608
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18328 28212 18380 28218
rect 18328 28154 18380 28160
rect 18340 27674 18368 28154
rect 18328 27668 18380 27674
rect 18328 27610 18380 27616
rect 17868 27532 17920 27538
rect 17868 27474 17920 27480
rect 17776 26580 17828 26586
rect 17776 26522 17828 26528
rect 17592 26444 17644 26450
rect 17592 26386 17644 26392
rect 17500 25900 17552 25906
rect 17500 25842 17552 25848
rect 17604 25786 17632 26386
rect 17880 25922 17908 27474
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 18432 27062 18460 28358
rect 18524 28150 18552 30602
rect 18616 28558 18644 30874
rect 18708 30666 18736 32302
rect 18892 31822 18920 34054
rect 18984 31822 19012 34190
rect 18880 31816 18932 31822
rect 18880 31758 18932 31764
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 18788 31680 18840 31686
rect 18788 31622 18840 31628
rect 18696 30660 18748 30666
rect 18696 30602 18748 30608
rect 18696 30388 18748 30394
rect 18696 30330 18748 30336
rect 18604 28552 18656 28558
rect 18604 28494 18656 28500
rect 18512 28144 18564 28150
rect 18512 28086 18564 28092
rect 18512 28008 18564 28014
rect 18512 27950 18564 27956
rect 18420 27056 18472 27062
rect 18420 26998 18472 27004
rect 18420 26512 18472 26518
rect 18420 26454 18472 26460
rect 18326 26344 18382 26353
rect 18326 26279 18382 26288
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 17512 25758 17632 25786
rect 17788 25894 17908 25922
rect 17512 24750 17540 25758
rect 17788 24954 17816 25894
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 18236 25832 18288 25838
rect 18236 25774 18288 25780
rect 17880 25158 17908 25774
rect 18248 25498 18276 25774
rect 18236 25492 18288 25498
rect 18236 25434 18288 25440
rect 18340 25294 18368 26279
rect 18328 25288 18380 25294
rect 18328 25230 18380 25236
rect 17868 25152 17920 25158
rect 17868 25094 17920 25100
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 18340 24954 18368 25230
rect 17776 24948 17828 24954
rect 17776 24890 17828 24896
rect 18328 24948 18380 24954
rect 18328 24890 18380 24896
rect 18432 24818 18460 26454
rect 18524 25480 18552 27950
rect 18604 27328 18656 27334
rect 18604 27270 18656 27276
rect 18616 27062 18644 27270
rect 18604 27056 18656 27062
rect 18604 26998 18656 27004
rect 18524 25452 18644 25480
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18616 24750 18644 25452
rect 18708 24750 18736 30330
rect 18800 29714 18828 31622
rect 18788 29708 18840 29714
rect 18788 29650 18840 29656
rect 18800 28150 18828 29650
rect 18788 28144 18840 28150
rect 18788 28086 18840 28092
rect 18788 27668 18840 27674
rect 18788 27610 18840 27616
rect 17500 24744 17552 24750
rect 17500 24686 17552 24692
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 17512 24138 17540 24686
rect 17684 24676 17736 24682
rect 17684 24618 17736 24624
rect 17500 24132 17552 24138
rect 17500 24074 17552 24080
rect 17512 23866 17540 24074
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17314 20632 17370 20641
rect 17314 20567 17316 20576
rect 17368 20567 17370 20576
rect 17316 20538 17368 20544
rect 17316 19780 17368 19786
rect 17316 19722 17368 19728
rect 17328 19514 17356 19722
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 16868 16374 16988 16402
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 16856 14884 16908 14890
rect 16856 14826 16908 14832
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16408 14482 16620 14498
rect 16396 14476 16620 14482
rect 16448 14470 16620 14476
rect 16396 14418 16448 14424
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16408 11778 16436 14214
rect 16500 13258 16528 14214
rect 16592 13938 16620 14470
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16500 12986 16528 13194
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16500 11898 16528 12922
rect 16488 11892 16540 11898
rect 16684 11880 16712 14758
rect 16488 11834 16540 11840
rect 16592 11852 16712 11880
rect 16408 11750 16528 11778
rect 16316 6886 16436 6914
rect 16408 6390 16436 6886
rect 16500 6798 16528 11750
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16396 6384 16448 6390
rect 16396 6326 16448 6332
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16316 3641 16344 3946
rect 16302 3632 16358 3641
rect 16302 3567 16358 3576
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16408 800 16436 4014
rect 16592 3670 16620 11852
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16684 4146 16712 11290
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16776 3058 16804 11494
rect 16868 11354 16896 14826
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16776 800 16804 2790
rect 16868 2446 16896 9862
rect 16960 3058 16988 16374
rect 17144 16182 17172 17682
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17052 12918 17080 15098
rect 17144 14618 17172 16118
rect 17236 15706 17264 19450
rect 17512 18358 17540 22714
rect 17592 21480 17644 21486
rect 17592 21422 17644 21428
rect 17604 20942 17632 21422
rect 17696 20942 17724 24618
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18420 24132 18472 24138
rect 18420 24074 18472 24080
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 17788 21010 17816 21422
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 17774 19952 17830 19961
rect 17880 19922 17908 24006
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17960 23792 18012 23798
rect 17958 23760 17960 23769
rect 18012 23760 18014 23769
rect 17958 23695 18014 23704
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18432 22166 18460 24074
rect 18420 22160 18472 22166
rect 18420 22102 18472 22108
rect 18524 22098 18552 24550
rect 18616 24138 18644 24686
rect 18604 24132 18656 24138
rect 18604 24074 18656 24080
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18616 23186 18644 23598
rect 18604 23180 18656 23186
rect 18604 23122 18656 23128
rect 18616 22710 18644 23122
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 18512 22092 18564 22098
rect 18512 22034 18564 22040
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18696 21412 18748 21418
rect 18696 21354 18748 21360
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 17774 19887 17830 19896
rect 17868 19916 17920 19922
rect 17788 19854 17816 19887
rect 17868 19858 17920 19864
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17788 18970 17816 19110
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 18326 18728 18382 18737
rect 18326 18663 18382 18672
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18340 18426 18368 18663
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17512 17882 17540 18294
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17972 16998 18000 17206
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 17144 12306 17172 13874
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17236 12986 17264 13126
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17328 12170 17356 16934
rect 17972 16504 18000 16934
rect 17880 16476 18000 16504
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17420 14006 17448 15506
rect 17512 14890 17540 16390
rect 17880 16182 17908 16476
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17868 16176 17920 16182
rect 17920 16136 18092 16164
rect 17868 16118 17920 16124
rect 18064 16096 18092 16136
rect 18144 16108 18196 16114
rect 18064 16068 18144 16096
rect 18144 16050 18196 16056
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17408 14000 17460 14006
rect 17460 13960 17540 13988
rect 17408 13942 17460 13948
rect 17512 12442 17540 13960
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17328 7478 17356 12106
rect 17420 11694 17448 12378
rect 17498 11928 17554 11937
rect 17498 11863 17500 11872
rect 17552 11863 17554 11872
rect 17500 11834 17552 11840
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17604 11150 17632 14010
rect 18340 13462 18368 18362
rect 18328 13456 18380 13462
rect 18328 13398 18380 13404
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17696 10742 17724 12582
rect 17684 10736 17736 10742
rect 17684 10678 17736 10684
rect 17788 10606 17816 13126
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18340 12102 18368 13194
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18432 11898 18460 12786
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18248 10130 18276 10406
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18432 9994 18460 20198
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18524 18902 18552 19654
rect 18512 18896 18564 18902
rect 18512 18838 18564 18844
rect 18524 14906 18552 18838
rect 18708 17134 18736 21354
rect 18800 19990 18828 27610
rect 18892 25786 18920 31758
rect 18972 31680 19024 31686
rect 18972 31622 19024 31628
rect 18984 28014 19012 31622
rect 19076 31278 19104 45766
rect 19352 45626 19380 46446
rect 19524 46368 19576 46374
rect 19524 46310 19576 46316
rect 19340 45620 19392 45626
rect 19340 45562 19392 45568
rect 19536 44878 19564 46310
rect 19628 45898 19656 53382
rect 19720 53242 19748 54062
rect 19904 53582 19932 56200
rect 19892 53576 19944 53582
rect 19892 53518 19944 53524
rect 19708 53236 19760 53242
rect 19708 53178 19760 53184
rect 20272 53106 20300 56200
rect 20640 55214 20668 56200
rect 20640 55186 20760 55214
rect 20732 54194 20760 55186
rect 20720 54188 20772 54194
rect 20720 54130 20772 54136
rect 20444 53508 20496 53514
rect 20444 53450 20496 53456
rect 20260 53100 20312 53106
rect 20260 53042 20312 53048
rect 20168 52896 20220 52902
rect 20168 52838 20220 52844
rect 20180 46034 20208 52838
rect 20456 47258 20484 53450
rect 20732 53174 20760 54130
rect 20904 53984 20956 53990
rect 20904 53926 20956 53932
rect 20720 53168 20772 53174
rect 20720 53110 20772 53116
rect 20444 47252 20496 47258
rect 20444 47194 20496 47200
rect 20456 47161 20484 47194
rect 20442 47152 20498 47161
rect 20442 47087 20498 47096
rect 20536 46504 20588 46510
rect 20536 46446 20588 46452
rect 20168 46028 20220 46034
rect 20168 45970 20220 45976
rect 20444 46028 20496 46034
rect 20444 45970 20496 45976
rect 19616 45892 19668 45898
rect 19616 45834 19668 45840
rect 19892 45824 19944 45830
rect 19892 45766 19944 45772
rect 19524 44872 19576 44878
rect 19524 44814 19576 44820
rect 19536 44334 19564 44814
rect 19800 44804 19852 44810
rect 19800 44746 19852 44752
rect 19812 44538 19840 44746
rect 19800 44532 19852 44538
rect 19800 44474 19852 44480
rect 19524 44328 19576 44334
rect 19524 44270 19576 44276
rect 19524 43648 19576 43654
rect 19524 43590 19576 43596
rect 19248 43104 19300 43110
rect 19248 43046 19300 43052
rect 19156 42560 19208 42566
rect 19156 42502 19208 42508
rect 19168 38962 19196 42502
rect 19260 42158 19288 43046
rect 19248 42152 19300 42158
rect 19248 42094 19300 42100
rect 19260 41682 19288 42094
rect 19340 41744 19392 41750
rect 19340 41686 19392 41692
rect 19248 41676 19300 41682
rect 19248 41618 19300 41624
rect 19260 41274 19288 41618
rect 19248 41268 19300 41274
rect 19248 41210 19300 41216
rect 19248 39840 19300 39846
rect 19248 39782 19300 39788
rect 19156 38956 19208 38962
rect 19156 38898 19208 38904
rect 19156 38820 19208 38826
rect 19156 38762 19208 38768
rect 19168 38554 19196 38762
rect 19156 38548 19208 38554
rect 19156 38490 19208 38496
rect 19260 35698 19288 39782
rect 19352 38554 19380 41686
rect 19432 40928 19484 40934
rect 19432 40870 19484 40876
rect 19444 39506 19472 40870
rect 19536 39982 19564 43590
rect 19708 43172 19760 43178
rect 19708 43114 19760 43120
rect 19616 42356 19668 42362
rect 19616 42298 19668 42304
rect 19524 39976 19576 39982
rect 19524 39918 19576 39924
rect 19432 39500 19484 39506
rect 19432 39442 19484 39448
rect 19524 39296 19576 39302
rect 19524 39238 19576 39244
rect 19340 38548 19392 38554
rect 19340 38490 19392 38496
rect 19430 38448 19486 38457
rect 19430 38383 19432 38392
rect 19484 38383 19486 38392
rect 19432 38354 19484 38360
rect 19340 38208 19392 38214
rect 19340 38150 19392 38156
rect 19248 35692 19300 35698
rect 19248 35634 19300 35640
rect 19248 33856 19300 33862
rect 19248 33798 19300 33804
rect 19156 31680 19208 31686
rect 19156 31622 19208 31628
rect 19064 31272 19116 31278
rect 19064 31214 19116 31220
rect 19062 30288 19118 30297
rect 19062 30223 19064 30232
rect 19116 30223 19118 30232
rect 19064 30194 19116 30200
rect 19076 30054 19104 30194
rect 19064 30048 19116 30054
rect 19064 29990 19116 29996
rect 19064 29504 19116 29510
rect 19064 29446 19116 29452
rect 19076 29034 19104 29446
rect 19064 29028 19116 29034
rect 19064 28970 19116 28976
rect 19076 28014 19104 28970
rect 18972 28008 19024 28014
rect 18972 27950 19024 27956
rect 19064 28008 19116 28014
rect 19064 27950 19116 27956
rect 18972 27872 19024 27878
rect 18972 27814 19024 27820
rect 19064 27872 19116 27878
rect 19064 27814 19116 27820
rect 18984 26450 19012 27814
rect 18972 26444 19024 26450
rect 18972 26386 19024 26392
rect 18892 25758 19012 25786
rect 18880 25696 18932 25702
rect 18880 25638 18932 25644
rect 18788 19984 18840 19990
rect 18788 19926 18840 19932
rect 18892 19854 18920 25638
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18788 19780 18840 19786
rect 18788 19722 18840 19728
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18616 16250 18644 17070
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18616 15026 18644 16186
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18708 15162 18736 15302
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18524 14878 18736 14906
rect 18602 14512 18658 14521
rect 18602 14447 18658 14456
rect 18616 14414 18644 14447
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18524 13938 18552 14214
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18524 12986 18552 13330
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18524 11830 18552 12922
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17684 9444 17736 9450
rect 17684 9386 17736 9392
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17144 800 17172 2858
rect 17512 800 17540 4014
rect 17696 2514 17724 9386
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18524 6914 18552 13126
rect 18708 12434 18736 17054
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18616 12406 18736 12434
rect 18616 8974 18644 12406
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18800 7886 18828 16730
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18524 6886 18644 6914
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18432 6322 18460 8298
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17788 4758 17816 5170
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 18524 4622 18552 6598
rect 18616 4622 18644 12582
rect 18708 9654 18736 14878
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18800 6914 18828 19722
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18892 18086 18920 19110
rect 18984 18970 19012 25758
rect 19076 25362 19104 27814
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 18984 18766 19012 18906
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18892 17762 18920 18022
rect 18984 17898 19012 18566
rect 19076 18204 19104 21286
rect 19168 20466 19196 31622
rect 19260 30938 19288 33798
rect 19248 30932 19300 30938
rect 19248 30874 19300 30880
rect 19248 30048 19300 30054
rect 19248 29990 19300 29996
rect 19260 27554 19288 29990
rect 19352 29578 19380 38150
rect 19430 38040 19486 38049
rect 19430 37975 19486 37984
rect 19444 36310 19472 37975
rect 19432 36304 19484 36310
rect 19432 36246 19484 36252
rect 19432 34196 19484 34202
rect 19432 34138 19484 34144
rect 19444 33998 19472 34138
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 19432 33380 19484 33386
rect 19432 33322 19484 33328
rect 19444 31754 19472 33322
rect 19536 32366 19564 39238
rect 19628 36922 19656 42298
rect 19720 41070 19748 43114
rect 19800 42628 19852 42634
rect 19800 42570 19852 42576
rect 19708 41064 19760 41070
rect 19708 41006 19760 41012
rect 19812 40662 19840 42570
rect 19904 41206 19932 45766
rect 20076 45416 20128 45422
rect 20076 45358 20128 45364
rect 20088 43450 20116 45358
rect 20456 44538 20484 45970
rect 20548 45558 20576 46446
rect 20916 45966 20944 53926
rect 21008 53582 21036 56200
rect 21376 54194 21404 56200
rect 21364 54188 21416 54194
rect 21364 54130 21416 54136
rect 21548 53984 21600 53990
rect 21548 53926 21600 53932
rect 20996 53576 21048 53582
rect 20996 53518 21048 53524
rect 21008 53242 21036 53518
rect 21364 53440 21416 53446
rect 21364 53382 21416 53388
rect 20996 53236 21048 53242
rect 20996 53178 21048 53184
rect 20996 49972 21048 49978
rect 20996 49914 21048 49920
rect 20904 45960 20956 45966
rect 20904 45902 20956 45908
rect 20720 45824 20772 45830
rect 20720 45766 20772 45772
rect 20536 45552 20588 45558
rect 20536 45494 20588 45500
rect 20548 45286 20576 45494
rect 20536 45280 20588 45286
rect 20536 45222 20588 45228
rect 20548 44946 20576 45222
rect 20536 44940 20588 44946
rect 20536 44882 20588 44888
rect 20444 44532 20496 44538
rect 20444 44474 20496 44480
rect 20548 44470 20576 44882
rect 20628 44736 20680 44742
rect 20628 44678 20680 44684
rect 20260 44464 20312 44470
rect 20536 44464 20588 44470
rect 20312 44412 20536 44418
rect 20260 44406 20588 44412
rect 20272 44390 20576 44406
rect 20076 43444 20128 43450
rect 20076 43386 20128 43392
rect 19984 42152 20036 42158
rect 19984 42094 20036 42100
rect 19996 41546 20024 42094
rect 19984 41540 20036 41546
rect 19984 41482 20036 41488
rect 19892 41200 19944 41206
rect 19892 41142 19944 41148
rect 19984 41064 20036 41070
rect 19984 41006 20036 41012
rect 19800 40656 19852 40662
rect 19800 40598 19852 40604
rect 19800 39976 19852 39982
rect 19800 39918 19852 39924
rect 19708 38004 19760 38010
rect 19708 37946 19760 37952
rect 19720 37806 19748 37946
rect 19708 37800 19760 37806
rect 19708 37742 19760 37748
rect 19706 37224 19762 37233
rect 19706 37159 19762 37168
rect 19616 36916 19668 36922
rect 19616 36858 19668 36864
rect 19720 36281 19748 37159
rect 19812 36666 19840 39918
rect 19892 38956 19944 38962
rect 19892 38898 19944 38904
rect 19904 38282 19932 38898
rect 19892 38276 19944 38282
rect 19892 38218 19944 38224
rect 19904 36854 19932 38218
rect 19892 36848 19944 36854
rect 19892 36790 19944 36796
rect 19996 36786 20024 41006
rect 20088 39506 20116 43386
rect 20548 43382 20576 44390
rect 20536 43376 20588 43382
rect 20536 43318 20588 43324
rect 20548 43110 20576 43318
rect 20640 43246 20668 44678
rect 20628 43240 20680 43246
rect 20628 43182 20680 43188
rect 20536 43104 20588 43110
rect 20536 43046 20588 43052
rect 20352 42900 20404 42906
rect 20352 42842 20404 42848
rect 20260 42016 20312 42022
rect 20260 41958 20312 41964
rect 20168 41268 20220 41274
rect 20168 41210 20220 41216
rect 20180 40458 20208 41210
rect 20168 40452 20220 40458
rect 20168 40394 20220 40400
rect 20076 39500 20128 39506
rect 20076 39442 20128 39448
rect 20168 38548 20220 38554
rect 20168 38490 20220 38496
rect 20180 37874 20208 38490
rect 20272 38418 20300 41958
rect 20364 39982 20392 42842
rect 20548 42634 20576 43046
rect 20536 42628 20588 42634
rect 20536 42570 20588 42576
rect 20732 42362 20760 45766
rect 20916 45554 20944 45902
rect 20824 45526 20944 45554
rect 20824 45286 20852 45526
rect 20812 45280 20864 45286
rect 20812 45222 20864 45228
rect 20824 44305 20852 45222
rect 20810 44296 20866 44305
rect 20810 44231 20866 44240
rect 20812 43648 20864 43654
rect 20812 43590 20864 43596
rect 20720 42356 20772 42362
rect 20720 42298 20772 42304
rect 20628 42220 20680 42226
rect 20628 42162 20680 42168
rect 20536 40656 20588 40662
rect 20536 40598 20588 40604
rect 20548 40361 20576 40598
rect 20534 40352 20590 40361
rect 20534 40287 20590 40296
rect 20352 39976 20404 39982
rect 20352 39918 20404 39924
rect 20352 39432 20404 39438
rect 20352 39374 20404 39380
rect 20442 39400 20498 39409
rect 20260 38412 20312 38418
rect 20260 38354 20312 38360
rect 20364 38010 20392 39374
rect 20442 39335 20444 39344
rect 20496 39335 20498 39344
rect 20444 39306 20496 39312
rect 20456 38894 20484 39306
rect 20444 38888 20496 38894
rect 20444 38830 20496 38836
rect 20444 38276 20496 38282
rect 20444 38218 20496 38224
rect 20456 38185 20484 38218
rect 20442 38176 20498 38185
rect 20442 38111 20498 38120
rect 20352 38004 20404 38010
rect 20352 37946 20404 37952
rect 20258 37904 20314 37913
rect 20168 37868 20220 37874
rect 20456 37890 20484 38111
rect 20258 37839 20260 37848
rect 20168 37810 20220 37816
rect 20312 37839 20314 37848
rect 20364 37862 20484 37890
rect 20260 37810 20312 37816
rect 20364 37670 20392 37862
rect 20444 37800 20496 37806
rect 20444 37742 20496 37748
rect 20352 37664 20404 37670
rect 20352 37606 20404 37612
rect 20456 37369 20484 37742
rect 20442 37360 20498 37369
rect 20442 37295 20444 37304
rect 20496 37295 20498 37304
rect 20444 37266 20496 37272
rect 20076 37188 20128 37194
rect 20076 37130 20128 37136
rect 20168 37188 20220 37194
rect 20168 37130 20220 37136
rect 19984 36780 20036 36786
rect 19984 36722 20036 36728
rect 19812 36638 19932 36666
rect 19706 36272 19762 36281
rect 19706 36207 19762 36216
rect 19616 35012 19668 35018
rect 19616 34954 19668 34960
rect 19628 33658 19656 34954
rect 19720 33998 19748 36207
rect 19800 35488 19852 35494
rect 19800 35430 19852 35436
rect 19812 34746 19840 35430
rect 19800 34740 19852 34746
rect 19800 34682 19852 34688
rect 19800 34468 19852 34474
rect 19800 34410 19852 34416
rect 19708 33992 19760 33998
rect 19708 33934 19760 33940
rect 19616 33652 19668 33658
rect 19616 33594 19668 33600
rect 19524 32360 19576 32366
rect 19524 32302 19576 32308
rect 19628 31890 19656 33594
rect 19616 31884 19668 31890
rect 19616 31826 19668 31832
rect 19444 31726 19656 31754
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19340 29572 19392 29578
rect 19340 29514 19392 29520
rect 19260 27526 19380 27554
rect 19352 27282 19380 27526
rect 19260 27254 19380 27282
rect 19260 24857 19288 27254
rect 19340 26920 19392 26926
rect 19340 26862 19392 26868
rect 19352 26042 19380 26862
rect 19340 26036 19392 26042
rect 19340 25978 19392 25984
rect 19444 25294 19472 30534
rect 19522 29336 19578 29345
rect 19522 29271 19524 29280
rect 19576 29271 19578 29280
rect 19524 29242 19576 29248
rect 19628 29034 19656 31726
rect 19812 30190 19840 34410
rect 19904 33386 19932 36638
rect 20088 36582 20116 37130
rect 20076 36576 20128 36582
rect 20076 36518 20128 36524
rect 20088 33930 20116 36518
rect 20180 35154 20208 37130
rect 20352 36032 20404 36038
rect 20352 35974 20404 35980
rect 20444 36032 20496 36038
rect 20444 35974 20496 35980
rect 20168 35148 20220 35154
rect 20168 35090 20220 35096
rect 20260 34672 20312 34678
rect 20260 34614 20312 34620
rect 20272 34134 20300 34614
rect 20260 34128 20312 34134
rect 20260 34070 20312 34076
rect 20076 33924 20128 33930
rect 20076 33866 20128 33872
rect 19892 33380 19944 33386
rect 19892 33322 19944 33328
rect 20076 32224 20128 32230
rect 20076 32166 20128 32172
rect 19892 31408 19944 31414
rect 19892 31350 19944 31356
rect 19904 31142 19932 31350
rect 19984 31272 20036 31278
rect 19982 31240 19984 31249
rect 20036 31240 20038 31249
rect 19982 31175 20038 31184
rect 19892 31136 19944 31142
rect 19892 31078 19944 31084
rect 19984 30796 20036 30802
rect 19984 30738 20036 30744
rect 19800 30184 19852 30190
rect 19800 30126 19852 30132
rect 19616 29028 19668 29034
rect 19616 28970 19668 28976
rect 19812 28490 19840 30126
rect 19800 28484 19852 28490
rect 19800 28426 19852 28432
rect 19524 28076 19576 28082
rect 19524 28018 19576 28024
rect 19536 27402 19564 28018
rect 19616 28008 19668 28014
rect 19616 27950 19668 27956
rect 19524 27396 19576 27402
rect 19524 27338 19576 27344
rect 19524 26784 19576 26790
rect 19524 26726 19576 26732
rect 19536 26042 19564 26726
rect 19524 26036 19576 26042
rect 19524 25978 19576 25984
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19524 25152 19576 25158
rect 19524 25094 19576 25100
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 19246 24848 19302 24857
rect 19246 24783 19302 24792
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19260 19446 19288 22374
rect 19352 22030 19380 24890
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19444 23050 19472 23258
rect 19432 23044 19484 23050
rect 19432 22986 19484 22992
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 19352 20602 19380 21014
rect 19444 21010 19472 21966
rect 19432 21004 19484 21010
rect 19432 20946 19484 20952
rect 19536 20602 19564 25094
rect 19628 24954 19656 27950
rect 19812 26926 19840 28426
rect 19996 28014 20024 30738
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19800 26920 19852 26926
rect 19800 26862 19852 26868
rect 19708 26512 19760 26518
rect 19708 26454 19760 26460
rect 19616 24948 19668 24954
rect 19616 24890 19668 24896
rect 19720 22710 19748 26454
rect 19892 24132 19944 24138
rect 19892 24074 19944 24080
rect 19800 23656 19852 23662
rect 19800 23598 19852 23604
rect 19708 22704 19760 22710
rect 19708 22646 19760 22652
rect 19616 22636 19668 22642
rect 19616 22578 19668 22584
rect 19628 21894 19656 22578
rect 19812 22574 19840 23598
rect 19904 22930 19932 24074
rect 19996 23050 20024 27950
rect 20088 25974 20116 32166
rect 20168 30796 20220 30802
rect 20168 30738 20220 30744
rect 20180 29102 20208 30738
rect 20272 30734 20300 34070
rect 20260 30728 20312 30734
rect 20260 30670 20312 30676
rect 20364 30410 20392 35974
rect 20456 31822 20484 35974
rect 20548 35766 20576 40287
rect 20640 40186 20668 42162
rect 20720 41064 20772 41070
rect 20720 41006 20772 41012
rect 20628 40180 20680 40186
rect 20628 40122 20680 40128
rect 20732 39098 20760 41006
rect 20720 39092 20772 39098
rect 20720 39034 20772 39040
rect 20628 38208 20680 38214
rect 20628 38150 20680 38156
rect 20536 35760 20588 35766
rect 20536 35702 20588 35708
rect 20640 34610 20668 38150
rect 20720 37460 20772 37466
rect 20720 37402 20772 37408
rect 20732 37194 20760 37402
rect 20720 37188 20772 37194
rect 20720 37130 20772 37136
rect 20732 34746 20760 37130
rect 20720 34740 20772 34746
rect 20720 34682 20772 34688
rect 20628 34604 20680 34610
rect 20628 34546 20680 34552
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20536 34128 20588 34134
rect 20536 34070 20588 34076
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 20548 31754 20576 34070
rect 20628 33856 20680 33862
rect 20628 33798 20680 33804
rect 20640 33658 20668 33798
rect 20628 33652 20680 33658
rect 20628 33594 20680 33600
rect 20536 31748 20588 31754
rect 20536 31690 20588 31696
rect 20628 31680 20680 31686
rect 20628 31622 20680 31628
rect 20536 31272 20588 31278
rect 20536 31214 20588 31220
rect 20442 30968 20498 30977
rect 20442 30903 20444 30912
rect 20496 30903 20498 30912
rect 20444 30874 20496 30880
rect 20364 30394 20484 30410
rect 20364 30388 20496 30394
rect 20364 30382 20444 30388
rect 20444 30330 20496 30336
rect 20352 29504 20404 29510
rect 20352 29446 20404 29452
rect 20168 29096 20220 29102
rect 20168 29038 20220 29044
rect 20076 25968 20128 25974
rect 20076 25910 20128 25916
rect 20076 25356 20128 25362
rect 20076 25298 20128 25304
rect 20088 23322 20116 25298
rect 20180 24682 20208 29038
rect 20258 28248 20314 28257
rect 20258 28183 20260 28192
rect 20312 28183 20314 28192
rect 20260 28154 20312 28160
rect 20260 26444 20312 26450
rect 20260 26386 20312 26392
rect 20168 24676 20220 24682
rect 20168 24618 20220 24624
rect 20272 24070 20300 26386
rect 20364 26042 20392 29446
rect 20456 27470 20484 30330
rect 20548 27538 20576 31214
rect 20536 27532 20588 27538
rect 20536 27474 20588 27480
rect 20444 27464 20496 27470
rect 20444 27406 20496 27412
rect 20548 26858 20576 27474
rect 20536 26852 20588 26858
rect 20536 26794 20588 26800
rect 20640 26314 20668 31622
rect 20732 29646 20760 34342
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20824 29306 20852 43590
rect 20904 43104 20956 43110
rect 20904 43046 20956 43052
rect 20916 42362 20944 43046
rect 20904 42356 20956 42362
rect 20904 42298 20956 42304
rect 20916 41682 20944 42298
rect 20904 41676 20956 41682
rect 20904 41618 20956 41624
rect 21008 41070 21036 49914
rect 21376 46034 21404 53382
rect 21560 49314 21588 53926
rect 21640 53712 21692 53718
rect 21640 53654 21692 53660
rect 21652 49450 21680 53654
rect 21744 53582 21772 56200
rect 22112 53582 22140 56200
rect 22480 54194 22508 56200
rect 22468 54188 22520 54194
rect 22468 54130 22520 54136
rect 22480 54074 22508 54130
rect 22480 54046 22600 54074
rect 22192 53984 22244 53990
rect 22192 53926 22244 53932
rect 21732 53576 21784 53582
rect 21732 53518 21784 53524
rect 22100 53576 22152 53582
rect 22100 53518 22152 53524
rect 21744 53242 21772 53518
rect 22112 53242 22140 53518
rect 21732 53236 21784 53242
rect 21732 53178 21784 53184
rect 22100 53236 22152 53242
rect 22100 53178 22152 53184
rect 22204 52986 22232 53926
rect 22376 53712 22428 53718
rect 22376 53654 22428 53660
rect 22112 52958 22232 52986
rect 21652 49422 21772 49450
rect 21560 49286 21680 49314
rect 21364 46028 21416 46034
rect 21364 45970 21416 45976
rect 21548 46028 21600 46034
rect 21548 45970 21600 45976
rect 21560 45558 21588 45970
rect 21548 45552 21600 45558
rect 21548 45494 21600 45500
rect 21456 44940 21508 44946
rect 21456 44882 21508 44888
rect 21468 44538 21496 44882
rect 21456 44532 21508 44538
rect 21456 44474 21508 44480
rect 21180 44328 21232 44334
rect 21180 44270 21232 44276
rect 21192 41818 21220 44270
rect 21560 42906 21588 45494
rect 21652 43314 21680 49286
rect 21744 43722 21772 49422
rect 22008 46912 22060 46918
rect 22008 46854 22060 46860
rect 21916 46708 21968 46714
rect 21916 46650 21968 46656
rect 21928 46617 21956 46650
rect 21914 46608 21970 46617
rect 21914 46543 21970 46552
rect 21732 43716 21784 43722
rect 21732 43658 21784 43664
rect 21916 43648 21968 43654
rect 21916 43590 21968 43596
rect 21640 43308 21692 43314
rect 21640 43250 21692 43256
rect 21652 43110 21680 43250
rect 21640 43104 21692 43110
rect 21638 43072 21640 43081
rect 21692 43072 21694 43081
rect 21638 43007 21694 43016
rect 21548 42900 21600 42906
rect 21548 42842 21600 42848
rect 21272 42560 21324 42566
rect 21272 42502 21324 42508
rect 21824 42560 21876 42566
rect 21824 42502 21876 42508
rect 21284 42158 21312 42502
rect 21272 42152 21324 42158
rect 21272 42094 21324 42100
rect 21180 41812 21232 41818
rect 21180 41754 21232 41760
rect 21088 41540 21140 41546
rect 21088 41482 21140 41488
rect 21100 41274 21128 41482
rect 21088 41268 21140 41274
rect 21088 41210 21140 41216
rect 21088 41132 21140 41138
rect 21088 41074 21140 41080
rect 20996 41064 21048 41070
rect 20996 41006 21048 41012
rect 21100 40934 21128 41074
rect 20904 40928 20956 40934
rect 20904 40870 20956 40876
rect 21088 40928 21140 40934
rect 21088 40870 21140 40876
rect 20916 39030 20944 40870
rect 20996 40384 21048 40390
rect 20996 40326 21048 40332
rect 21008 40118 21036 40326
rect 20996 40112 21048 40118
rect 20996 40054 21048 40060
rect 21008 39302 21036 40054
rect 20996 39296 21048 39302
rect 20996 39238 21048 39244
rect 20904 39024 20956 39030
rect 20904 38966 20956 38972
rect 20904 38888 20956 38894
rect 20904 38830 20956 38836
rect 20916 35290 20944 38830
rect 20996 38208 21048 38214
rect 20996 38150 21048 38156
rect 21008 36310 21036 38150
rect 20996 36304 21048 36310
rect 20996 36246 21048 36252
rect 21100 36038 21128 40870
rect 21192 38418 21220 41754
rect 21548 41268 21600 41274
rect 21548 41210 21600 41216
rect 21454 40624 21510 40633
rect 21364 40588 21416 40594
rect 21454 40559 21456 40568
rect 21364 40530 21416 40536
rect 21508 40559 21510 40568
rect 21456 40530 21508 40536
rect 21376 40497 21404 40530
rect 21362 40488 21418 40497
rect 21362 40423 21418 40432
rect 21456 40452 21508 40458
rect 21456 40394 21508 40400
rect 21468 40186 21496 40394
rect 21456 40180 21508 40186
rect 21456 40122 21508 40128
rect 21364 39500 21416 39506
rect 21364 39442 21416 39448
rect 21272 38752 21324 38758
rect 21272 38694 21324 38700
rect 21180 38412 21232 38418
rect 21180 38354 21232 38360
rect 21284 36242 21312 38694
rect 21376 37806 21404 39442
rect 21468 38554 21496 40122
rect 21456 38548 21508 38554
rect 21456 38490 21508 38496
rect 21364 37800 21416 37806
rect 21364 37742 21416 37748
rect 21272 36236 21324 36242
rect 21272 36178 21324 36184
rect 21180 36168 21232 36174
rect 21180 36110 21232 36116
rect 21088 36032 21140 36038
rect 21088 35974 21140 35980
rect 21088 35692 21140 35698
rect 21088 35634 21140 35640
rect 20996 35488 21048 35494
rect 20996 35430 21048 35436
rect 20904 35284 20956 35290
rect 20904 35226 20956 35232
rect 21008 35018 21036 35430
rect 21100 35290 21128 35634
rect 21088 35284 21140 35290
rect 21088 35226 21140 35232
rect 20996 35012 21048 35018
rect 20996 34954 21048 34960
rect 21192 34950 21220 36110
rect 21180 34944 21232 34950
rect 21180 34886 21232 34892
rect 21192 34066 21220 34886
rect 21180 34060 21232 34066
rect 21180 34002 21232 34008
rect 20904 33924 20956 33930
rect 20904 33866 20956 33872
rect 20916 33114 20944 33866
rect 20996 33448 21048 33454
rect 20996 33390 21048 33396
rect 20904 33108 20956 33114
rect 20904 33050 20956 33056
rect 21008 32910 21036 33390
rect 21192 33318 21220 34002
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 21284 33318 21312 33458
rect 21376 33318 21404 37742
rect 21560 37738 21588 41210
rect 21836 40497 21864 42502
rect 21638 40488 21694 40497
rect 21638 40423 21640 40432
rect 21692 40423 21694 40432
rect 21822 40488 21878 40497
rect 21822 40423 21878 40432
rect 21640 40394 21692 40400
rect 21732 38820 21784 38826
rect 21732 38762 21784 38768
rect 21640 38548 21692 38554
rect 21640 38490 21692 38496
rect 21652 38350 21680 38490
rect 21640 38344 21692 38350
rect 21640 38286 21692 38292
rect 21548 37732 21600 37738
rect 21548 37674 21600 37680
rect 21548 35556 21600 35562
rect 21548 35498 21600 35504
rect 21456 33856 21508 33862
rect 21456 33798 21508 33804
rect 21468 33658 21496 33798
rect 21456 33652 21508 33658
rect 21456 33594 21508 33600
rect 21180 33312 21232 33318
rect 21180 33254 21232 33260
rect 21272 33312 21324 33318
rect 21272 33254 21324 33260
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21180 33108 21232 33114
rect 21180 33050 21232 33056
rect 20996 32904 21048 32910
rect 20996 32846 21048 32852
rect 20904 32768 20956 32774
rect 21088 32768 21140 32774
rect 20904 32710 20956 32716
rect 21008 32716 21088 32722
rect 21008 32710 21140 32716
rect 20916 31686 20944 32710
rect 21008 32694 21128 32710
rect 20904 31680 20956 31686
rect 20904 31622 20956 31628
rect 20904 29504 20956 29510
rect 20904 29446 20956 29452
rect 20916 29306 20944 29446
rect 20812 29300 20864 29306
rect 20812 29242 20864 29248
rect 20904 29300 20956 29306
rect 20904 29242 20956 29248
rect 20824 29186 20852 29242
rect 20824 29158 20944 29186
rect 20916 29034 20944 29158
rect 20812 29028 20864 29034
rect 20812 28970 20864 28976
rect 20904 29028 20956 29034
rect 20904 28970 20956 28976
rect 20628 26308 20680 26314
rect 20628 26250 20680 26256
rect 20352 26036 20404 26042
rect 20352 25978 20404 25984
rect 20720 24744 20772 24750
rect 20720 24686 20772 24692
rect 20628 24676 20680 24682
rect 20628 24618 20680 24624
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 20180 23202 20208 23462
rect 20088 23174 20208 23202
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 19904 22902 20024 22930
rect 19800 22568 19852 22574
rect 19800 22510 19852 22516
rect 19812 22094 19840 22510
rect 19812 22066 19932 22094
rect 19904 21894 19932 22066
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 19996 21554 20024 22902
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19982 21176 20038 21185
rect 19982 21111 19984 21120
rect 20036 21111 20038 21120
rect 19984 21082 20036 21088
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 19352 19394 19380 19654
rect 19444 19514 19472 19654
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19536 19394 19564 19450
rect 19352 19366 19564 19394
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19156 18216 19208 18222
rect 19076 18176 19156 18204
rect 19156 18158 19208 18164
rect 18984 17870 19196 17898
rect 18892 17734 19012 17762
rect 18880 17604 18932 17610
rect 18880 17546 18932 17552
rect 18892 15162 18920 17546
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18892 12918 18920 13398
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18984 12434 19012 17734
rect 19168 13870 19196 17870
rect 19260 16250 19288 19178
rect 19352 18426 19380 19246
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19352 17134 19380 18362
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19168 13462 19196 13806
rect 19156 13456 19208 13462
rect 19156 13398 19208 13404
rect 18892 12406 19012 12434
rect 18892 8566 18920 12406
rect 19352 12238 19380 14758
rect 19444 14550 19472 19366
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19536 17338 19564 17614
rect 19524 17332 19576 17338
rect 19524 17274 19576 17280
rect 19536 16522 19564 17274
rect 19524 16516 19576 16522
rect 19524 16458 19576 16464
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19536 14414 19564 16458
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19444 13326 19472 14214
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19536 12782 19564 14350
rect 19628 14074 19656 15302
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19536 11898 19564 12718
rect 19720 12434 19748 18566
rect 19812 15026 19840 20198
rect 20088 16538 20116 23174
rect 20272 22234 20300 24006
rect 20640 23798 20668 24618
rect 20732 23866 20760 24686
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20628 23792 20680 23798
rect 20628 23734 20680 23740
rect 20444 23316 20496 23322
rect 20444 23258 20496 23264
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20180 20874 20208 21422
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20272 21162 20300 21354
rect 20364 21332 20392 22714
rect 20456 21486 20484 23258
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 20444 21344 20496 21350
rect 20364 21304 20444 21332
rect 20444 21286 20496 21292
rect 20272 21134 20392 21162
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20180 17610 20208 18022
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 20180 16658 20208 17546
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 19996 16510 20116 16538
rect 19996 15638 20024 16510
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20088 16250 20116 16390
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 19892 15632 19944 15638
rect 19892 15574 19944 15580
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19904 13394 19932 15574
rect 19996 15502 20024 15574
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 20272 14278 20300 19926
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 19996 14006 20024 14214
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 20364 13938 20392 21134
rect 20456 18766 20484 21286
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20732 20754 20760 20946
rect 20640 20726 20760 20754
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20456 16590 20484 17070
rect 20548 16590 20576 19382
rect 20640 18902 20668 20726
rect 20824 20058 20852 28970
rect 20916 21418 20944 28970
rect 21008 27674 21036 32694
rect 21088 32428 21140 32434
rect 21088 32370 21140 32376
rect 21100 32337 21128 32370
rect 21086 32328 21142 32337
rect 21086 32263 21142 32272
rect 21100 30122 21128 32263
rect 21192 32026 21220 33050
rect 21284 32774 21312 33254
rect 21560 32978 21588 35498
rect 21652 34746 21680 38286
rect 21640 34740 21692 34746
rect 21640 34682 21692 34688
rect 21640 34604 21692 34610
rect 21640 34546 21692 34552
rect 21456 32972 21508 32978
rect 21456 32914 21508 32920
rect 21548 32972 21600 32978
rect 21548 32914 21600 32920
rect 21468 32881 21496 32914
rect 21454 32872 21510 32881
rect 21454 32807 21510 32816
rect 21272 32768 21324 32774
rect 21272 32710 21324 32716
rect 21272 32564 21324 32570
rect 21272 32506 21324 32512
rect 21180 32020 21232 32026
rect 21180 31962 21232 31968
rect 21192 31754 21220 31962
rect 21284 31754 21312 32506
rect 21560 32366 21588 32914
rect 21652 32434 21680 34546
rect 21744 33998 21772 38762
rect 21928 38418 21956 43590
rect 22020 42770 22048 46854
rect 22112 46714 22140 52958
rect 22192 52896 22244 52902
rect 22192 52838 22244 52844
rect 22100 46708 22152 46714
rect 22100 46650 22152 46656
rect 22100 45076 22152 45082
rect 22100 45018 22152 45024
rect 22112 44470 22140 45018
rect 22100 44464 22152 44470
rect 22100 44406 22152 44412
rect 22008 42764 22060 42770
rect 22008 42706 22060 42712
rect 22008 41472 22060 41478
rect 22008 41414 22060 41420
rect 22020 41274 22048 41414
rect 22008 41268 22060 41274
rect 22008 41210 22060 41216
rect 22008 40656 22060 40662
rect 22008 40598 22060 40604
rect 22020 40118 22048 40598
rect 22112 40186 22140 44406
rect 22204 43858 22232 52838
rect 22284 45280 22336 45286
rect 22284 45222 22336 45228
rect 22296 44878 22324 45222
rect 22284 44872 22336 44878
rect 22284 44814 22336 44820
rect 22296 44334 22324 44814
rect 22284 44328 22336 44334
rect 22284 44270 22336 44276
rect 22296 44198 22324 44270
rect 22284 44192 22336 44198
rect 22284 44134 22336 44140
rect 22192 43852 22244 43858
rect 22192 43794 22244 43800
rect 22192 42696 22244 42702
rect 22296 42650 22324 44134
rect 22388 43450 22416 53654
rect 22468 53440 22520 53446
rect 22468 53382 22520 53388
rect 22480 47122 22508 53382
rect 22572 53242 22600 54046
rect 22744 53984 22796 53990
rect 22742 53952 22744 53961
rect 22796 53952 22798 53961
rect 22742 53887 22798 53896
rect 22848 53582 22876 56200
rect 23216 55214 23244 56200
rect 23386 56128 23442 56137
rect 23386 56063 23442 56072
rect 23216 55186 23336 55214
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 22836 53576 22888 53582
rect 22836 53518 22888 53524
rect 23308 53242 23336 55186
rect 23400 53582 23428 56063
rect 23388 53576 23440 53582
rect 23388 53518 23440 53524
rect 22560 53236 22612 53242
rect 22560 53178 22612 53184
rect 23296 53236 23348 53242
rect 23296 53178 23348 53184
rect 23584 53106 23612 56200
rect 24490 55448 24546 55457
rect 24490 55383 24546 55392
rect 24504 54330 24532 55383
rect 24766 54632 24822 54641
rect 24766 54567 24822 54576
rect 24492 54324 24544 54330
rect 24492 54266 24544 54272
rect 24124 53984 24176 53990
rect 24124 53926 24176 53932
rect 23572 53100 23624 53106
rect 23572 53042 23624 53048
rect 23940 52896 23992 52902
rect 23940 52838 23992 52844
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 23492 52494 23520 52838
rect 23952 52698 23980 54130
rect 24136 54126 24164 56200
rect 24504 55214 24532 56200
rect 24412 55186 24532 55214
rect 24124 54120 24176 54126
rect 24124 54062 24176 54068
rect 24032 53576 24084 53582
rect 24032 53518 24084 53524
rect 23940 52692 23992 52698
rect 23940 52634 23992 52640
rect 23480 52488 23532 52494
rect 23480 52430 23532 52436
rect 23296 52352 23348 52358
rect 23296 52294 23348 52300
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22744 51264 22796 51270
rect 22744 51206 22796 51212
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 23848 47592 23900 47598
rect 23848 47534 23900 47540
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22468 47116 22520 47122
rect 22468 47058 22520 47064
rect 22560 47116 22612 47122
rect 22560 47058 22612 47064
rect 22572 45082 22600 47058
rect 22652 46436 22704 46442
rect 22652 46378 22704 46384
rect 22560 45076 22612 45082
rect 22560 45018 22612 45024
rect 22664 44962 22692 46378
rect 23296 46368 23348 46374
rect 23296 46310 23348 46316
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22744 45416 22796 45422
rect 22744 45358 22796 45364
rect 22480 44934 22692 44962
rect 22376 43444 22428 43450
rect 22376 43386 22428 43392
rect 22244 42644 22324 42650
rect 22192 42638 22324 42644
rect 22204 42622 22324 42638
rect 22192 42560 22244 42566
rect 22192 42502 22244 42508
rect 22204 40730 22232 42502
rect 22296 42158 22324 42622
rect 22284 42152 22336 42158
rect 22284 42094 22336 42100
rect 22480 41970 22508 44934
rect 22560 44804 22612 44810
rect 22560 44746 22612 44752
rect 22572 44538 22600 44746
rect 22756 44742 22784 45358
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 22744 44736 22796 44742
rect 22744 44678 22796 44684
rect 22560 44532 22612 44538
rect 22560 44474 22612 44480
rect 22572 42770 22600 44474
rect 22652 44464 22704 44470
rect 22652 44406 22704 44412
rect 22664 44334 22692 44406
rect 22652 44328 22704 44334
rect 22652 44270 22704 44276
rect 22652 43240 22704 43246
rect 22652 43182 22704 43188
rect 22560 42764 22612 42770
rect 22560 42706 22612 42712
rect 22388 41942 22508 41970
rect 22284 41540 22336 41546
rect 22284 41482 22336 41488
rect 22192 40724 22244 40730
rect 22192 40666 22244 40672
rect 22192 40452 22244 40458
rect 22192 40394 22244 40400
rect 22100 40180 22152 40186
rect 22100 40122 22152 40128
rect 22008 40112 22060 40118
rect 22008 40054 22060 40060
rect 22204 39370 22232 40394
rect 22296 39642 22324 41482
rect 22388 41206 22416 41942
rect 22572 41834 22600 42706
rect 22480 41806 22600 41834
rect 22480 41682 22508 41806
rect 22560 41744 22612 41750
rect 22560 41686 22612 41692
rect 22468 41676 22520 41682
rect 22468 41618 22520 41624
rect 22376 41200 22428 41206
rect 22376 41142 22428 41148
rect 22284 39636 22336 39642
rect 22284 39578 22336 39584
rect 22388 39506 22416 41142
rect 22468 40656 22520 40662
rect 22468 40598 22520 40604
rect 22376 39500 22428 39506
rect 22376 39442 22428 39448
rect 22192 39364 22244 39370
rect 22192 39306 22244 39312
rect 22100 38888 22152 38894
rect 22100 38830 22152 38836
rect 21916 38412 21968 38418
rect 21916 38354 21968 38360
rect 22112 37262 22140 38830
rect 22376 38480 22428 38486
rect 22376 38422 22428 38428
rect 22284 38208 22336 38214
rect 22284 38150 22336 38156
rect 22100 37256 22152 37262
rect 22100 37198 22152 37204
rect 22112 36786 22140 37198
rect 22100 36780 22152 36786
rect 22100 36722 22152 36728
rect 21916 36712 21968 36718
rect 21916 36654 21968 36660
rect 21824 36304 21876 36310
rect 21824 36246 21876 36252
rect 21732 33992 21784 33998
rect 21732 33934 21784 33940
rect 21836 33114 21864 36246
rect 21824 33108 21876 33114
rect 21824 33050 21876 33056
rect 21928 32994 21956 36654
rect 22100 36100 22152 36106
rect 22100 36042 22152 36048
rect 22112 34746 22140 36042
rect 22192 35692 22244 35698
rect 22192 35634 22244 35640
rect 22204 35086 22232 35634
rect 22192 35080 22244 35086
rect 22192 35022 22244 35028
rect 22100 34740 22152 34746
rect 22100 34682 22152 34688
rect 22100 34468 22152 34474
rect 22100 34410 22152 34416
rect 22008 34400 22060 34406
rect 22008 34342 22060 34348
rect 21836 32966 21956 32994
rect 21640 32428 21692 32434
rect 21640 32370 21692 32376
rect 21548 32360 21600 32366
rect 21548 32302 21600 32308
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 21376 31890 21404 32166
rect 21364 31884 21416 31890
rect 21364 31826 21416 31832
rect 21560 31754 21588 32302
rect 21836 31822 21864 32966
rect 21914 32600 21970 32609
rect 21914 32535 21916 32544
rect 21968 32535 21970 32544
rect 21916 32506 21968 32512
rect 21824 31816 21876 31822
rect 21824 31758 21876 31764
rect 21180 31748 21232 31754
rect 21284 31726 21404 31754
rect 21560 31726 21680 31754
rect 21180 31690 21232 31696
rect 21088 30116 21140 30122
rect 21088 30058 21140 30064
rect 21180 29708 21232 29714
rect 21180 29650 21232 29656
rect 21192 28694 21220 29650
rect 21272 28756 21324 28762
rect 21272 28698 21324 28704
rect 21180 28688 21232 28694
rect 21180 28630 21232 28636
rect 20996 27668 21048 27674
rect 20996 27610 21048 27616
rect 21088 27600 21140 27606
rect 21088 27542 21140 27548
rect 20996 26240 21048 26246
rect 20996 26182 21048 26188
rect 21008 25702 21036 26182
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21008 24206 21036 25638
rect 21100 25362 21128 27542
rect 21192 26926 21220 28630
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 21192 26314 21220 26862
rect 21180 26308 21232 26314
rect 21180 26250 21232 26256
rect 21180 25696 21232 25702
rect 21180 25638 21232 25644
rect 21088 25356 21140 25362
rect 21088 25298 21140 25304
rect 20996 24200 21048 24206
rect 20996 24142 21048 24148
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20904 21412 20956 21418
rect 20904 21354 20956 21360
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20824 19514 20852 19994
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20628 18896 20680 18902
rect 20628 18838 20680 18844
rect 20640 18358 20668 18838
rect 20628 18352 20680 18358
rect 20628 18294 20680 18300
rect 20640 17610 20668 18294
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20640 17202 20668 17546
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 19628 12406 19748 12434
rect 19524 11892 19576 11898
rect 19628 11880 19656 12406
rect 19628 11852 19748 11880
rect 19524 11834 19576 11840
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19628 10810 19656 10950
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 18880 8560 18932 8566
rect 18880 8502 18932 8508
rect 18708 6886 18828 6914
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18708 4146 18736 6886
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17684 2508 17736 2514
rect 17684 2450 17736 2456
rect 17880 800 17908 3538
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18340 1170 18368 2314
rect 18248 1142 18368 1170
rect 18248 800 18276 1142
rect 18616 800 18644 3062
rect 18984 800 19012 3402
rect 19352 800 19380 5102
rect 19444 2446 19472 9998
rect 19720 6914 19748 11852
rect 19812 10062 19840 13126
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19904 11762 19932 12038
rect 19996 11898 20024 12242
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19996 10606 20024 11834
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 19536 6886 19748 6914
rect 19536 5234 19564 6886
rect 19616 5296 19668 5302
rect 19616 5238 19668 5244
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19628 3942 19656 5238
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19708 4616 19760 4622
rect 19708 4558 19760 4564
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19720 800 19748 4558
rect 19904 3126 19932 4626
rect 20076 4072 20128 4078
rect 20180 4049 20208 13806
rect 20364 13530 20392 13874
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20456 11694 20484 14758
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20456 7886 20484 11630
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20548 5710 20576 13806
rect 20640 11082 20668 15302
rect 20732 14006 20760 19110
rect 21100 17270 21128 21626
rect 21192 19514 21220 25638
rect 21284 22094 21312 28698
rect 21376 27946 21404 31726
rect 21456 31476 21508 31482
rect 21456 31418 21508 31424
rect 21468 29578 21496 31418
rect 21652 31414 21680 31726
rect 21836 31482 21864 31758
rect 21824 31476 21876 31482
rect 21824 31418 21876 31424
rect 21640 31408 21692 31414
rect 21640 31350 21692 31356
rect 21824 30048 21876 30054
rect 21824 29990 21876 29996
rect 21732 29844 21784 29850
rect 21732 29786 21784 29792
rect 21744 29578 21772 29786
rect 21456 29572 21508 29578
rect 21456 29514 21508 29520
rect 21732 29572 21784 29578
rect 21732 29514 21784 29520
rect 21548 29504 21600 29510
rect 21548 29446 21600 29452
rect 21454 29200 21510 29209
rect 21454 29135 21456 29144
rect 21508 29135 21510 29144
rect 21456 29106 21508 29112
rect 21456 28756 21508 28762
rect 21456 28698 21508 28704
rect 21468 28490 21496 28698
rect 21456 28484 21508 28490
rect 21456 28426 21508 28432
rect 21364 27940 21416 27946
rect 21364 27882 21416 27888
rect 21560 24206 21588 29446
rect 21732 27056 21784 27062
rect 21732 26998 21784 27004
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21652 25294 21680 25774
rect 21640 25288 21692 25294
rect 21640 25230 21692 25236
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 21468 23526 21496 24142
rect 21456 23520 21508 23526
rect 21456 23462 21508 23468
rect 21468 22982 21496 23462
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21468 22166 21496 22918
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21456 22160 21508 22166
rect 21456 22102 21508 22108
rect 21284 22066 21404 22094
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21284 17882 21312 19246
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 21088 17264 21140 17270
rect 21088 17206 21140 17212
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 20824 15366 20852 15642
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20812 14884 20864 14890
rect 20812 14826 20864 14832
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 20824 12434 20852 14826
rect 21008 14056 21036 15642
rect 21192 15570 21220 16390
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21192 14482 21220 15506
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 20732 12406 20852 12434
rect 20916 14028 21036 14056
rect 20732 11830 20760 12406
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20640 7886 20668 11018
rect 20824 10538 20852 11018
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 20916 8566 20944 14028
rect 21100 13410 21128 14282
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21192 13938 21220 14010
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 21008 13382 21128 13410
rect 20904 8560 20956 8566
rect 20904 8502 20956 8508
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20640 5710 20668 7210
rect 20824 6798 20852 7686
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20916 5914 20944 7346
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20628 4548 20680 4554
rect 20628 4490 20680 4496
rect 20076 4014 20128 4020
rect 20166 4040 20222 4049
rect 19892 3120 19944 3126
rect 19892 3062 19944 3068
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19904 2514 19932 2790
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 20088 800 20116 4014
rect 20166 3975 20222 3984
rect 20640 2922 20668 4490
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20732 2802 20760 5714
rect 21008 3534 21036 13382
rect 21284 12306 21312 15370
rect 21376 13870 21404 22066
rect 21468 21962 21496 22102
rect 21456 21956 21508 21962
rect 21456 21898 21508 21904
rect 21468 21078 21496 21898
rect 21548 21140 21600 21146
rect 21548 21082 21600 21088
rect 21456 21072 21508 21078
rect 21456 21014 21508 21020
rect 21468 20942 21496 21014
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21560 20754 21588 21082
rect 21652 20806 21680 22510
rect 21744 21894 21772 26998
rect 21836 24138 21864 29990
rect 22020 29646 22048 34342
rect 22112 31278 22140 34410
rect 22204 33522 22232 35022
rect 22296 34066 22324 38150
rect 22388 37874 22416 38422
rect 22376 37868 22428 37874
rect 22376 37810 22428 37816
rect 22388 35494 22416 37810
rect 22480 37233 22508 40598
rect 22572 40526 22600 41686
rect 22560 40520 22612 40526
rect 22560 40462 22612 40468
rect 22560 39976 22612 39982
rect 22560 39918 22612 39924
rect 22572 39506 22600 39918
rect 22560 39500 22612 39506
rect 22560 39442 22612 39448
rect 22560 38412 22612 38418
rect 22560 38354 22612 38360
rect 22466 37224 22522 37233
rect 22466 37159 22522 37168
rect 22376 35488 22428 35494
rect 22376 35430 22428 35436
rect 22376 35284 22428 35290
rect 22376 35226 22428 35232
rect 22284 34060 22336 34066
rect 22284 34002 22336 34008
rect 22192 33516 22244 33522
rect 22192 33458 22244 33464
rect 22204 31278 22232 33458
rect 22388 32910 22416 35226
rect 22572 35018 22600 38354
rect 22664 37738 22692 43182
rect 22756 40662 22784 44678
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22836 42152 22888 42158
rect 22836 42094 22888 42100
rect 22848 41070 22876 42094
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 23204 41812 23256 41818
rect 23204 41754 23256 41760
rect 22836 41064 22888 41070
rect 22836 41006 22888 41012
rect 22744 40656 22796 40662
rect 22744 40598 22796 40604
rect 22848 40118 22876 41006
rect 23216 40984 23244 41754
rect 23308 41682 23336 46310
rect 23480 45960 23532 45966
rect 23480 45902 23532 45908
rect 23492 45665 23520 45902
rect 23478 45656 23534 45665
rect 23478 45591 23534 45600
rect 23388 43852 23440 43858
rect 23388 43794 23440 43800
rect 23400 42362 23428 43794
rect 23572 43376 23624 43382
rect 23572 43318 23624 43324
rect 23480 43240 23532 43246
rect 23480 43182 23532 43188
rect 23388 42356 23440 42362
rect 23388 42298 23440 42304
rect 23296 41676 23348 41682
rect 23296 41618 23348 41624
rect 23216 40956 23336 40984
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 23112 40656 23164 40662
rect 23110 40624 23112 40633
rect 23164 40624 23166 40633
rect 23308 40610 23336 40956
rect 23110 40559 23166 40568
rect 23216 40582 23336 40610
rect 22928 40520 22980 40526
rect 22926 40488 22928 40497
rect 22980 40488 22982 40497
rect 22926 40423 22982 40432
rect 22836 40112 22888 40118
rect 22836 40054 22888 40060
rect 23216 39930 23244 40582
rect 23296 40520 23348 40526
rect 23296 40462 23348 40468
rect 23308 40390 23336 40462
rect 23296 40384 23348 40390
rect 23296 40326 23348 40332
rect 22848 39902 23244 39930
rect 22848 38486 22876 39902
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22836 38480 22888 38486
rect 22836 38422 22888 38428
rect 22744 37868 22796 37874
rect 22744 37810 22796 37816
rect 22652 37732 22704 37738
rect 22652 37674 22704 37680
rect 22664 36854 22692 37674
rect 22652 36848 22704 36854
rect 22652 36790 22704 36796
rect 22756 35894 22784 37810
rect 22848 37806 22876 38422
rect 23308 37874 23336 40326
rect 23400 38894 23428 42298
rect 23492 42158 23520 43182
rect 23480 42152 23532 42158
rect 23480 42094 23532 42100
rect 23584 41970 23612 43318
rect 23664 42696 23716 42702
rect 23664 42638 23716 42644
rect 23756 42696 23808 42702
rect 23756 42638 23808 42644
rect 23492 41942 23612 41970
rect 23492 41682 23520 41942
rect 23480 41676 23532 41682
rect 23480 41618 23532 41624
rect 23572 41676 23624 41682
rect 23572 41618 23624 41624
rect 23492 41274 23520 41618
rect 23480 41268 23532 41274
rect 23480 41210 23532 41216
rect 23492 39506 23520 41210
rect 23584 40458 23612 41618
rect 23676 41070 23704 42638
rect 23768 42294 23796 42638
rect 23756 42288 23808 42294
rect 23756 42230 23808 42236
rect 23664 41064 23716 41070
rect 23664 41006 23716 41012
rect 23860 40662 23888 47534
rect 23952 46714 23980 52838
rect 23940 46708 23992 46714
rect 23940 46650 23992 46656
rect 24032 45484 24084 45490
rect 24032 45426 24084 45432
rect 24044 45286 24072 45426
rect 24032 45280 24084 45286
rect 24032 45222 24084 45228
rect 24044 44878 24072 45222
rect 24032 44872 24084 44878
rect 24032 44814 24084 44820
rect 23940 44328 23992 44334
rect 23940 44270 23992 44276
rect 23848 40656 23900 40662
rect 23848 40598 23900 40604
rect 23572 40452 23624 40458
rect 23572 40394 23624 40400
rect 23756 39840 23808 39846
rect 23756 39782 23808 39788
rect 23480 39500 23532 39506
rect 23480 39442 23532 39448
rect 23572 39432 23624 39438
rect 23572 39374 23624 39380
rect 23388 38888 23440 38894
rect 23388 38830 23440 38836
rect 23400 38486 23428 38830
rect 23584 38826 23612 39374
rect 23768 39030 23796 39782
rect 23756 39024 23808 39030
rect 23756 38966 23808 38972
rect 23572 38820 23624 38826
rect 23572 38762 23624 38768
rect 23388 38480 23440 38486
rect 23388 38422 23440 38428
rect 23480 38276 23532 38282
rect 23480 38218 23532 38224
rect 23492 37942 23520 38218
rect 23584 38214 23612 38762
rect 23664 38752 23716 38758
rect 23664 38694 23716 38700
rect 23676 38418 23704 38694
rect 23664 38412 23716 38418
rect 23664 38354 23716 38360
rect 23768 38298 23796 38966
rect 23848 38412 23900 38418
rect 23848 38354 23900 38360
rect 23676 38270 23796 38298
rect 23676 38214 23704 38270
rect 23572 38208 23624 38214
rect 23572 38150 23624 38156
rect 23664 38208 23716 38214
rect 23664 38150 23716 38156
rect 23756 38208 23808 38214
rect 23756 38150 23808 38156
rect 23480 37936 23532 37942
rect 23480 37878 23532 37884
rect 23296 37868 23348 37874
rect 23296 37810 23348 37816
rect 22836 37800 22888 37806
rect 22836 37742 22888 37748
rect 22836 37664 22888 37670
rect 22836 37606 22888 37612
rect 22848 36786 22876 37606
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 23584 37466 23612 38150
rect 23572 37460 23624 37466
rect 23572 37402 23624 37408
rect 23388 36848 23440 36854
rect 23388 36790 23440 36796
rect 22836 36780 22888 36786
rect 22836 36722 22888 36728
rect 22664 35866 22784 35894
rect 22560 35012 22612 35018
rect 22560 34954 22612 34960
rect 22466 34912 22522 34921
rect 22466 34847 22522 34856
rect 22480 34746 22508 34847
rect 22468 34740 22520 34746
rect 22468 34682 22520 34688
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22376 32904 22428 32910
rect 22376 32846 22428 32852
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 22192 31272 22244 31278
rect 22192 31214 22244 31220
rect 22204 30258 22232 31214
rect 22284 31136 22336 31142
rect 22284 31078 22336 31084
rect 22296 30734 22324 31078
rect 22480 30734 22508 33798
rect 22572 33046 22600 34954
rect 22560 33040 22612 33046
rect 22560 32982 22612 32988
rect 22664 32337 22692 35866
rect 22848 35698 22876 36722
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 23296 36032 23348 36038
rect 23296 35974 23348 35980
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22744 35624 22796 35630
rect 22744 35566 22796 35572
rect 22756 34746 22784 35566
rect 22836 35488 22888 35494
rect 22836 35430 22888 35436
rect 22744 34740 22796 34746
rect 22744 34682 22796 34688
rect 22744 32904 22796 32910
rect 22742 32872 22744 32881
rect 22848 32892 22876 35430
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23020 35148 23072 35154
rect 23020 35090 23072 35096
rect 23032 35018 23060 35090
rect 23020 35012 23072 35018
rect 23020 34954 23072 34960
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 22796 32872 22876 32892
rect 22798 32864 22876 32872
rect 22742 32807 22798 32816
rect 22650 32328 22706 32337
rect 22650 32263 22706 32272
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22468 30728 22520 30734
rect 22468 30670 22520 30676
rect 22284 30592 22336 30598
rect 22284 30534 22336 30540
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 22008 28620 22060 28626
rect 22008 28562 22060 28568
rect 22020 28082 22048 28562
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 22020 27554 22048 28018
rect 22100 27872 22152 27878
rect 22100 27814 22152 27820
rect 21928 27538 22048 27554
rect 21916 27532 22048 27538
rect 21968 27526 22048 27532
rect 21916 27474 21968 27480
rect 22020 26926 22048 27526
rect 22008 26920 22060 26926
rect 22008 26862 22060 26868
rect 22020 26518 22048 26862
rect 22008 26512 22060 26518
rect 22008 26454 22060 26460
rect 22020 24818 22048 26454
rect 22112 24970 22140 27814
rect 22192 27396 22244 27402
rect 22192 27338 22244 27344
rect 22204 26586 22232 27338
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 22204 25906 22232 26522
rect 22296 26382 22324 30534
rect 22560 29708 22612 29714
rect 22560 29650 22612 29656
rect 22374 29336 22430 29345
rect 22374 29271 22430 29280
rect 22284 26376 22336 26382
rect 22284 26318 22336 26324
rect 22388 26042 22416 29271
rect 22468 29232 22520 29238
rect 22468 29174 22520 29180
rect 22480 26450 22508 29174
rect 22572 26602 22600 29650
rect 22572 26586 22692 26602
rect 22572 26580 22704 26586
rect 22572 26574 22652 26580
rect 22652 26522 22704 26528
rect 22560 26512 22612 26518
rect 22560 26454 22612 26460
rect 22468 26444 22520 26450
rect 22468 26386 22520 26392
rect 22376 26036 22428 26042
rect 22376 25978 22428 25984
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22388 25378 22416 25978
rect 22388 25350 22508 25378
rect 22376 25220 22428 25226
rect 22376 25162 22428 25168
rect 22112 24942 22324 24970
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 22112 24274 22140 24754
rect 22100 24268 22152 24274
rect 22100 24210 22152 24216
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 22112 23730 22140 24210
rect 22192 24132 22244 24138
rect 22192 24074 22244 24080
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22020 22642 22048 23666
rect 22204 23066 22232 24074
rect 22112 23038 22232 23066
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 22020 22098 22048 22578
rect 22008 22092 22060 22098
rect 22008 22034 22060 22040
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 22020 21622 22048 22034
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21468 20726 21588 20754
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21468 14074 21496 20726
rect 21652 20398 21680 20742
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21560 16046 21588 19654
rect 21824 19508 21876 19514
rect 21824 19450 21876 19456
rect 21836 19310 21864 19450
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 21732 18692 21784 18698
rect 21732 18634 21784 18640
rect 21744 17746 21772 18634
rect 21732 17740 21784 17746
rect 21732 17682 21784 17688
rect 21744 16590 21772 17682
rect 21836 16794 21864 19246
rect 22020 18698 22048 19246
rect 22008 18692 22060 18698
rect 22008 18634 22060 18640
rect 22112 18290 22140 23038
rect 22296 22094 22324 24942
rect 22204 22066 22324 22094
rect 22204 20942 22232 22066
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 22112 16674 22140 18022
rect 22020 16646 22140 16674
rect 21732 16584 21784 16590
rect 22020 16574 22048 16646
rect 22020 16546 22140 16574
rect 21732 16526 21784 16532
rect 22112 16182 22140 16546
rect 22100 16176 22152 16182
rect 22100 16118 22152 16124
rect 21548 16040 21600 16046
rect 21548 15982 21600 15988
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 21376 12918 21404 13126
rect 21364 12912 21416 12918
rect 21364 12854 21416 12860
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 21100 9586 21128 12038
rect 21376 11558 21404 12854
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21560 10606 21588 15302
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21732 14000 21784 14006
rect 21732 13942 21784 13948
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21744 10554 21772 13942
rect 21836 12782 21864 14214
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21836 12306 21864 12718
rect 21928 12306 21956 15846
rect 22112 15706 22140 15846
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22204 14006 22232 18090
rect 22296 15502 22324 21286
rect 22388 20466 22416 25162
rect 22480 25158 22508 25350
rect 22468 25152 22520 25158
rect 22468 25094 22520 25100
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22480 16182 22508 24006
rect 22572 21486 22600 26454
rect 22664 25362 22692 26522
rect 22756 26042 22784 32807
rect 23204 32360 23256 32366
rect 23202 32328 23204 32337
rect 23256 32328 23258 32337
rect 23202 32263 23258 32272
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23308 31482 23336 35974
rect 23400 35894 23428 36790
rect 23664 36372 23716 36378
rect 23664 36314 23716 36320
rect 23676 36122 23704 36314
rect 23768 36242 23796 38150
rect 23860 37942 23888 38354
rect 23952 38350 23980 44270
rect 24032 40520 24084 40526
rect 24032 40462 24084 40468
rect 24044 40390 24072 40462
rect 24032 40384 24084 40390
rect 24032 40326 24084 40332
rect 24044 40118 24072 40326
rect 24032 40112 24084 40118
rect 24032 40054 24084 40060
rect 24044 38962 24072 40054
rect 24032 38956 24084 38962
rect 24032 38898 24084 38904
rect 23940 38344 23992 38350
rect 23940 38286 23992 38292
rect 23848 37936 23900 37942
rect 23848 37878 23900 37884
rect 23860 36922 23888 37878
rect 24044 37398 24072 38898
rect 24032 37392 24084 37398
rect 24032 37334 24084 37340
rect 24030 37224 24086 37233
rect 24030 37159 24086 37168
rect 23848 36916 23900 36922
rect 23848 36858 23900 36864
rect 23756 36236 23808 36242
rect 23756 36178 23808 36184
rect 23676 36094 23796 36122
rect 23768 36038 23796 36094
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23756 36032 23808 36038
rect 23756 35974 23808 35980
rect 23676 35894 23704 35974
rect 23400 35866 23520 35894
rect 23388 35624 23440 35630
rect 23388 35566 23440 35572
rect 23400 34950 23428 35566
rect 23492 35494 23520 35866
rect 23584 35866 23704 35894
rect 23480 35488 23532 35494
rect 23480 35430 23532 35436
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 23400 34066 23428 34886
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23492 33386 23520 35430
rect 23584 34542 23612 35866
rect 23572 34536 23624 34542
rect 23572 34478 23624 34484
rect 23664 34536 23716 34542
rect 23664 34478 23716 34484
rect 23676 33590 23704 34478
rect 23664 33584 23716 33590
rect 23664 33526 23716 33532
rect 23768 33538 23796 35974
rect 23860 34474 23888 36858
rect 23940 35760 23992 35766
rect 23940 35702 23992 35708
rect 23952 35630 23980 35702
rect 23940 35624 23992 35630
rect 23940 35566 23992 35572
rect 23952 35154 23980 35566
rect 23940 35148 23992 35154
rect 23940 35090 23992 35096
rect 24044 34610 24072 37159
rect 24032 34604 24084 34610
rect 24032 34546 24084 34552
rect 23848 34468 23900 34474
rect 23848 34410 23900 34416
rect 23768 33510 23888 33538
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 23480 33380 23532 33386
rect 23480 33322 23532 33328
rect 23388 31952 23440 31958
rect 23388 31894 23440 31900
rect 23296 31476 23348 31482
rect 23296 31418 23348 31424
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 22744 29708 22796 29714
rect 22744 29650 22796 29656
rect 22744 29504 22796 29510
rect 22744 29446 22796 29452
rect 22652 28212 22704 28218
rect 22652 28154 22704 28160
rect 22468 25968 22520 25974
rect 22468 25910 22520 25916
rect 22652 25968 22704 25974
rect 22652 25910 22704 25916
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22560 25832 22612 25838
rect 22560 25774 22612 25780
rect 22284 25764 22336 25770
rect 22284 25706 22336 25712
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 22020 25242 22048 25298
rect 22020 25214 22232 25242
rect 21732 25152 21784 25158
rect 21732 25094 21784 25100
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 21916 23112 21968 23118
rect 21916 23054 21968 23060
rect 21640 22704 21692 22710
rect 21640 22646 21692 22652
rect 21928 22574 21956 23054
rect 21916 22568 21968 22574
rect 21916 22510 21968 22516
rect 21640 22500 21692 22506
rect 21640 22442 21692 22448
rect 21652 21622 21680 22442
rect 22112 22166 22140 24686
rect 22204 24682 22232 25214
rect 22192 24676 22244 24682
rect 22192 24618 22244 24624
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22112 21010 22140 21490
rect 22204 21078 22232 22714
rect 22192 21072 22244 21078
rect 22192 21014 22244 21020
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21836 20602 21864 20878
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21732 19712 21784 19718
rect 21732 19654 21784 19660
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20732 17270 20760 17546
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20732 17134 20760 17206
rect 21192 17134 21220 17478
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21192 16658 21220 17070
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21364 16448 21416 16454
rect 21364 16390 21416 16396
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 19996 12406 20116 12434
rect 19996 12374 20024 12406
rect 19984 12368 20036 12374
rect 19984 12310 20036 12316
rect 20364 11626 20392 14758
rect 21008 14074 21036 15302
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 20916 13190 20944 13738
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20916 12918 20944 13126
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19720 5234 19748 6666
rect 19996 5710 20024 11562
rect 21100 10674 21128 13466
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20260 7812 20312 7818
rect 20260 7754 20312 7760
rect 20168 6316 20220 6322
rect 20168 6258 20220 6264
rect 20180 5914 20208 6258
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20272 5846 20300 7754
rect 20260 5840 20312 5846
rect 20260 5782 20312 5788
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19800 5296 19852 5302
rect 19800 5238 19852 5244
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19708 5228 19760 5234
rect 19708 5170 19760 5176
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 18972 2576 19024 2582
rect 18972 2518 19024 2524
rect 19168 800 19196 3402
rect 19536 800 19564 5102
rect 19812 3670 19840 5238
rect 20536 5092 20588 5098
rect 20536 5034 20588 5040
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19800 3664 19852 3670
rect 19800 3606 19852 3612
rect 19904 2854 19932 4626
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19996 2258 20024 2858
rect 19904 2230 20024 2258
rect 19904 800 19932 2230
rect 20272 800 20300 4014
rect 20548 2990 20576 5034
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20640 800 20668 5714
rect 20732 5710 20760 8842
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 21008 3942 21036 7278
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 21100 3534 21128 7754
rect 21192 4622 21220 13398
rect 21284 7886 21312 14758
rect 21376 13870 21404 16390
rect 21468 14414 21496 18566
rect 21548 17128 21600 17134
rect 21548 17070 21600 17076
rect 21560 16794 21588 17070
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 13190 21404 13670
rect 21560 13394 21588 16730
rect 21640 16448 21692 16454
rect 21640 16390 21692 16396
rect 21652 15609 21680 16390
rect 21638 15600 21694 15609
rect 21638 15535 21694 15544
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 21376 12986 21404 13126
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21376 12102 21404 12922
rect 21456 12776 21508 12782
rect 21560 12764 21588 13330
rect 21652 13190 21680 15535
rect 21744 14346 21772 19654
rect 22100 19440 22152 19446
rect 22100 19382 22152 19388
rect 22112 19281 22140 19382
rect 22296 19378 22324 25706
rect 22376 23316 22428 23322
rect 22376 23258 22428 23264
rect 22388 22642 22416 23258
rect 22376 22636 22428 22642
rect 22376 22578 22428 22584
rect 22388 22234 22416 22578
rect 22376 22228 22428 22234
rect 22376 22170 22428 22176
rect 22376 21956 22428 21962
rect 22376 21898 22428 21904
rect 22388 20602 22416 21898
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22098 19272 22154 19281
rect 22098 19207 22154 19216
rect 22572 18970 22600 25774
rect 22664 25226 22692 25910
rect 22652 25220 22704 25226
rect 22652 25162 22704 25168
rect 22756 24954 22784 29446
rect 22848 27402 22876 30126
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 23400 29714 23428 31894
rect 23480 31884 23532 31890
rect 23480 31826 23532 31832
rect 23492 31226 23520 31826
rect 23492 31198 23612 31226
rect 23584 31142 23612 31198
rect 23572 31136 23624 31142
rect 23572 31078 23624 31084
rect 23480 30932 23532 30938
rect 23480 30874 23532 30880
rect 23492 30598 23520 30874
rect 23480 30592 23532 30598
rect 23480 30534 23532 30540
rect 23584 30326 23612 31078
rect 23572 30320 23624 30326
rect 23572 30262 23624 30268
rect 23388 29708 23440 29714
rect 23388 29650 23440 29656
rect 22836 29504 22888 29510
rect 22836 29446 22888 29452
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 22848 28626 22876 29446
rect 23308 29034 23336 29446
rect 23584 29102 23612 30262
rect 23768 30190 23796 33390
rect 23860 30938 23888 33510
rect 23940 33108 23992 33114
rect 23940 33050 23992 33056
rect 23848 30932 23900 30938
rect 23848 30874 23900 30880
rect 23756 30184 23808 30190
rect 23756 30126 23808 30132
rect 23768 29714 23796 30126
rect 23756 29708 23808 29714
rect 23756 29650 23808 29656
rect 23848 29572 23900 29578
rect 23848 29514 23900 29520
rect 23860 29306 23888 29514
rect 23848 29300 23900 29306
rect 23848 29242 23900 29248
rect 23572 29096 23624 29102
rect 23572 29038 23624 29044
rect 23296 29028 23348 29034
rect 23296 28970 23348 28976
rect 23480 29028 23532 29034
rect 23480 28970 23532 28976
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 22836 28620 22888 28626
rect 22836 28562 22888 28568
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 23388 27532 23440 27538
rect 23388 27474 23440 27480
rect 23112 27328 23164 27334
rect 23112 27270 23164 27276
rect 23124 27062 23152 27270
rect 23400 27062 23428 27474
rect 23112 27056 23164 27062
rect 23112 26998 23164 27004
rect 23388 27056 23440 27062
rect 23388 26998 23440 27004
rect 23124 26926 23152 26998
rect 23112 26920 23164 26926
rect 23112 26862 23164 26868
rect 23204 26920 23256 26926
rect 23256 26880 23336 26908
rect 23204 26862 23256 26868
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 22744 26036 22796 26042
rect 22744 25978 22796 25984
rect 22756 25922 22784 25978
rect 22756 25894 22876 25922
rect 22744 25832 22796 25838
rect 22744 25774 22796 25780
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 22664 24886 22692 25298
rect 22652 24880 22704 24886
rect 22652 24822 22704 24828
rect 22652 24676 22704 24682
rect 22652 24618 22704 24624
rect 22664 23050 22692 24618
rect 22652 23044 22704 23050
rect 22652 22986 22704 22992
rect 22652 22092 22704 22098
rect 22652 22034 22704 22040
rect 22664 21486 22692 22034
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22560 21072 22612 21078
rect 22560 21014 22612 21020
rect 22572 19446 22600 21014
rect 22560 19440 22612 19446
rect 22560 19382 22612 19388
rect 22572 18850 22600 19382
rect 22756 19310 22784 25774
rect 22848 25498 22876 25894
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 22836 25492 22888 25498
rect 22836 25434 22888 25440
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23308 23118 23336 26880
rect 23400 26518 23428 26998
rect 23388 26512 23440 26518
rect 23388 26454 23440 26460
rect 23400 26314 23428 26454
rect 23388 26308 23440 26314
rect 23388 26250 23440 26256
rect 23492 24206 23520 28970
rect 23848 26784 23900 26790
rect 23848 26726 23900 26732
rect 23860 25906 23888 26726
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 23756 25764 23808 25770
rect 23756 25706 23808 25712
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23480 23792 23532 23798
rect 23532 23740 23612 23746
rect 23480 23734 23612 23740
rect 23492 23718 23612 23734
rect 23584 23662 23612 23718
rect 23572 23656 23624 23662
rect 23572 23598 23624 23604
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23294 22808 23350 22817
rect 23294 22743 23350 22752
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 22848 21554 22876 22034
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23308 20398 23336 22743
rect 23492 21690 23520 22918
rect 23584 22778 23612 23598
rect 23664 23248 23716 23254
rect 23664 23190 23716 23196
rect 23572 22772 23624 22778
rect 23572 22714 23624 22720
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 23584 22030 23612 22578
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23584 21690 23612 21966
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 23676 21622 23704 23190
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23386 21176 23442 21185
rect 23386 21111 23442 21120
rect 23400 20534 23428 21111
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22652 19168 22704 19174
rect 22652 19110 22704 19116
rect 22664 18850 22692 19110
rect 22756 18970 22784 19246
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22744 18964 22796 18970
rect 22744 18906 22796 18912
rect 22572 18822 22692 18850
rect 22664 18698 22692 18822
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 22652 18692 22704 18698
rect 22652 18634 22704 18640
rect 22572 17882 22600 18634
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22664 17610 22692 18634
rect 22756 18086 22784 18906
rect 23388 18216 23440 18222
rect 23388 18158 23440 18164
rect 22744 18080 22796 18086
rect 22744 18022 22796 18028
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23400 17921 23428 18158
rect 23386 17912 23442 17921
rect 22744 17876 22796 17882
rect 23386 17847 23442 17856
rect 22744 17818 22796 17824
rect 22652 17604 22704 17610
rect 22652 17546 22704 17552
rect 22652 17060 22704 17066
rect 22652 17002 22704 17008
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22388 15162 22416 16050
rect 22560 15972 22612 15978
rect 22560 15914 22612 15920
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 22008 13728 22060 13734
rect 22008 13670 22060 13676
rect 22020 13190 22048 13670
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 22020 12238 22048 12718
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 22572 11762 22600 15914
rect 22664 13326 22692 17002
rect 22756 16046 22784 17818
rect 22836 17604 22888 17610
rect 22836 17546 22888 17552
rect 22848 16674 22876 17546
rect 23768 17202 23796 25706
rect 23952 25294 23980 33050
rect 24136 32774 24164 53926
rect 24780 53582 24808 54567
rect 24952 54188 25004 54194
rect 24952 54130 25004 54136
rect 24964 53825 24992 54130
rect 25136 54052 25188 54058
rect 25136 53994 25188 54000
rect 24950 53816 25006 53825
rect 24950 53751 25006 53760
rect 24768 53576 24820 53582
rect 24768 53518 24820 53524
rect 24216 53508 24268 53514
rect 24216 53450 24268 53456
rect 24228 40474 24256 53450
rect 24780 52698 24808 53518
rect 24768 52692 24820 52698
rect 24768 52634 24820 52640
rect 24768 52488 24820 52494
rect 24768 52430 24820 52436
rect 24780 52193 24808 52430
rect 24766 52184 24822 52193
rect 24964 52154 24992 53751
rect 25044 53100 25096 53106
rect 25044 53042 25096 53048
rect 25056 53009 25084 53042
rect 25042 53000 25098 53009
rect 25042 52935 25098 52944
rect 24766 52119 24822 52128
rect 24952 52148 25004 52154
rect 24952 52090 25004 52096
rect 25044 50924 25096 50930
rect 25044 50866 25096 50872
rect 25056 50561 25084 50866
rect 25042 50552 25098 50561
rect 25042 50487 25098 50496
rect 25148 49722 25176 53994
rect 25872 53440 25924 53446
rect 25872 53382 25924 53388
rect 25228 52896 25280 52902
rect 25228 52838 25280 52844
rect 25056 49694 25176 49722
rect 24860 48000 24912 48006
rect 24860 47942 24912 47948
rect 24768 46980 24820 46986
rect 24768 46922 24820 46928
rect 24492 46504 24544 46510
rect 24492 46446 24544 46452
rect 24676 46504 24728 46510
rect 24780 46481 24808 46922
rect 24676 46446 24728 46452
rect 24766 46472 24822 46481
rect 24504 46170 24532 46446
rect 24492 46164 24544 46170
rect 24492 46106 24544 46112
rect 24400 45484 24452 45490
rect 24400 45426 24452 45432
rect 24228 40446 24348 40474
rect 24216 40384 24268 40390
rect 24216 40326 24268 40332
rect 24228 38962 24256 40326
rect 24216 38956 24268 38962
rect 24216 38898 24268 38904
rect 24320 38282 24348 40446
rect 24308 38276 24360 38282
rect 24308 38218 24360 38224
rect 24308 37936 24360 37942
rect 24228 37884 24308 37890
rect 24228 37878 24360 37884
rect 24228 37862 24348 37878
rect 24228 37398 24256 37862
rect 24216 37392 24268 37398
rect 24216 37334 24268 37340
rect 24228 36786 24256 37334
rect 24216 36780 24268 36786
rect 24216 36722 24268 36728
rect 24228 35154 24256 36722
rect 24412 36038 24440 45426
rect 24492 45416 24544 45422
rect 24492 45358 24544 45364
rect 24504 44742 24532 45358
rect 24584 44872 24636 44878
rect 24584 44814 24636 44820
rect 24492 44736 24544 44742
rect 24492 44678 24544 44684
rect 24596 44470 24624 44814
rect 24584 44464 24636 44470
rect 24584 44406 24636 44412
rect 24596 43654 24624 44406
rect 24584 43648 24636 43654
rect 24584 43590 24636 43596
rect 24596 43382 24624 43590
rect 24584 43376 24636 43382
rect 24584 43318 24636 43324
rect 24596 42634 24624 43318
rect 24584 42628 24636 42634
rect 24584 42570 24636 42576
rect 24596 42514 24624 42570
rect 24504 42486 24624 42514
rect 24504 42294 24532 42486
rect 24492 42288 24544 42294
rect 24492 42230 24544 42236
rect 24504 41460 24532 42230
rect 24584 41472 24636 41478
rect 24504 41432 24584 41460
rect 24504 41206 24532 41432
rect 24584 41414 24636 41420
rect 24492 41200 24544 41206
rect 24492 41142 24544 41148
rect 24504 40526 24532 41142
rect 24492 40520 24544 40526
rect 24492 40462 24544 40468
rect 24584 40384 24636 40390
rect 24582 40352 24584 40361
rect 24636 40352 24638 40361
rect 24582 40287 24638 40296
rect 24492 39976 24544 39982
rect 24492 39918 24544 39924
rect 24504 37806 24532 39918
rect 24584 39296 24636 39302
rect 24584 39238 24636 39244
rect 24492 37800 24544 37806
rect 24492 37742 24544 37748
rect 24504 36242 24532 37742
rect 24492 36236 24544 36242
rect 24492 36178 24544 36184
rect 24400 36032 24452 36038
rect 24400 35974 24452 35980
rect 24400 35828 24452 35834
rect 24400 35770 24452 35776
rect 24216 35148 24268 35154
rect 24216 35090 24268 35096
rect 24216 33448 24268 33454
rect 24216 33390 24268 33396
rect 24124 32768 24176 32774
rect 24124 32710 24176 32716
rect 24032 32496 24084 32502
rect 24032 32438 24084 32444
rect 24044 25362 24072 32438
rect 24228 32026 24256 33390
rect 24216 32020 24268 32026
rect 24216 31962 24268 31968
rect 24228 31414 24256 31962
rect 24412 31482 24440 35770
rect 24596 33998 24624 39238
rect 24688 38298 24716 46446
rect 24766 46407 24822 46416
rect 24768 46164 24820 46170
rect 24768 46106 24820 46112
rect 24780 44849 24808 46106
rect 24766 44840 24822 44849
rect 24766 44775 24822 44784
rect 24872 42702 24900 47942
rect 24952 45824 25004 45830
rect 24952 45766 25004 45772
rect 24964 45665 24992 45766
rect 24950 45656 25006 45665
rect 24950 45591 25006 45600
rect 24952 43104 25004 43110
rect 24952 43046 25004 43052
rect 24860 42696 24912 42702
rect 24860 42638 24912 42644
rect 24860 42560 24912 42566
rect 24860 42502 24912 42508
rect 24872 42401 24900 42502
rect 24858 42392 24914 42401
rect 24858 42327 24914 42336
rect 24860 42016 24912 42022
rect 24860 41958 24912 41964
rect 24872 40730 24900 41958
rect 24860 40724 24912 40730
rect 24860 40666 24912 40672
rect 24768 40520 24820 40526
rect 24768 40462 24820 40468
rect 24780 39953 24808 40462
rect 24766 39944 24822 39953
rect 24766 39879 24822 39888
rect 24858 39128 24914 39137
rect 24858 39063 24914 39072
rect 24872 38962 24900 39063
rect 24860 38956 24912 38962
rect 24860 38898 24912 38904
rect 24964 38350 24992 43046
rect 25056 42022 25084 49694
rect 25136 49088 25188 49094
rect 25136 49030 25188 49036
rect 25148 42770 25176 49030
rect 25240 43194 25268 52838
rect 25596 52624 25648 52630
rect 25596 52566 25648 52572
rect 25504 51808 25556 51814
rect 25504 51750 25556 51756
rect 25516 51406 25544 51750
rect 25504 51400 25556 51406
rect 25502 51368 25504 51377
rect 25556 51368 25558 51377
rect 25502 51303 25558 51312
rect 25412 50720 25464 50726
rect 25412 50662 25464 50668
rect 25320 50176 25372 50182
rect 25320 50118 25372 50124
rect 25332 49842 25360 50118
rect 25320 49836 25372 49842
rect 25320 49778 25372 49784
rect 25332 49745 25360 49778
rect 25318 49736 25374 49745
rect 25318 49671 25374 49680
rect 25320 49224 25372 49230
rect 25320 49166 25372 49172
rect 25332 48929 25360 49166
rect 25318 48920 25374 48929
rect 25318 48855 25374 48864
rect 25320 48136 25372 48142
rect 25318 48104 25320 48113
rect 25372 48104 25374 48113
rect 25318 48039 25374 48048
rect 25320 44396 25372 44402
rect 25320 44338 25372 44344
rect 25332 43654 25360 44338
rect 25320 43648 25372 43654
rect 25320 43590 25372 43596
rect 25240 43166 25360 43194
rect 25136 42764 25188 42770
rect 25136 42706 25188 42712
rect 25044 42016 25096 42022
rect 25044 41958 25096 41964
rect 25332 41818 25360 43166
rect 25320 41812 25372 41818
rect 25320 41754 25372 41760
rect 25044 41744 25096 41750
rect 25044 41686 25096 41692
rect 25056 39506 25084 41686
rect 25320 41608 25372 41614
rect 25318 41576 25320 41585
rect 25372 41576 25374 41585
rect 25318 41511 25374 41520
rect 25136 41472 25188 41478
rect 25136 41414 25188 41420
rect 25320 41472 25372 41478
rect 25320 41414 25372 41420
rect 25148 39642 25176 41414
rect 25332 41138 25360 41414
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 25332 40769 25360 41074
rect 25318 40760 25374 40769
rect 25318 40695 25374 40704
rect 25424 40594 25452 50662
rect 25608 47274 25636 52566
rect 25688 51264 25740 51270
rect 25688 51206 25740 51212
rect 25516 47246 25636 47274
rect 25516 44878 25544 47246
rect 25596 47184 25648 47190
rect 25596 47126 25648 47132
rect 25504 44872 25556 44878
rect 25504 44814 25556 44820
rect 25504 44736 25556 44742
rect 25504 44678 25556 44684
rect 25516 44033 25544 44678
rect 25502 44024 25558 44033
rect 25502 43959 25558 43968
rect 25504 43648 25556 43654
rect 25504 43590 25556 43596
rect 25516 43217 25544 43590
rect 25502 43208 25558 43217
rect 25502 43143 25558 43152
rect 25504 43104 25556 43110
rect 25504 43046 25556 43052
rect 25516 42158 25544 43046
rect 25504 42152 25556 42158
rect 25504 42094 25556 42100
rect 25412 40588 25464 40594
rect 25412 40530 25464 40536
rect 25320 40384 25372 40390
rect 25320 40326 25372 40332
rect 25136 39636 25188 39642
rect 25136 39578 25188 39584
rect 25044 39500 25096 39506
rect 25044 39442 25096 39448
rect 25332 38962 25360 40326
rect 25516 39506 25544 42094
rect 25504 39500 25556 39506
rect 25504 39442 25556 39448
rect 25320 38956 25372 38962
rect 25320 38898 25372 38904
rect 25136 38752 25188 38758
rect 25136 38694 25188 38700
rect 24952 38344 25004 38350
rect 24688 38270 24808 38298
rect 24952 38286 25004 38292
rect 24676 38208 24728 38214
rect 24676 38150 24728 38156
rect 24688 38010 24716 38150
rect 24676 38004 24728 38010
rect 24676 37946 24728 37952
rect 24676 37188 24728 37194
rect 24676 37130 24728 37136
rect 24688 36786 24716 37130
rect 24676 36780 24728 36786
rect 24676 36722 24728 36728
rect 24780 36718 24808 38270
rect 24768 36712 24820 36718
rect 24768 36654 24820 36660
rect 25148 36106 25176 38694
rect 25332 38321 25360 38898
rect 25608 38554 25636 47126
rect 25700 41682 25728 51206
rect 25780 48544 25832 48550
rect 25780 48486 25832 48492
rect 25792 47666 25820 48486
rect 25780 47660 25832 47666
rect 25780 47602 25832 47608
rect 25792 47297 25820 47602
rect 25778 47288 25834 47297
rect 25778 47223 25834 47232
rect 25780 44872 25832 44878
rect 25780 44814 25832 44820
rect 25688 41676 25740 41682
rect 25688 41618 25740 41624
rect 25792 39030 25820 44814
rect 25780 39024 25832 39030
rect 25780 38966 25832 38972
rect 25884 38826 25912 53382
rect 25872 38820 25924 38826
rect 25872 38762 25924 38768
rect 25596 38548 25648 38554
rect 25596 38490 25648 38496
rect 25318 38312 25374 38321
rect 25318 38247 25374 38256
rect 25318 37496 25374 37505
rect 25318 37431 25374 37440
rect 25332 37262 25360 37431
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 25320 36780 25372 36786
rect 25320 36722 25372 36728
rect 25332 36689 25360 36722
rect 25318 36680 25374 36689
rect 25318 36615 25374 36624
rect 25320 36168 25372 36174
rect 25320 36110 25372 36116
rect 25136 36100 25188 36106
rect 25136 36042 25188 36048
rect 25332 35873 25360 36110
rect 25318 35864 25374 35873
rect 25318 35799 25374 35808
rect 25412 35624 25464 35630
rect 25412 35566 25464 35572
rect 25320 35488 25372 35494
rect 25320 35430 25372 35436
rect 25332 35086 25360 35430
rect 25320 35080 25372 35086
rect 25318 35048 25320 35057
rect 25372 35048 25374 35057
rect 25318 34983 25374 34992
rect 24952 34944 25004 34950
rect 24952 34886 25004 34892
rect 24676 34740 24728 34746
rect 24676 34682 24728 34688
rect 24584 33992 24636 33998
rect 24584 33934 24636 33940
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24492 32564 24544 32570
rect 24492 32506 24544 32512
rect 24400 31476 24452 31482
rect 24400 31418 24452 31424
rect 24216 31408 24268 31414
rect 24216 31350 24268 31356
rect 24228 30326 24256 31350
rect 24400 31136 24452 31142
rect 24400 31078 24452 31084
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 24228 30054 24256 30262
rect 24216 30048 24268 30054
rect 24268 30008 24348 30036
rect 24216 29990 24268 29996
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 24136 27713 24164 29106
rect 24320 28762 24348 30008
rect 24308 28756 24360 28762
rect 24308 28698 24360 28704
rect 24216 28484 24268 28490
rect 24216 28426 24268 28432
rect 24122 27704 24178 27713
rect 24228 27674 24256 28426
rect 24320 28218 24348 28698
rect 24308 28212 24360 28218
rect 24308 28154 24360 28160
rect 24122 27639 24178 27648
rect 24216 27668 24268 27674
rect 24216 27610 24268 27616
rect 24320 27606 24348 28154
rect 24308 27600 24360 27606
rect 24308 27542 24360 27548
rect 24412 26382 24440 31078
rect 24504 27470 24532 32506
rect 24596 29238 24624 33798
rect 24584 29232 24636 29238
rect 24584 29174 24636 29180
rect 24584 28416 24636 28422
rect 24584 28358 24636 28364
rect 24492 27464 24544 27470
rect 24492 27406 24544 27412
rect 24596 27130 24624 28358
rect 24688 28150 24716 34682
rect 24766 33416 24822 33425
rect 24766 33351 24822 33360
rect 24780 32570 24808 33351
rect 24768 32564 24820 32570
rect 24768 32506 24820 32512
rect 24964 31278 24992 34886
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25332 34241 25360 34546
rect 25318 34232 25374 34241
rect 25424 34202 25452 35566
rect 25318 34167 25320 34176
rect 25372 34167 25374 34176
rect 25412 34196 25464 34202
rect 25320 34138 25372 34144
rect 25412 34138 25464 34144
rect 25136 33924 25188 33930
rect 25136 33866 25188 33872
rect 25148 32026 25176 33866
rect 25424 33590 25452 34138
rect 25412 33584 25464 33590
rect 25412 33526 25464 33532
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 25332 32609 25360 32846
rect 25318 32600 25374 32609
rect 25318 32535 25374 32544
rect 25136 32020 25188 32026
rect 25136 31962 25188 31968
rect 25320 31816 25372 31822
rect 25318 31784 25320 31793
rect 25372 31784 25374 31793
rect 25318 31719 25374 31728
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 24952 31272 25004 31278
rect 24952 31214 25004 31220
rect 25332 30977 25360 31282
rect 25318 30968 25374 30977
rect 25318 30903 25320 30912
rect 25372 30903 25374 30912
rect 25320 30874 25372 30880
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 25044 30592 25096 30598
rect 25044 30534 25096 30540
rect 25136 30592 25188 30598
rect 25136 30534 25188 30540
rect 24858 28520 24914 28529
rect 24858 28455 24860 28464
rect 24912 28455 24914 28464
rect 24860 28426 24912 28432
rect 24676 28144 24728 28150
rect 24676 28086 24728 28092
rect 24676 28008 24728 28014
rect 24676 27950 24728 27956
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24596 26586 24624 26726
rect 24584 26580 24636 26586
rect 24584 26522 24636 26528
rect 24584 26444 24636 26450
rect 24584 26386 24636 26392
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 24032 25356 24084 25362
rect 24032 25298 24084 25304
rect 23940 25288 23992 25294
rect 23940 25230 23992 25236
rect 24032 25220 24084 25226
rect 24032 25162 24084 25168
rect 23846 23624 23902 23633
rect 23846 23559 23902 23568
rect 23860 23118 23888 23559
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23296 17060 23348 17066
rect 23296 17002 23348 17008
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22848 16658 23060 16674
rect 22848 16652 23072 16658
rect 22848 16646 23020 16652
rect 23020 16594 23072 16600
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22652 13320 22704 13326
rect 22652 13262 22704 13268
rect 22848 12850 22876 16186
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23308 15570 23336 17274
rect 23676 16114 23704 18634
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22940 13734 22968 14214
rect 22928 13728 22980 13734
rect 22928 13670 22980 13676
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23308 12850 23336 17002
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23400 14346 23428 16594
rect 23860 15026 23888 19722
rect 24044 18290 24072 25162
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 24320 23730 24348 24754
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24320 22778 24348 23666
rect 24596 23662 24624 26386
rect 24688 24750 24716 27950
rect 25056 27062 25084 30534
rect 25148 30394 25176 30534
rect 25136 30388 25188 30394
rect 25136 30330 25188 30336
rect 25318 30152 25374 30161
rect 25318 30087 25374 30096
rect 25332 29646 25360 30087
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25332 29306 25360 29582
rect 25516 29345 25544 30670
rect 25502 29336 25558 29345
rect 25320 29300 25372 29306
rect 25502 29271 25504 29280
rect 25320 29242 25372 29248
rect 25556 29271 25558 29280
rect 25504 29242 25556 29248
rect 25228 27396 25280 27402
rect 25228 27338 25280 27344
rect 25044 27056 25096 27062
rect 25044 26998 25096 27004
rect 24952 26512 25004 26518
rect 24952 26454 25004 26460
rect 24964 25498 24992 26454
rect 25044 26308 25096 26314
rect 25044 26250 25096 26256
rect 24952 25492 25004 25498
rect 24952 25434 25004 25440
rect 24860 25424 24912 25430
rect 24860 25366 24912 25372
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 24688 24342 24716 24686
rect 24676 24336 24728 24342
rect 24676 24278 24728 24284
rect 24872 24070 24900 25366
rect 24964 24886 24992 25434
rect 24952 24880 25004 24886
rect 24952 24822 25004 24828
rect 24950 24440 25006 24449
rect 24950 24375 25006 24384
rect 24964 24274 24992 24375
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 24596 23254 24624 23598
rect 24584 23248 24636 23254
rect 24584 23190 24636 23196
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 24858 21992 24914 22001
rect 24858 21927 24914 21936
rect 24216 21888 24268 21894
rect 24216 21830 24268 21836
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24228 16114 24256 21830
rect 24872 21010 24900 21927
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24766 19544 24822 19553
rect 24766 19479 24822 19488
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24412 18970 24440 19110
rect 24400 18964 24452 18970
rect 24400 18906 24452 18912
rect 24674 18728 24730 18737
rect 24674 18663 24730 18672
rect 24308 17536 24360 17542
rect 24308 17478 24360 17484
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 24320 15502 24348 17478
rect 24688 17134 24716 18663
rect 24780 18222 24808 19479
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24872 17678 24900 20810
rect 25056 20466 25084 26250
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25148 25265 25176 25774
rect 25134 25256 25190 25265
rect 25134 25191 25190 25200
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 24950 20360 25006 20369
rect 24950 20295 25006 20304
rect 24964 19922 24992 20295
rect 24952 19916 25004 19922
rect 24952 19858 25004 19864
rect 25240 19854 25268 27338
rect 25502 26888 25558 26897
rect 25502 26823 25558 26832
rect 25318 26072 25374 26081
rect 25318 26007 25374 26016
rect 25332 23730 25360 26007
rect 25516 25498 25544 26823
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 25516 24818 25544 25434
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 25332 22778 25360 23666
rect 25320 22772 25372 22778
rect 25320 22714 25372 22720
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24676 17128 24728 17134
rect 24676 17070 24728 17076
rect 24766 17096 24822 17105
rect 24766 17031 24822 17040
rect 24674 16280 24730 16289
rect 24674 16215 24730 16224
rect 24308 15496 24360 15502
rect 24308 15438 24360 15444
rect 23848 15020 23900 15026
rect 23848 14962 23900 14968
rect 24688 14958 24716 16215
rect 24780 16046 24808 17031
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24950 15464 25006 15473
rect 24950 15399 24952 15408
rect 25004 15399 25006 15408
rect 24952 15370 25004 15376
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 25134 14648 25190 14657
rect 25134 14583 25190 14592
rect 23388 14340 23440 14346
rect 23388 14282 23440 14288
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22100 11620 22152 11626
rect 22100 11562 22152 11568
rect 21744 10526 21864 10554
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21744 8974 21772 10406
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21100 6322 21128 7686
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21284 4622 21312 8366
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21180 4004 21232 4010
rect 21180 3946 21232 3952
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20456 2774 20760 2802
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 20456 800 20484 2774
rect 20824 800 20852 2790
rect 21192 800 21220 3946
rect 21560 800 21588 5714
rect 21836 5234 21864 10526
rect 22008 8356 22060 8362
rect 22008 8298 22060 8304
rect 22020 7410 22048 8298
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21928 800 21956 6190
rect 22020 3398 22048 6666
rect 22112 6322 22140 11562
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22560 10192 22612 10198
rect 22560 10134 22612 10140
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22112 4049 22140 4082
rect 22098 4040 22154 4049
rect 22098 3975 22154 3984
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22204 2417 22232 7278
rect 22190 2408 22246 2417
rect 22190 2343 22246 2352
rect 22296 800 22324 7278
rect 22388 5250 22416 8366
rect 22572 5710 22600 10134
rect 23308 9994 23336 12310
rect 23296 9988 23348 9994
rect 23296 9930 23348 9936
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22652 6384 22704 6390
rect 22652 6326 22704 6332
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22388 5222 22600 5250
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22374 4040 22430 4049
rect 22374 3975 22430 3984
rect 22388 3942 22416 3975
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22480 2854 22508 5102
rect 22572 3233 22600 5222
rect 22558 3224 22614 3233
rect 22558 3159 22614 3168
rect 22468 2848 22520 2854
rect 22468 2790 22520 2796
rect 22664 800 22692 6326
rect 22756 4690 22784 9318
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22836 9104 22888 9110
rect 22836 9046 22888 9052
rect 22848 6798 22876 9046
rect 23400 8974 23428 14010
rect 25148 14006 25176 14583
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 24766 13832 24822 13841
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23296 8832 23348 8838
rect 23296 8774 23348 8780
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 22836 6180 22888 6186
rect 22836 6122 22888 6128
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 22848 3738 22876 6122
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23308 4622 23336 8774
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23400 4865 23428 7890
rect 23492 7886 23520 8774
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23386 4856 23442 4865
rect 23386 4791 23442 4800
rect 23296 4616 23348 4622
rect 23296 4558 23348 4564
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 22848 2530 22876 3334
rect 23584 3126 23612 3334
rect 23572 3120 23624 3126
rect 23572 3062 23624 3068
rect 23388 2916 23440 2922
rect 23388 2858 23440 2864
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22848 2502 23060 2530
rect 23032 800 23060 2502
rect 23400 800 23428 2858
rect 23768 800 23796 13806
rect 24766 13767 24822 13776
rect 24780 12782 24808 13767
rect 25688 13252 25740 13258
rect 25688 13194 25740 13200
rect 25700 13025 25728 13194
rect 25686 13016 25742 13025
rect 25686 12951 25742 12960
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23860 9586 23888 11018
rect 23940 10464 23992 10470
rect 23940 10406 23992 10412
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23848 9444 23900 9450
rect 23848 9386 23900 9392
rect 23860 4146 23888 9386
rect 23952 8498 23980 10406
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23940 7404 23992 7410
rect 23940 7346 23992 7352
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23952 3641 23980 7346
rect 24044 6322 24072 9862
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 24136 5234 24164 7686
rect 24504 6914 24532 11494
rect 24596 8974 24624 12582
rect 25134 12200 25190 12209
rect 25134 12135 25190 12144
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24766 11384 24822 11393
rect 24766 11319 24822 11328
rect 24780 10606 24808 11319
rect 24768 10600 24820 10606
rect 24674 10568 24730 10577
rect 24768 10542 24820 10548
rect 24674 10503 24730 10512
rect 24688 9518 24716 10503
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24872 7886 24900 12038
rect 25148 11830 25176 12135
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24964 9761 24992 9998
rect 24950 9752 25006 9761
rect 24950 9687 25006 9696
rect 25134 8936 25190 8945
rect 25134 8871 25190 8880
rect 25148 8566 25176 8871
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24860 7880 24912 7886
rect 24860 7822 24912 7828
rect 24964 6914 24992 8366
rect 25134 8120 25190 8129
rect 25134 8055 25190 8064
rect 25148 7478 25176 8055
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 25134 7304 25190 7313
rect 25134 7239 25190 7248
rect 24504 6886 24716 6914
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 23938 3632 23994 3641
rect 23938 3567 23994 3576
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24136 800 24164 3334
rect 24688 3194 24716 6886
rect 24872 6886 24992 6914
rect 24766 5672 24822 5681
rect 24766 5607 24822 5616
rect 24780 5166 24808 5607
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24872 4758 24900 6886
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 24964 6497 24992 6666
rect 24950 6488 25006 6497
rect 24950 6423 25006 6432
rect 25148 6390 25176 7239
rect 25136 6384 25188 6390
rect 25136 6326 25188 6332
rect 24860 4752 24912 4758
rect 24860 4694 24912 4700
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 13188 734 13400 762
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 24964 785 24992 3674
rect 25320 2440 25372 2446
rect 25320 2382 25372 2388
rect 25332 1601 25360 2382
rect 25318 1592 25374 1601
rect 25318 1527 25374 1536
rect 24950 776 25006 785
rect 24950 711 25006 720
<< via2 >>
rect 1306 52944 1362 53000
rect 1306 50496 1362 50552
rect 2778 55392 2834 55448
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 1306 48068 1362 48104
rect 1306 48048 1308 48068
rect 1308 48048 1360 48068
rect 1360 48048 1362 48068
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 1306 45620 1362 45656
rect 1306 45600 1308 45620
rect 1308 45600 1360 45620
rect 1360 45600 1362 45620
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 1306 43152 1362 43208
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 1306 40704 1362 40760
rect 1306 38292 1308 38312
rect 1308 38292 1360 38312
rect 1360 38292 1362 38312
rect 1306 38256 1362 38292
rect 1306 33360 1362 33416
rect 1306 30912 1362 30968
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 1306 36488 1362 36544
rect 1582 34176 1638 34232
rect 1306 31864 1362 31920
rect 1306 29552 1362 29608
rect 1306 27240 1362 27296
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 1766 35808 1822 35864
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 1306 24928 1362 24984
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 1306 28464 1362 28520
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 1306 23604 1308 23624
rect 1308 23604 1360 23624
rect 1360 23604 1362 23624
rect 1306 23568 1362 23604
rect 2778 26016 2834 26072
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 938 22616 994 22672
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 1306 21120 1362 21176
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 1306 18672 1362 18728
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 1306 15680 1362 15736
rect 1766 13368 1822 13424
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2502 16496 2558 16552
rect 1306 16224 1362 16280
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 1306 13812 1308 13832
rect 1308 13812 1360 13832
rect 1360 13812 1362 13832
rect 1306 13776 1362 13812
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3054 8880 3110 8936
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3054 6432 3110 6488
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3146 4020 3148 4040
rect 3148 4020 3200 4040
rect 3200 4020 3202 4040
rect 3146 3984 3202 4020
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 4066 16496 4122 16552
rect 3882 11600 3938 11656
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 2870 1536 2926 1592
rect 5906 6296 5962 6352
rect 7102 35672 7158 35728
rect 7286 38256 7342 38312
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 8482 42472 8538 42528
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7654 40432 7710 40488
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 8206 38256 8262 38312
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 9678 44684 9680 44704
rect 9680 44684 9732 44704
rect 9732 44684 9734 44704
rect 9678 44648 9734 44684
rect 9862 36896 9918 36952
rect 8758 35808 8814 35864
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 9402 44240 9458 44296
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 9586 40452 9642 40488
rect 9586 40432 9588 40452
rect 9588 40432 9640 40452
rect 9640 40432 9642 40452
rect 9586 38836 9588 38856
rect 9588 38836 9640 38856
rect 9640 38836 9642 38856
rect 9586 38800 9642 38836
rect 10414 42508 10416 42528
rect 10416 42508 10468 42528
rect 10468 42508 10470 42528
rect 10414 42472 10470 42508
rect 9770 36760 9826 36816
rect 9954 36760 10010 36816
rect 8850 33904 8906 33960
rect 9402 33904 9458 33960
rect 9632 33924 9688 33926
rect 9632 33872 9680 33924
rect 9680 33872 9688 33924
rect 9632 33870 9688 33872
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 7010 5616 7066 5672
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 10598 41248 10654 41304
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12254 45228 12256 45248
rect 12256 45228 12308 45248
rect 12308 45228 12310 45248
rect 12254 45192 12310 45228
rect 11334 41248 11390 41304
rect 10598 30640 10654 30696
rect 10874 31728 10930 31784
rect 12070 37168 12126 37224
rect 12070 33632 12126 33688
rect 11058 21684 11114 21720
rect 11058 21664 11060 21684
rect 11060 21664 11112 21684
rect 11112 21664 11114 21684
rect 11610 24112 11666 24168
rect 11702 21528 11758 21584
rect 11702 21020 11704 21040
rect 11704 21020 11756 21040
rect 11756 21020 11758 21040
rect 11702 20984 11758 21020
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 11518 44512 11574 44568
rect 11334 38256 11390 38312
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 9494 16496 9550 16552
rect 11426 38120 11482 38176
rect 12438 40452 12494 40488
rect 12438 40432 12440 40452
rect 12440 40432 12492 40452
rect 12492 40432 12494 40452
rect 12162 36216 12218 36272
rect 12438 37712 12494 37768
rect 14002 52536 14058 52592
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 13450 40704 13506 40760
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12622 38392 12678 38448
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12714 36624 12770 36680
rect 12438 35808 12494 35864
rect 10874 19116 10876 19136
rect 10876 19116 10928 19136
rect 10928 19116 10930 19136
rect 10874 19080 10930 19116
rect 11058 18164 11060 18184
rect 11060 18164 11112 18184
rect 11112 18164 11114 18184
rect 11058 18128 11114 18164
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 13450 38392 13506 38448
rect 13450 35808 13506 35864
rect 13358 35400 13414 35456
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 13358 35128 13414 35184
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12622 30912 12678 30968
rect 12162 23976 12218 24032
rect 12162 22752 12218 22808
rect 12162 19352 12218 19408
rect 12346 19216 12402 19272
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 13818 38256 13874 38312
rect 14462 52944 14518 53000
rect 14370 38800 14426 38856
rect 13818 36236 13874 36272
rect 13818 36216 13820 36236
rect 13820 36216 13872 36236
rect 13872 36216 13874 36236
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 14002 35284 14058 35320
rect 14002 35264 14004 35284
rect 14004 35264 14056 35284
rect 14056 35264 14058 35284
rect 14002 33360 14058 33416
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 13542 30504 13598 30560
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 14370 30252 14426 30288
rect 14370 30232 14372 30252
rect 14372 30232 14424 30252
rect 14424 30232 14426 30252
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12990 19252 12992 19272
rect 12992 19252 13044 19272
rect 13044 19252 13046 19272
rect 12990 19216 13046 19252
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12714 17856 12770 17912
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12806 17876 12862 17912
rect 12806 17856 12808 17876
rect 12808 17856 12860 17876
rect 12860 17856 12862 17876
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12806 15952 12862 16008
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 13818 21800 13874 21836
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 13818 18128 13874 18184
rect 14186 16108 14242 16144
rect 14186 16088 14188 16108
rect 14188 16088 14240 16108
rect 14240 16088 14242 16108
rect 15198 30368 15254 30424
rect 15198 28364 15200 28384
rect 15200 28364 15252 28384
rect 15252 28364 15254 28384
rect 15198 28328 15254 28364
rect 17038 53932 17040 53952
rect 17040 53932 17092 53952
rect 17092 53932 17094 53952
rect 17038 53896 17094 53932
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 16394 52536 16450 52592
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 15842 40432 15898 40488
rect 16026 38700 16028 38720
rect 16028 38700 16080 38720
rect 16080 38700 16082 38720
rect 16026 38664 16082 38700
rect 15750 35980 15752 36000
rect 15752 35980 15804 36000
rect 15804 35980 15806 36000
rect 15750 35944 15806 35980
rect 15382 29008 15438 29064
rect 15382 27240 15438 27296
rect 15658 32816 15714 32872
rect 15750 29008 15806 29064
rect 14554 19252 14556 19272
rect 14556 19252 14608 19272
rect 14608 19252 14610 19272
rect 14554 19216 14610 19252
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 14554 36760 14610 36816
rect 14462 34448 14518 34504
rect 15658 53896 15714 53952
rect 15290 38700 15292 38720
rect 15292 38700 15344 38720
rect 15344 38700 15346 38720
rect 15290 38664 15346 38700
rect 14738 29008 14794 29064
rect 14738 21836 14740 21856
rect 14740 21836 14792 21856
rect 14792 21836 14794 21856
rect 14738 21800 14794 21836
rect 14554 21392 14610 21448
rect 14646 20168 14702 20224
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 16394 38120 16450 38176
rect 16762 36780 16818 36816
rect 16762 36760 16764 36780
rect 16764 36760 16816 36780
rect 16816 36760 16818 36780
rect 17222 38256 17278 38312
rect 16486 30368 16542 30424
rect 15934 28212 15990 28248
rect 15934 28192 15936 28212
rect 15936 28192 15988 28212
rect 15988 28192 15990 28212
rect 16026 20712 16082 20768
rect 16394 29008 16450 29064
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 18786 47676 18788 47696
rect 18788 47676 18840 47696
rect 18840 47676 18842 47696
rect 18786 47640 18842 47676
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17590 39344 17646 39400
rect 17590 38664 17646 38720
rect 17590 38528 17646 38584
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17774 37204 17776 37224
rect 17776 37204 17828 37224
rect 17828 37204 17830 37224
rect 17774 37168 17830 37204
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 18418 38836 18420 38856
rect 18420 38836 18472 38856
rect 18472 38836 18474 38856
rect 18418 38800 18474 38836
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 16394 16244 16450 16280
rect 16394 16224 16396 16244
rect 16396 16224 16448 16244
rect 16448 16224 16450 16244
rect 17222 27396 17278 27432
rect 17222 27376 17224 27396
rect 17224 27376 17276 27396
rect 17276 27376 17278 27396
rect 17222 26288 17278 26344
rect 18694 37712 18750 37768
rect 18878 38528 18934 38584
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 19522 44240 19578 44296
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 18142 30796 18198 30832
rect 18142 30776 18144 30796
rect 18144 30776 18196 30796
rect 18196 30776 18198 30796
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 18234 29708 18290 29744
rect 18234 29688 18236 29708
rect 18236 29688 18288 29708
rect 18288 29688 18290 29708
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 18326 28464 18382 28520
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 18786 37304 18842 37360
rect 18970 36644 19026 36680
rect 18970 36624 18972 36644
rect 18972 36624 19024 36644
rect 19024 36624 19026 36644
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 18326 26288 18382 26344
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17314 20596 17370 20632
rect 17314 20576 17316 20596
rect 17316 20576 17368 20596
rect 17368 20576 17370 20596
rect 16302 3576 16358 3632
rect 17774 19896 17830 19952
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17958 23740 17960 23760
rect 17960 23740 18012 23760
rect 18012 23740 18014 23760
rect 17958 23704 18014 23740
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17222 19896 17278 19952
rect 15658 2624 15714 2680
rect 17590 18828 17646 18864
rect 17590 18808 17592 18828
rect 17592 18808 17644 18828
rect 17644 18808 17646 18828
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18326 18672 18382 18728
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18510 18264 18566 18320
rect 17866 17584 17922 17640
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17498 11892 17554 11928
rect 17498 11872 17500 11892
rect 17500 11872 17552 11892
rect 17552 11872 17554 11892
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 20442 47096 20498 47152
rect 19430 38412 19486 38448
rect 19430 38392 19432 38412
rect 19432 38392 19484 38412
rect 19484 38392 19486 38412
rect 19062 30252 19118 30288
rect 19062 30232 19064 30252
rect 19064 30232 19116 30252
rect 19116 30232 19118 30252
rect 18602 14456 18658 14512
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 19430 37984 19486 38040
rect 19706 37168 19762 37224
rect 20810 44240 20866 44296
rect 20534 40296 20590 40352
rect 20442 39364 20498 39400
rect 20442 39344 20444 39364
rect 20444 39344 20496 39364
rect 20496 39344 20498 39364
rect 20442 38120 20498 38176
rect 20258 37868 20314 37904
rect 20258 37848 20260 37868
rect 20260 37848 20312 37868
rect 20312 37848 20314 37868
rect 20442 37324 20498 37360
rect 20442 37304 20444 37324
rect 20444 37304 20496 37324
rect 20496 37304 20498 37324
rect 19706 36216 19762 36272
rect 19522 29300 19578 29336
rect 19522 29280 19524 29300
rect 19524 29280 19576 29300
rect 19576 29280 19578 29300
rect 19982 31220 19984 31240
rect 19984 31220 20036 31240
rect 20036 31220 20038 31240
rect 19982 31184 20038 31220
rect 19246 24792 19302 24848
rect 20442 30932 20498 30968
rect 20442 30912 20444 30932
rect 20444 30912 20496 30932
rect 20496 30912 20498 30932
rect 20258 28212 20314 28248
rect 20258 28192 20260 28212
rect 20260 28192 20312 28212
rect 20312 28192 20314 28212
rect 21914 46552 21970 46608
rect 21638 43052 21640 43072
rect 21640 43052 21692 43072
rect 21692 43052 21694 43072
rect 21638 43016 21694 43052
rect 21454 40588 21510 40624
rect 21454 40568 21456 40588
rect 21456 40568 21508 40588
rect 21508 40568 21510 40588
rect 21362 40432 21418 40488
rect 21638 40452 21694 40488
rect 21638 40432 21640 40452
rect 21640 40432 21692 40452
rect 21692 40432 21694 40452
rect 21822 40432 21878 40488
rect 19982 21140 20038 21176
rect 19982 21120 19984 21140
rect 19984 21120 20036 21140
rect 20036 21120 20038 21140
rect 21086 32272 21142 32328
rect 21454 32816 21510 32872
rect 22742 53932 22744 53952
rect 22744 53932 22796 53952
rect 22796 53932 22798 53952
rect 22742 53896 22798 53932
rect 23386 56072 23442 56128
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 24490 55392 24546 55448
rect 24766 54576 24822 54632
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22650 45484 22706 45520
rect 22650 45464 22652 45484
rect 22652 45464 22704 45484
rect 22704 45464 22706 45484
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 21914 32564 21970 32600
rect 21914 32544 21916 32564
rect 21916 32544 21968 32564
rect 21968 32544 21970 32564
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 21454 29164 21510 29200
rect 21454 29144 21456 29164
rect 21456 29144 21508 29164
rect 21508 29144 21510 29164
rect 20166 3984 20222 4040
rect 22466 37168 22522 37224
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 23478 45600 23534 45656
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 23110 40604 23112 40624
rect 23112 40604 23164 40624
rect 23164 40604 23166 40624
rect 23110 40568 23166 40604
rect 22926 40468 22928 40488
rect 22928 40468 22980 40488
rect 22980 40468 22982 40488
rect 22926 40432 22982 40468
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 23386 40296 23442 40352
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22466 34856 22522 34912
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 24674 52536 24730 52592
rect 24766 49136 24822 49192
rect 24766 47776 24822 47832
rect 25226 51856 25282 51912
rect 25318 51176 25374 51232
rect 24858 46436 24914 46472
rect 24858 46416 24860 46436
rect 24860 46416 24912 46436
rect 24912 46416 24914 46436
rect 24766 45736 24822 45792
rect 24766 44376 24822 44432
rect 24674 43696 24730 43752
rect 23662 37168 23718 37224
rect 23938 36760 23994 36816
rect 24766 40976 24822 41032
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22742 32852 22744 32872
rect 22744 32852 22796 32872
rect 22796 32852 22798 32872
rect 22742 32816 22798 32852
rect 22650 32272 22706 32328
rect 22374 29280 22430 29336
rect 23202 32308 23204 32328
rect 23204 32308 23256 32328
rect 23256 32308 23258 32328
rect 23202 32272 23258 32308
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 24030 37168 24086 37224
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 21638 15544 21694 15600
rect 22098 19216 22154 19272
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 23294 22752 23350 22808
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 24122 28736 24178 28792
rect 23386 23296 23442 23352
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23386 21120 23442 21176
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23386 17856 23442 17912
rect 24950 53760 25006 53816
rect 24766 52128 24822 52184
rect 25042 52944 25098 53000
rect 25042 50496 25098 50552
rect 24582 40332 24584 40352
rect 24584 40332 24636 40352
rect 24636 40332 24638 40352
rect 24582 40296 24638 40332
rect 24766 46416 24822 46472
rect 24766 44784 24822 44840
rect 24950 45600 25006 45656
rect 24858 42336 24914 42392
rect 24766 39888 24822 39944
rect 24858 39072 24914 39128
rect 25502 51348 25504 51368
rect 25504 51348 25556 51368
rect 25556 51348 25558 51368
rect 25502 51312 25558 51348
rect 25318 49680 25374 49736
rect 25318 48864 25374 48920
rect 25318 48084 25320 48104
rect 25320 48084 25372 48104
rect 25372 48084 25374 48104
rect 25318 48048 25374 48084
rect 25318 41556 25320 41576
rect 25320 41556 25372 41576
rect 25372 41556 25374 41576
rect 25318 41520 25374 41556
rect 25318 40704 25374 40760
rect 25502 43968 25558 44024
rect 25502 43152 25558 43208
rect 25778 47232 25834 47288
rect 25318 38256 25374 38312
rect 25318 37440 25374 37496
rect 25318 36624 25374 36680
rect 25318 35808 25374 35864
rect 25318 35028 25320 35048
rect 25320 35028 25372 35048
rect 25372 35028 25374 35048
rect 25318 34992 25374 35028
rect 24122 27648 24178 27704
rect 24766 33360 24822 33416
rect 25318 34196 25374 34232
rect 25318 34176 25320 34196
rect 25320 34176 25372 34196
rect 25372 34176 25374 34196
rect 25318 32544 25374 32600
rect 25318 31764 25320 31784
rect 25320 31764 25372 31784
rect 25372 31764 25374 31784
rect 25318 31728 25374 31764
rect 25318 30932 25374 30968
rect 25318 30912 25320 30932
rect 25320 30912 25372 30932
rect 25372 30912 25374 30932
rect 24858 28484 24914 28520
rect 24858 28464 24860 28484
rect 24860 28464 24912 28484
rect 24912 28464 24914 28484
rect 23846 23568 23902 23624
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 25318 30096 25374 30152
rect 25502 29300 25558 29336
rect 25502 29280 25504 29300
rect 25504 29280 25556 29300
rect 25556 29280 25558 29300
rect 24950 24384 25006 24440
rect 24858 21936 24914 21992
rect 24766 19488 24822 19544
rect 24674 18672 24730 18728
rect 25134 25200 25190 25256
rect 24950 20304 25006 20360
rect 25502 26832 25558 26888
rect 25318 26016 25374 26072
rect 24766 17040 24822 17096
rect 24674 16224 24730 16280
rect 24950 15428 25006 15464
rect 24950 15408 24952 15428
rect 24952 15408 25004 15428
rect 25004 15408 25006 15428
rect 25134 14592 25190 14648
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 24766 38256 24822 38312
rect 25318 50496 25374 50552
rect 25318 49816 25374 49872
rect 25318 48456 25374 48512
rect 25502 47096 25558 47152
rect 24950 39616 25006 39672
rect 24950 36896 25006 36952
rect 24766 35536 24822 35592
rect 24858 28056 24914 28112
rect 24674 26696 24730 26752
rect 24490 21256 24546 21312
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22098 3984 22154 4040
rect 22190 2352 22246 2408
rect 22374 3984 22430 4040
rect 22558 3168 22614 3224
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 23386 4800 23442 4856
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24766 13776 24822 13832
rect 25686 12960 25742 13016
rect 25134 12144 25190 12200
rect 24766 11328 24822 11384
rect 24674 10512 24730 10568
rect 24950 9696 25006 9752
rect 25134 8880 25190 8936
rect 25134 8064 25190 8120
rect 25134 7248 25190 7304
rect 23938 3576 23994 3632
rect 24766 5616 24822 5672
rect 24950 6432 25006 6488
rect 25318 1536 25374 1592
rect 24950 720 25006 776
<< metal3 >>
rect 26200 56266 27000 56296
rect 23430 56206 27000 56266
rect 23430 56133 23490 56206
rect 26200 56176 27000 56206
rect 23381 56128 23490 56133
rect 23381 56072 23386 56128
rect 23442 56072 23490 56128
rect 23381 56070 23490 56072
rect 23381 56067 23447 56070
rect 0 55450 800 55480
rect 2773 55450 2839 55453
rect 0 55448 2839 55450
rect 0 55392 2778 55448
rect 2834 55392 2839 55448
rect 0 55390 2839 55392
rect 0 55360 800 55390
rect 2773 55387 2839 55390
rect 24485 55450 24551 55453
rect 26200 55450 27000 55480
rect 24485 55448 27000 55450
rect 24485 55392 24490 55448
rect 24546 55392 27000 55448
rect 24485 55390 27000 55392
rect 24485 55387 24551 55390
rect 26200 55360 27000 55390
rect 24761 54634 24827 54637
rect 26200 54634 27000 54664
rect 24761 54632 27000 54634
rect 24761 54576 24766 54632
rect 24822 54576 27000 54632
rect 24761 54574 27000 54576
rect 24761 54571 24827 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 17033 53954 17099 53957
rect 22737 53956 22803 53957
rect 17166 53954 17172 53956
rect 17033 53952 17172 53954
rect 17033 53896 17038 53952
rect 17094 53896 17172 53952
rect 17033 53894 17172 53896
rect 17033 53891 17099 53894
rect 17166 53892 17172 53894
rect 17236 53892 17242 53956
rect 22686 53954 22692 53956
rect 22646 53894 22692 53954
rect 22756 53952 22803 53956
rect 22798 53896 22803 53952
rect 22686 53892 22692 53894
rect 22756 53892 22803 53896
rect 22737 53891 22803 53892
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 24945 53818 25011 53821
rect 26200 53818 27000 53848
rect 24945 53816 27000 53818
rect 24945 53760 24950 53816
rect 25006 53760 27000 53816
rect 24945 53758 27000 53760
rect 24945 53755 25011 53758
rect 26200 53728 27000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 0 53002 800 53032
rect 1301 53002 1367 53005
rect 0 53000 1367 53002
rect 0 52944 1306 53000
rect 1362 52944 1367 53000
rect 0 52942 1367 52944
rect 0 52912 800 52942
rect 1301 52939 1367 52942
rect 14457 53002 14523 53005
rect 14590 53002 14596 53004
rect 14457 53000 14596 53002
rect 14457 52944 14462 53000
rect 14518 52944 14596 53000
rect 14457 52942 14596 52944
rect 14457 52939 14523 52942
rect 14590 52940 14596 52942
rect 14660 52940 14666 53004
rect 25037 53002 25103 53005
rect 26200 53002 27000 53032
rect 25037 53000 27000 53002
rect 25037 52944 25042 53000
rect 25098 52944 27000 53000
rect 25037 52942 27000 52944
rect 25037 52939 25103 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 13997 52596 14063 52597
rect 16389 52596 16455 52597
rect 13997 52592 14044 52596
rect 14108 52594 14114 52596
rect 13997 52536 14002 52592
rect 13997 52532 14044 52536
rect 14108 52534 14154 52594
rect 16389 52592 16436 52596
rect 16500 52594 16506 52596
rect 16389 52536 16394 52592
rect 14108 52532 14114 52534
rect 16389 52532 16436 52536
rect 16500 52534 16546 52594
rect 16500 52532 16506 52534
rect 13997 52531 14063 52532
rect 16389 52531 16455 52532
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 24761 52186 24827 52189
rect 26200 52186 27000 52216
rect 24761 52184 27000 52186
rect 24761 52128 24766 52184
rect 24822 52128 27000 52184
rect 24761 52126 27000 52128
rect 24761 52123 24827 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 25497 51370 25563 51373
rect 26200 51370 27000 51400
rect 25497 51368 27000 51370
rect 25497 51312 25502 51368
rect 25558 51312 27000 51368
rect 25497 51310 27000 51312
rect 25497 51307 25563 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 0 50554 800 50584
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 1301 50554 1367 50557
rect 0 50552 1367 50554
rect 0 50496 1306 50552
rect 1362 50496 1367 50552
rect 0 50494 1367 50496
rect 0 50464 800 50494
rect 1301 50491 1367 50494
rect 25037 50554 25103 50557
rect 26200 50554 27000 50584
rect 25313 50552 27000 50554
rect 25313 50496 25318 50552
rect 25374 50496 27000 50552
rect 25313 50494 27000 50496
rect 25313 50491 25379 50494
rect 26200 50464 27000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25313 49738 25379 49741
rect 26200 49738 27000 49768
rect 25313 49736 27000 49738
rect 25313 49680 25318 49736
rect 25374 49680 27000 49736
rect 25313 49678 27000 49680
rect 25313 49675 25379 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25313 48922 25379 48925
rect 26200 48922 27000 48952
rect 25313 48920 27000 48922
rect 25313 48864 25318 48920
rect 25374 48864 27000 48920
rect 25313 48862 27000 48864
rect 25313 48859 25379 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 0 48106 800 48136
rect 1301 48106 1367 48109
rect 0 48104 1367 48106
rect 0 48048 1306 48104
rect 1362 48048 1367 48104
rect 0 48046 1367 48048
rect 0 48016 800 48046
rect 1301 48043 1367 48046
rect 25313 48106 25379 48109
rect 26200 48106 27000 48136
rect 25313 48104 27000 48106
rect 25313 48048 25318 48104
rect 25374 48048 27000 48104
rect 25313 48046 27000 48048
rect 25313 48043 25379 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 18781 47700 18847 47701
rect 18781 47696 18828 47700
rect 18892 47698 18898 47700
rect 18781 47640 18786 47696
rect 18781 47636 18828 47640
rect 18892 47638 18938 47698
rect 18892 47636 18898 47638
rect 18781 47635 18847 47636
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25773 47290 25839 47293
rect 26200 47290 27000 47320
rect 25773 47288 27000 47290
rect 25773 47232 25778 47288
rect 25834 47232 27000 47288
rect 25773 47230 27000 47232
rect 25773 47227 25839 47230
rect 26200 47200 27000 47230
rect 19190 47092 19196 47156
rect 19260 47154 19266 47156
rect 20437 47154 20503 47157
rect 19260 47152 20503 47154
rect 19260 47096 20442 47152
rect 20498 47096 20503 47152
rect 19260 47094 20503 47096
rect 19260 47092 19266 47094
rect 20437 47091 20503 47094
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 21909 46612 21975 46613
rect 21909 46608 21956 46612
rect 22020 46610 22026 46612
rect 21909 46552 21914 46608
rect 21909 46548 21956 46552
rect 22020 46550 22066 46610
rect 22020 46548 22026 46550
rect 21909 46547 21975 46548
rect 24761 46474 24827 46477
rect 26200 46474 27000 46504
rect 24761 46472 27000 46474
rect 24761 46416 24766 46472
rect 24822 46416 27000 46472
rect 24761 46414 27000 46416
rect 24761 46411 24827 46414
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 7946 45728 8262 45729
rect 0 45658 800 45688
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 1301 45658 1367 45661
rect 0 45656 1367 45658
rect 0 45600 1306 45656
rect 1362 45600 1367 45656
rect 0 45598 1367 45600
rect 0 45568 800 45598
rect 1301 45595 1367 45598
rect 23473 45658 23539 45661
rect 23606 45658 23612 45660
rect 23473 45656 23612 45658
rect 23473 45600 23478 45656
rect 23534 45600 23612 45656
rect 23473 45598 23612 45600
rect 23473 45595 23539 45598
rect 23606 45596 23612 45598
rect 23676 45596 23682 45660
rect 24945 45658 25011 45661
rect 26200 45658 27000 45688
rect 24945 45656 27000 45658
rect 24945 45600 24950 45656
rect 25006 45600 27000 45656
rect 24945 45598 27000 45600
rect 24945 45595 25011 45598
rect 26200 45568 27000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 24761 44842 24827 44845
rect 26200 44842 27000 44872
rect 24761 44840 27000 44842
rect 24761 44784 24766 44840
rect 24822 44784 27000 44840
rect 24761 44782 27000 44784
rect 24761 44779 24827 44782
rect 26200 44752 27000 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 11513 44570 11579 44573
rect 12382 44570 12388 44572
rect 11513 44568 12388 44570
rect 11513 44512 11518 44568
rect 11574 44512 12388 44568
rect 11513 44510 12388 44512
rect 11513 44507 11579 44510
rect 12382 44508 12388 44510
rect 12452 44508 12458 44572
rect 9397 44298 9463 44301
rect 9622 44298 9628 44300
rect 9397 44296 9628 44298
rect 9397 44240 9402 44296
rect 9458 44240 9628 44296
rect 9397 44238 9628 44240
rect 9397 44235 9463 44238
rect 9622 44236 9628 44238
rect 9692 44236 9698 44300
rect 20662 44236 20668 44300
rect 20732 44298 20738 44300
rect 20805 44298 20871 44301
rect 20732 44296 20871 44298
rect 20732 44240 20810 44296
rect 20866 44240 20871 44296
rect 20732 44238 20871 44240
rect 20732 44236 20738 44238
rect 20805 44235 20871 44238
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 25497 44026 25563 44029
rect 26200 44026 27000 44056
rect 25497 44024 27000 44026
rect 25497 43968 25502 44024
rect 25558 43968 27000 44024
rect 25497 43966 27000 43968
rect 25497 43963 25563 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 0 43210 800 43240
rect 1301 43210 1367 43213
rect 0 43208 1367 43210
rect 0 43152 1306 43208
rect 1362 43152 1367 43208
rect 0 43150 1367 43152
rect 0 43120 800 43150
rect 1301 43147 1367 43150
rect 25497 43210 25563 43213
rect 26200 43210 27000 43240
rect 25497 43208 27000 43210
rect 25497 43152 25502 43208
rect 25558 43152 27000 43208
rect 25497 43150 27000 43152
rect 25497 43147 25563 43150
rect 26200 43120 27000 43150
rect 21633 43076 21699 43077
rect 21582 43012 21588 43076
rect 21652 43074 21699 43076
rect 21652 43072 21744 43074
rect 21694 43016 21744 43072
rect 21652 43014 21744 43016
rect 21652 43012 21699 43014
rect 21633 43011 21699 43012
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 8477 42530 8543 42533
rect 9254 42530 9260 42532
rect 8477 42528 9260 42530
rect 8477 42472 8482 42528
rect 8538 42472 9260 42528
rect 8477 42470 9260 42472
rect 8477 42467 8543 42470
rect 9254 42468 9260 42470
rect 9324 42468 9330 42532
rect 10409 42530 10475 42533
rect 10542 42530 10548 42532
rect 10409 42528 10548 42530
rect 10409 42472 10414 42528
rect 10470 42472 10548 42528
rect 10409 42470 10548 42472
rect 10409 42467 10475 42470
rect 10542 42468 10548 42470
rect 10612 42468 10618 42532
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 24853 42394 24919 42397
rect 26200 42394 27000 42424
rect 24853 42392 27000 42394
rect 24853 42336 24858 42392
rect 24914 42336 27000 42392
rect 24853 42334 27000 42336
rect 24853 42331 24919 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 25313 41578 25379 41581
rect 26200 41578 27000 41608
rect 25313 41576 27000 41578
rect 25313 41520 25318 41576
rect 25374 41520 27000 41576
rect 25313 41518 27000 41520
rect 25313 41515 25379 41518
rect 26200 41488 27000 41518
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 10593 41306 10659 41309
rect 11646 41306 11652 41308
rect 10593 41304 11652 41306
rect 10593 41248 10598 41304
rect 10654 41248 11652 41304
rect 10593 41246 11652 41248
rect 10593 41243 10659 41246
rect 11646 41244 11652 41246
rect 11716 41244 11722 41308
rect 2946 40832 3262 40833
rect 0 40762 800 40792
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 1301 40762 1367 40765
rect 0 40760 1367 40762
rect 0 40704 1306 40760
rect 1362 40704 1367 40760
rect 0 40702 1367 40704
rect 0 40672 800 40702
rect 1301 40699 1367 40702
rect 25313 40762 25379 40765
rect 26200 40762 27000 40792
rect 25313 40760 27000 40762
rect 25313 40704 25318 40760
rect 25374 40704 27000 40760
rect 25313 40702 27000 40704
rect 25313 40699 25379 40702
rect 26200 40672 27000 40702
rect 21449 40626 21515 40629
rect 22502 40626 22508 40628
rect 21449 40624 22508 40626
rect 21449 40568 21454 40624
rect 21510 40568 22508 40624
rect 21449 40566 22508 40568
rect 21449 40563 21515 40566
rect 22502 40564 22508 40566
rect 22572 40626 22578 40628
rect 23105 40626 23171 40629
rect 22572 40624 23171 40626
rect 22572 40568 23110 40624
rect 23166 40568 23171 40624
rect 22572 40566 23171 40568
rect 22572 40564 22578 40566
rect 23105 40563 23171 40566
rect 7649 40490 7715 40493
rect 9581 40490 9647 40493
rect 12433 40490 12499 40493
rect 15837 40492 15903 40493
rect 15837 40490 15884 40492
rect 7649 40488 12499 40490
rect 7649 40432 7654 40488
rect 7710 40432 9586 40488
rect 9642 40432 12438 40488
rect 12494 40432 12499 40488
rect 7649 40430 12499 40432
rect 15792 40488 15884 40490
rect 15792 40432 15842 40488
rect 15792 40430 15884 40432
rect 7649 40427 7715 40430
rect 9581 40427 9647 40430
rect 12433 40427 12499 40430
rect 15837 40428 15884 40430
rect 15948 40428 15954 40492
rect 21357 40490 21423 40493
rect 21633 40490 21699 40493
rect 21357 40488 21699 40490
rect 21357 40432 21362 40488
rect 21418 40432 21638 40488
rect 21694 40432 21699 40488
rect 21357 40430 21699 40432
rect 15837 40427 15903 40428
rect 21357 40427 21423 40430
rect 21633 40427 21699 40430
rect 21817 40490 21883 40493
rect 22921 40490 22987 40493
rect 21817 40488 22987 40490
rect 21817 40432 21822 40488
rect 21878 40432 22926 40488
rect 22982 40432 22987 40488
rect 21817 40430 22987 40432
rect 21817 40427 21883 40430
rect 22921 40427 22987 40430
rect 20529 40354 20595 40357
rect 24577 40354 24643 40357
rect 20529 40352 24643 40354
rect 20529 40296 20534 40352
rect 20590 40296 24582 40352
rect 24638 40296 24643 40352
rect 20529 40294 24643 40296
rect 20529 40291 20595 40294
rect 24577 40291 24643 40294
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 24761 39946 24827 39949
rect 26200 39946 27000 39976
rect 24761 39944 27000 39946
rect 24761 39888 24766 39944
rect 24822 39888 27000 39944
rect 24761 39886 27000 39888
rect 24761 39883 24827 39886
rect 26200 39856 27000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 17585 39402 17651 39405
rect 20437 39402 20503 39405
rect 17585 39400 20503 39402
rect 17585 39344 17590 39400
rect 17646 39344 20442 39400
rect 20498 39344 20503 39400
rect 17585 39342 20503 39344
rect 17585 39339 17651 39342
rect 20437 39339 20503 39342
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 24853 39130 24919 39133
rect 26200 39130 27000 39160
rect 24853 39128 27000 39130
rect 24853 39072 24858 39128
rect 24914 39072 27000 39128
rect 24853 39070 27000 39072
rect 24853 39067 24919 39070
rect 26200 39040 27000 39070
rect 9581 38858 9647 38861
rect 14365 38858 14431 38861
rect 9581 38856 14431 38858
rect 9581 38800 9586 38856
rect 9642 38800 14370 38856
rect 14426 38800 14431 38856
rect 9581 38798 14431 38800
rect 9581 38795 9647 38798
rect 14365 38795 14431 38798
rect 18413 38858 18479 38861
rect 18822 38858 18828 38860
rect 18413 38856 18828 38858
rect 18413 38800 18418 38856
rect 18474 38800 18828 38856
rect 18413 38798 18828 38800
rect 18413 38795 18479 38798
rect 18822 38796 18828 38798
rect 18892 38796 18898 38860
rect 16021 38724 16087 38725
rect 16021 38722 16068 38724
rect 15976 38720 16068 38722
rect 15976 38664 16026 38720
rect 15976 38662 16068 38664
rect 16021 38660 16068 38662
rect 16132 38660 16138 38724
rect 17350 38660 17356 38724
rect 17420 38722 17426 38724
rect 17585 38722 17651 38725
rect 17420 38720 17651 38722
rect 17420 38664 17590 38720
rect 17646 38664 17651 38720
rect 17420 38662 17651 38664
rect 17420 38660 17426 38662
rect 16021 38659 16087 38660
rect 17585 38659 17651 38662
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 17585 38586 17651 38589
rect 18873 38586 18939 38589
rect 17585 38584 18939 38586
rect 17585 38528 17590 38584
rect 17646 38528 18878 38584
rect 18934 38528 18939 38584
rect 17585 38526 18939 38528
rect 17585 38523 17651 38526
rect 18873 38523 18939 38526
rect 12617 38450 12683 38453
rect 13445 38450 13511 38453
rect 19425 38450 19491 38453
rect 12617 38448 19491 38450
rect 12617 38392 12622 38448
rect 12678 38392 13450 38448
rect 13506 38392 19430 38448
rect 19486 38392 19491 38448
rect 12617 38390 19491 38392
rect 12617 38387 12683 38390
rect 13445 38387 13511 38390
rect 19425 38387 19491 38390
rect 0 38314 800 38344
rect 1301 38314 1367 38317
rect 0 38312 1367 38314
rect 0 38256 1306 38312
rect 1362 38256 1367 38312
rect 0 38254 1367 38256
rect 0 38224 800 38254
rect 1301 38251 1367 38254
rect 7281 38314 7347 38317
rect 8201 38314 8267 38317
rect 11329 38314 11395 38317
rect 13813 38314 13879 38317
rect 7281 38312 13879 38314
rect 7281 38256 7286 38312
rect 7342 38256 8206 38312
rect 8262 38256 11334 38312
rect 11390 38256 13818 38312
rect 13874 38256 13879 38312
rect 7281 38254 13879 38256
rect 7281 38251 7347 38254
rect 8201 38251 8267 38254
rect 11329 38251 11395 38254
rect 13813 38251 13879 38254
rect 17217 38314 17283 38317
rect 25313 38314 25379 38317
rect 26200 38314 27000 38344
rect 17217 38312 18522 38314
rect 17217 38256 17222 38312
rect 17278 38256 18522 38312
rect 17217 38254 18522 38256
rect 17217 38251 17283 38254
rect 9806 38116 9812 38180
rect 9876 38178 9882 38180
rect 11421 38178 11487 38181
rect 16389 38178 16455 38181
rect 9876 38176 16455 38178
rect 9876 38120 11426 38176
rect 11482 38120 16394 38176
rect 16450 38120 16455 38176
rect 9876 38118 16455 38120
rect 9876 38116 9882 38118
rect 11421 38115 11487 38118
rect 16389 38115 16455 38118
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 18462 38042 18522 38254
rect 25313 38312 27000 38314
rect 25313 38256 25318 38312
rect 25374 38256 27000 38312
rect 25313 38254 27000 38256
rect 25313 38251 25379 38254
rect 26200 38224 27000 38254
rect 20294 38116 20300 38180
rect 20364 38178 20370 38180
rect 20437 38178 20503 38181
rect 20364 38176 20503 38178
rect 20364 38120 20442 38176
rect 20498 38120 20503 38176
rect 20364 38118 20503 38120
rect 20364 38116 20370 38118
rect 20437 38115 20503 38118
rect 19425 38042 19491 38045
rect 18462 38040 19491 38042
rect 18462 37984 19430 38040
rect 19486 37984 19491 38040
rect 18462 37982 19491 37984
rect 19425 37979 19491 37982
rect 12750 37844 12756 37908
rect 12820 37906 12826 37908
rect 20253 37906 20319 37909
rect 12820 37904 20319 37906
rect 12820 37848 20258 37904
rect 20314 37848 20319 37904
rect 12820 37846 20319 37848
rect 12820 37844 12826 37846
rect 20253 37843 20319 37846
rect 10542 37708 10548 37772
rect 10612 37770 10618 37772
rect 12433 37770 12499 37773
rect 18689 37770 18755 37773
rect 10612 37768 18755 37770
rect 10612 37712 12438 37768
rect 12494 37712 18694 37768
rect 18750 37712 18755 37768
rect 10612 37710 18755 37712
rect 10612 37708 10618 37710
rect 12433 37707 12499 37710
rect 18689 37707 18755 37710
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 25313 37498 25379 37501
rect 26200 37498 27000 37528
rect 25313 37496 27000 37498
rect 25313 37440 25318 37496
rect 25374 37440 27000 37496
rect 25313 37438 27000 37440
rect 25313 37435 25379 37438
rect 26200 37408 27000 37438
rect 18781 37362 18847 37365
rect 20437 37364 20503 37365
rect 19190 37362 19196 37364
rect 18781 37360 19196 37362
rect 18781 37304 18786 37360
rect 18842 37304 19196 37360
rect 18781 37302 19196 37304
rect 18781 37299 18847 37302
rect 19190 37300 19196 37302
rect 19260 37300 19266 37364
rect 20437 37362 20484 37364
rect 20392 37360 20484 37362
rect 20392 37304 20442 37360
rect 20392 37302 20484 37304
rect 20437 37300 20484 37302
rect 20548 37300 20554 37364
rect 20437 37299 20503 37300
rect 17769 37226 17835 37229
rect 19701 37226 19767 37229
rect 17769 37224 19767 37226
rect 17769 37168 17774 37224
rect 17830 37168 19706 37224
rect 19762 37168 19767 37224
rect 17769 37166 19767 37168
rect 17769 37163 17835 37166
rect 19701 37163 19767 37166
rect 22461 37226 22527 37229
rect 24025 37226 24091 37229
rect 22461 37224 24091 37226
rect 22461 37168 22466 37224
rect 22522 37168 24030 37224
rect 24086 37168 24091 37224
rect 22461 37166 24091 37168
rect 22461 37163 22527 37166
rect 24025 37163 24091 37166
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 9765 36818 9831 36821
rect 9949 36818 10015 36821
rect 16757 36818 16823 36821
rect 9765 36816 16823 36818
rect 9765 36760 9770 36816
rect 9826 36760 9954 36816
rect 10010 36760 16762 36816
rect 16818 36760 16823 36816
rect 9765 36758 16823 36760
rect 9765 36755 9831 36758
rect 9949 36755 10015 36758
rect 16757 36755 16823 36758
rect 12709 36682 12775 36685
rect 18965 36682 19031 36685
rect 12709 36680 19031 36682
rect 12709 36624 12714 36680
rect 12770 36624 18970 36680
rect 19026 36624 19031 36680
rect 12709 36622 19031 36624
rect 12709 36619 12775 36622
rect 18965 36619 19031 36622
rect 25313 36682 25379 36685
rect 26200 36682 27000 36712
rect 25313 36680 27000 36682
rect 25313 36624 25318 36680
rect 25374 36624 27000 36680
rect 25313 36622 27000 36624
rect 25313 36619 25379 36622
rect 26200 36592 27000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 11646 36212 11652 36276
rect 11716 36274 11722 36276
rect 12157 36274 12223 36277
rect 13813 36274 13879 36277
rect 11716 36272 13879 36274
rect 11716 36216 12162 36272
rect 12218 36216 13818 36272
rect 13874 36216 13879 36272
rect 11716 36214 13879 36216
rect 11716 36212 11722 36214
rect 12157 36211 12223 36214
rect 13813 36211 13879 36214
rect 19701 36274 19767 36277
rect 23606 36274 23612 36276
rect 19701 36272 23612 36274
rect 19701 36216 19706 36272
rect 19762 36216 23612 36272
rect 19701 36214 23612 36216
rect 19701 36211 19767 36214
rect 23606 36212 23612 36214
rect 23676 36212 23682 36276
rect 9254 35940 9260 36004
rect 9324 36002 9330 36004
rect 15745 36002 15811 36005
rect 9324 36000 15811 36002
rect 9324 35944 15750 36000
rect 15806 35944 15811 36000
rect 9324 35942 15811 35944
rect 9324 35940 9330 35942
rect 7946 35936 8262 35937
rect 0 35866 800 35896
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 1761 35866 1827 35869
rect 0 35864 1827 35866
rect 0 35808 1766 35864
rect 1822 35808 1827 35864
rect 0 35806 1827 35808
rect 0 35776 800 35806
rect 1761 35803 1827 35806
rect 7097 35730 7163 35733
rect 9446 35730 9506 35942
rect 15745 35939 15811 35942
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 12433 35866 12499 35869
rect 13445 35868 13511 35869
rect 12750 35866 12756 35868
rect 12433 35864 12756 35866
rect 12433 35808 12438 35864
rect 12494 35808 12756 35864
rect 12433 35806 12756 35808
rect 12433 35803 12499 35806
rect 12750 35804 12756 35806
rect 12820 35804 12826 35868
rect 13445 35866 13492 35868
rect 13400 35864 13492 35866
rect 13400 35808 13450 35864
rect 13400 35806 13492 35808
rect 13445 35804 13492 35806
rect 13556 35804 13562 35868
rect 25313 35866 25379 35869
rect 26200 35866 27000 35896
rect 25313 35864 27000 35866
rect 25313 35808 25318 35864
rect 25374 35808 27000 35864
rect 25313 35806 27000 35808
rect 13445 35803 13511 35804
rect 25313 35803 25379 35806
rect 26200 35776 27000 35806
rect 7097 35728 9506 35730
rect 7097 35672 7102 35728
rect 7158 35672 9506 35728
rect 7097 35670 9506 35672
rect 7097 35667 7163 35670
rect 13353 35458 13419 35461
rect 13353 35456 13554 35458
rect 13353 35400 13358 35456
rect 13414 35400 13554 35456
rect 13353 35398 13554 35400
rect 13353 35395 13419 35398
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 13353 35186 13419 35189
rect 13494 35186 13554 35398
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 13353 35184 13554 35186
rect 13353 35128 13358 35184
rect 13414 35128 13554 35184
rect 13353 35126 13554 35128
rect 13353 35123 13419 35126
rect 25313 35050 25379 35053
rect 26200 35050 27000 35080
rect 25313 35048 27000 35050
rect 25313 34992 25318 35048
rect 25374 34992 27000 35048
rect 25313 34990 27000 34992
rect 25313 34987 25379 34990
rect 26200 34960 27000 34990
rect 22461 34916 22527 34917
rect 22461 34914 22508 34916
rect 22416 34912 22508 34914
rect 22416 34856 22466 34912
rect 22416 34854 22508 34856
rect 22461 34852 22508 34854
rect 22572 34852 22578 34916
rect 22461 34851 22527 34852
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 25313 34234 25379 34237
rect 26200 34234 27000 34264
rect 25313 34232 27000 34234
rect 25313 34176 25318 34232
rect 25374 34176 27000 34232
rect 25313 34174 27000 34176
rect 25313 34171 25379 34174
rect 26200 34144 27000 34174
rect 8845 33962 8911 33965
rect 9397 33962 9463 33965
rect 8845 33960 9690 33962
rect 8845 33904 8850 33960
rect 8906 33904 9402 33960
rect 9458 33931 9690 33960
rect 9458 33926 9693 33931
rect 9458 33904 9632 33926
rect 8845 33902 9632 33904
rect 8845 33899 8911 33902
rect 9397 33899 9463 33902
rect 9627 33870 9632 33902
rect 9688 33870 9693 33926
rect 9627 33865 9693 33870
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 0 33418 800 33448
rect 1301 33418 1367 33421
rect 0 33416 1367 33418
rect 0 33360 1306 33416
rect 1362 33360 1367 33416
rect 0 33358 1367 33360
rect 0 33328 800 33358
rect 1301 33355 1367 33358
rect 24761 33418 24827 33421
rect 26200 33418 27000 33448
rect 24761 33416 27000 33418
rect 24761 33360 24766 33416
rect 24822 33360 27000 33416
rect 24761 33358 27000 33360
rect 24761 33355 24827 33358
rect 26200 33328 27000 33358
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 15653 32874 15719 32877
rect 21449 32874 21515 32877
rect 22737 32874 22803 32877
rect 15653 32872 22803 32874
rect 15653 32816 15658 32872
rect 15714 32816 21454 32872
rect 21510 32816 22742 32872
rect 22798 32816 22803 32872
rect 15653 32814 22803 32816
rect 15653 32811 15719 32814
rect 21449 32811 21515 32814
rect 22737 32811 22803 32814
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 21909 32602 21975 32605
rect 22686 32602 22692 32604
rect 21909 32600 22692 32602
rect 21909 32544 21914 32600
rect 21970 32544 22692 32600
rect 21909 32542 22692 32544
rect 21909 32539 21975 32542
rect 22686 32540 22692 32542
rect 22756 32540 22762 32604
rect 25313 32602 25379 32605
rect 26200 32602 27000 32632
rect 25313 32600 27000 32602
rect 25313 32544 25318 32600
rect 25374 32544 27000 32600
rect 25313 32542 27000 32544
rect 25313 32539 25379 32542
rect 26200 32512 27000 32542
rect 21081 32330 21147 32333
rect 22645 32330 22711 32333
rect 23197 32330 23263 32333
rect 21081 32328 23263 32330
rect 21081 32272 21086 32328
rect 21142 32272 22650 32328
rect 22706 32272 23202 32328
rect 23258 32272 23263 32328
rect 21081 32270 23263 32272
rect 21081 32267 21147 32270
rect 22645 32267 22711 32270
rect 23197 32267 23263 32270
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 25313 31786 25379 31789
rect 26200 31786 27000 31816
rect 25313 31784 27000 31786
rect 25313 31728 25318 31784
rect 25374 31728 27000 31784
rect 25313 31726 27000 31728
rect 25313 31723 25379 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 19977 31242 20043 31245
rect 20110 31242 20116 31244
rect 19977 31240 20116 31242
rect 19977 31184 19982 31240
rect 20038 31184 20116 31240
rect 19977 31182 20116 31184
rect 19977 31179 20043 31182
rect 20110 31180 20116 31182
rect 20180 31180 20186 31244
rect 2946 31040 3262 31041
rect 0 30970 800 31000
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 1301 30970 1367 30973
rect 12617 30972 12683 30973
rect 12566 30970 12572 30972
rect 0 30968 1367 30970
rect 0 30912 1306 30968
rect 1362 30912 1367 30968
rect 0 30910 1367 30912
rect 12526 30910 12572 30970
rect 12636 30968 12683 30972
rect 12678 30912 12683 30968
rect 0 30880 800 30910
rect 1301 30907 1367 30910
rect 12566 30908 12572 30910
rect 12636 30908 12683 30912
rect 20294 30908 20300 30972
rect 20364 30970 20370 30972
rect 20437 30970 20503 30973
rect 20364 30968 20503 30970
rect 20364 30912 20442 30968
rect 20498 30912 20503 30968
rect 20364 30910 20503 30912
rect 20364 30908 20370 30910
rect 12617 30907 12683 30908
rect 20437 30907 20503 30910
rect 25313 30970 25379 30973
rect 26200 30970 27000 31000
rect 25313 30968 27000 30970
rect 25313 30912 25318 30968
rect 25374 30912 27000 30968
rect 25313 30910 27000 30912
rect 25313 30907 25379 30910
rect 26200 30880 27000 30910
rect 13537 30564 13603 30565
rect 13486 30562 13492 30564
rect 13446 30502 13492 30562
rect 13556 30560 13603 30564
rect 13598 30504 13603 30560
rect 13486 30500 13492 30502
rect 13556 30500 13603 30504
rect 13537 30499 13603 30500
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 14038 30364 14044 30428
rect 14108 30426 14114 30428
rect 15193 30426 15259 30429
rect 16481 30426 16547 30429
rect 14108 30424 16547 30426
rect 14108 30368 15198 30424
rect 15254 30368 16486 30424
rect 16542 30368 16547 30424
rect 14108 30366 16547 30368
rect 14108 30364 14114 30366
rect 15193 30363 15259 30366
rect 16481 30363 16547 30366
rect 14365 30290 14431 30293
rect 14590 30290 14596 30292
rect 14365 30288 14596 30290
rect 14365 30232 14370 30288
rect 14426 30232 14596 30288
rect 14365 30230 14596 30232
rect 14365 30227 14431 30230
rect 14590 30228 14596 30230
rect 14660 30228 14666 30292
rect 19057 30290 19123 30293
rect 20662 30290 20668 30292
rect 19057 30288 20668 30290
rect 19057 30232 19062 30288
rect 19118 30232 20668 30288
rect 19057 30230 20668 30232
rect 19057 30227 19123 30230
rect 20662 30228 20668 30230
rect 20732 30228 20738 30292
rect 25313 30154 25379 30157
rect 26200 30154 27000 30184
rect 25313 30152 27000 30154
rect 25313 30096 25318 30152
rect 25374 30096 27000 30152
rect 25313 30094 27000 30096
rect 25313 30091 25379 30094
rect 26200 30064 27000 30094
rect 16113 30018 16179 30021
rect 16246 30018 16252 30020
rect 16113 30016 16252 30018
rect 16113 29960 16118 30016
rect 16174 29960 16252 30016
rect 16113 29958 16252 29960
rect 16113 29955 16179 29958
rect 16246 29956 16252 29958
rect 16316 29956 16322 30020
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 19517 29338 19583 29341
rect 20478 29338 20484 29340
rect 19517 29336 20484 29338
rect 19517 29280 19522 29336
rect 19578 29280 20484 29336
rect 19517 29278 20484 29280
rect 19517 29275 19583 29278
rect 20478 29276 20484 29278
rect 20548 29338 20554 29340
rect 22369 29338 22435 29341
rect 20548 29336 22435 29338
rect 20548 29280 22374 29336
rect 22430 29280 22435 29336
rect 20548 29278 22435 29280
rect 20548 29276 20554 29278
rect 22369 29275 22435 29278
rect 25497 29338 25563 29341
rect 26200 29338 27000 29368
rect 25497 29336 27000 29338
rect 25497 29280 25502 29336
rect 25558 29280 27000 29336
rect 25497 29278 27000 29280
rect 25497 29275 25563 29278
rect 26200 29248 27000 29278
rect 21449 29202 21515 29205
rect 16070 29200 21515 29202
rect 16070 29144 21454 29200
rect 21510 29144 21515 29200
rect 16070 29142 21515 29144
rect 15377 29066 15443 29069
rect 15745 29066 15811 29069
rect 16070 29066 16130 29142
rect 21449 29139 21515 29142
rect 15377 29064 16130 29066
rect 15377 29008 15382 29064
rect 15438 29008 15750 29064
rect 15806 29008 16130 29064
rect 15377 29006 16130 29008
rect 15377 29003 15443 29006
rect 15745 29003 15811 29006
rect 16246 29004 16252 29068
rect 16316 29066 16322 29068
rect 16389 29066 16455 29069
rect 16316 29064 16455 29066
rect 16316 29008 16394 29064
rect 16450 29008 16455 29064
rect 16316 29006 16455 29008
rect 16316 29004 16322 29006
rect 16389 29003 16455 29006
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 0 28522 800 28552
rect 1301 28522 1367 28525
rect 0 28520 1367 28522
rect 0 28464 1306 28520
rect 1362 28464 1367 28520
rect 0 28462 1367 28464
rect 0 28432 800 28462
rect 1301 28459 1367 28462
rect 18321 28522 18387 28525
rect 21582 28522 21588 28524
rect 18321 28520 21588 28522
rect 18321 28464 18326 28520
rect 18382 28464 21588 28520
rect 18321 28462 21588 28464
rect 18321 28459 18387 28462
rect 21582 28460 21588 28462
rect 21652 28460 21658 28524
rect 24853 28522 24919 28525
rect 26200 28522 27000 28552
rect 24853 28520 27000 28522
rect 24853 28464 24858 28520
rect 24914 28464 27000 28520
rect 24853 28462 27000 28464
rect 24853 28459 24919 28462
rect 26200 28432 27000 28462
rect 14222 28324 14228 28388
rect 14292 28386 14298 28388
rect 15193 28386 15259 28389
rect 14292 28384 15259 28386
rect 14292 28328 15198 28384
rect 15254 28328 15259 28384
rect 14292 28326 15259 28328
rect 14292 28324 14298 28326
rect 15193 28323 15259 28326
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 15929 28252 15995 28253
rect 15878 28188 15884 28252
rect 15948 28250 15995 28252
rect 15948 28248 16040 28250
rect 15990 28192 16040 28248
rect 15948 28190 16040 28192
rect 15948 28188 15995 28190
rect 19926 28188 19932 28252
rect 19996 28250 20002 28252
rect 20253 28250 20319 28253
rect 21950 28250 21956 28252
rect 19996 28248 21956 28250
rect 19996 28192 20258 28248
rect 20314 28192 21956 28248
rect 19996 28190 21956 28192
rect 19996 28188 20002 28190
rect 15929 28187 15995 28188
rect 20253 28187 20319 28190
rect 21950 28188 21956 28190
rect 22020 28188 22026 28252
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 24117 27706 24183 27709
rect 26200 27706 27000 27736
rect 24117 27704 27000 27706
rect 24117 27648 24122 27704
rect 24178 27648 27000 27704
rect 24117 27646 27000 27648
rect 24117 27643 24183 27646
rect 26200 27616 27000 27646
rect 17217 27436 17283 27437
rect 17166 27434 17172 27436
rect 17126 27374 17172 27434
rect 17236 27432 17283 27436
rect 17278 27376 17283 27432
rect 17166 27372 17172 27374
rect 17236 27372 17283 27376
rect 17217 27371 17283 27372
rect 14958 27236 14964 27300
rect 15028 27298 15034 27300
rect 15377 27298 15443 27301
rect 15028 27296 15443 27298
rect 15028 27240 15382 27296
rect 15438 27240 15443 27296
rect 15028 27238 15443 27240
rect 15028 27236 15034 27238
rect 15377 27235 15443 27238
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 25497 26890 25563 26893
rect 26200 26890 27000 26920
rect 25497 26888 27000 26890
rect 25497 26832 25502 26888
rect 25558 26832 27000 26888
rect 25497 26830 27000 26832
rect 25497 26827 25563 26830
rect 26200 26800 27000 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 15142 26284 15148 26348
rect 15212 26346 15218 26348
rect 17217 26346 17283 26349
rect 18321 26346 18387 26349
rect 15212 26344 18387 26346
rect 15212 26288 17222 26344
rect 17278 26288 18326 26344
rect 18382 26288 18387 26344
rect 15212 26286 18387 26288
rect 15212 26284 15218 26286
rect 17217 26283 17283 26286
rect 18321 26283 18387 26286
rect 7946 26144 8262 26145
rect 0 26074 800 26104
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 2773 26074 2839 26077
rect 0 26072 2839 26074
rect 0 26016 2778 26072
rect 2834 26016 2839 26072
rect 0 26014 2839 26016
rect 0 25984 800 26014
rect 2773 26011 2839 26014
rect 25313 26074 25379 26077
rect 26200 26074 27000 26104
rect 25313 26072 27000 26074
rect 25313 26016 25318 26072
rect 25374 26016 27000 26072
rect 25313 26014 27000 26016
rect 25313 26011 25379 26014
rect 26200 25984 27000 26014
rect 16113 25668 16179 25669
rect 16062 25604 16068 25668
rect 16132 25666 16179 25668
rect 16132 25664 16224 25666
rect 16174 25608 16224 25664
rect 16132 25606 16224 25608
rect 16132 25604 16179 25606
rect 16113 25603 16179 25604
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 25129 25258 25195 25261
rect 26200 25258 27000 25288
rect 25129 25256 27000 25258
rect 25129 25200 25134 25256
rect 25190 25200 27000 25256
rect 25129 25198 27000 25200
rect 25129 25195 25195 25198
rect 26200 25168 27000 25198
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 18638 24788 18644 24852
rect 18708 24850 18714 24852
rect 19241 24850 19307 24853
rect 18708 24848 19307 24850
rect 18708 24792 19246 24848
rect 19302 24792 19307 24848
rect 18708 24790 19307 24792
rect 18708 24788 18714 24790
rect 19241 24787 19307 24790
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 24945 24442 25011 24445
rect 26200 24442 27000 24472
rect 24945 24440 27000 24442
rect 24945 24384 24950 24440
rect 25006 24384 27000 24440
rect 24945 24382 27000 24384
rect 24945 24379 25011 24382
rect 26200 24352 27000 24382
rect 12157 24036 12223 24037
rect 12157 24032 12204 24036
rect 12268 24034 12274 24036
rect 12157 23976 12162 24032
rect 12157 23972 12204 23976
rect 12268 23974 12314 24034
rect 12268 23972 12274 23974
rect 12157 23971 12223 23972
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 17953 23762 18019 23765
rect 18638 23762 18644 23764
rect 17953 23760 18644 23762
rect 17953 23704 17958 23760
rect 18014 23704 18644 23760
rect 17953 23702 18644 23704
rect 17953 23699 18019 23702
rect 18638 23700 18644 23702
rect 18708 23700 18714 23764
rect 0 23626 800 23656
rect 1301 23626 1367 23629
rect 0 23624 1367 23626
rect 0 23568 1306 23624
rect 1362 23568 1367 23624
rect 0 23566 1367 23568
rect 0 23536 800 23566
rect 1301 23563 1367 23566
rect 23841 23626 23907 23629
rect 26200 23626 27000 23656
rect 23841 23624 27000 23626
rect 23841 23568 23846 23624
rect 23902 23568 27000 23624
rect 23841 23566 27000 23568
rect 23841 23563 23907 23566
rect 26200 23536 27000 23566
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 12157 22810 12223 22813
rect 15142 22810 15148 22812
rect 12157 22808 15148 22810
rect 12157 22752 12162 22808
rect 12218 22752 15148 22808
rect 12157 22750 15148 22752
rect 12157 22747 12223 22750
rect 15142 22748 15148 22750
rect 15212 22748 15218 22812
rect 23289 22810 23355 22813
rect 26200 22810 27000 22840
rect 23289 22808 27000 22810
rect 23289 22752 23294 22808
rect 23350 22752 27000 22808
rect 23289 22750 27000 22752
rect 23289 22747 23355 22750
rect 26200 22720 27000 22750
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 12382 22204 12388 22268
rect 12452 22266 12458 22268
rect 12750 22266 12756 22268
rect 12452 22206 12756 22266
rect 12452 22204 12458 22206
rect 12750 22204 12756 22206
rect 12820 22204 12826 22268
rect 24853 21994 24919 21997
rect 26200 21994 27000 22024
rect 24853 21992 27000 21994
rect 24853 21936 24858 21992
rect 24914 21936 27000 21992
rect 24853 21934 27000 21936
rect 24853 21931 24919 21934
rect 26200 21904 27000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 1301 21178 1367 21181
rect 19977 21180 20043 21181
rect 19926 21178 19932 21180
rect 0 21176 1367 21178
rect 0 21120 1306 21176
rect 1362 21120 1367 21176
rect 0 21118 1367 21120
rect 19886 21118 19932 21178
rect 19996 21176 20043 21180
rect 20038 21120 20043 21176
rect 0 21088 800 21118
rect 1301 21115 1367 21118
rect 19926 21116 19932 21118
rect 19996 21116 20043 21120
rect 19977 21115 20043 21116
rect 23381 21178 23447 21181
rect 26200 21178 27000 21208
rect 23381 21176 27000 21178
rect 23381 21120 23386 21176
rect 23442 21120 27000 21176
rect 23381 21118 27000 21120
rect 23381 21115 23447 21118
rect 26200 21088 27000 21118
rect 16021 20772 16087 20773
rect 16021 20768 16068 20772
rect 16132 20770 16138 20772
rect 16021 20712 16026 20768
rect 16021 20708 16068 20712
rect 16132 20710 16178 20770
rect 16132 20708 16138 20710
rect 16021 20707 16087 20708
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 17309 20636 17375 20637
rect 17309 20634 17356 20636
rect 17264 20632 17356 20634
rect 17264 20576 17314 20632
rect 17264 20574 17356 20576
rect 17309 20572 17356 20574
rect 17420 20572 17426 20636
rect 17309 20571 17375 20572
rect 24945 20362 25011 20365
rect 26200 20362 27000 20392
rect 24945 20360 27000 20362
rect 24945 20304 24950 20360
rect 25006 20304 27000 20360
rect 24945 20302 27000 20304
rect 24945 20299 25011 20302
rect 26200 20272 27000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 17769 19954 17835 19957
rect 18822 19954 18828 19956
rect 17769 19952 18828 19954
rect 17769 19896 17774 19952
rect 17830 19896 18828 19952
rect 17769 19894 18828 19896
rect 17769 19891 17835 19894
rect 18822 19892 18828 19894
rect 18892 19892 18898 19956
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 24761 19546 24827 19549
rect 26200 19546 27000 19576
rect 24761 19544 27000 19546
rect 24761 19488 24766 19544
rect 24822 19488 27000 19544
rect 24761 19486 27000 19488
rect 24761 19483 24827 19486
rect 26200 19456 27000 19486
rect 12157 19410 12223 19413
rect 14958 19410 14964 19412
rect 12157 19408 14964 19410
rect 12157 19352 12162 19408
rect 12218 19352 14964 19408
rect 12157 19350 14964 19352
rect 12157 19347 12223 19350
rect 14958 19348 14964 19350
rect 15028 19410 15034 19412
rect 17534 19410 17540 19412
rect 15028 19350 17540 19410
rect 15028 19348 15034 19350
rect 17534 19348 17540 19350
rect 17604 19348 17610 19412
rect 12341 19274 12407 19277
rect 12566 19274 12572 19276
rect 12341 19272 12572 19274
rect 12341 19216 12346 19272
rect 12402 19216 12572 19272
rect 12341 19214 12572 19216
rect 12341 19211 12407 19214
rect 12566 19212 12572 19214
rect 12636 19212 12642 19276
rect 12985 19274 13051 19277
rect 14549 19274 14615 19277
rect 12985 19272 14615 19274
rect 12985 19216 12990 19272
rect 13046 19216 14554 19272
rect 14610 19216 14615 19272
rect 12985 19214 14615 19216
rect 12985 19211 13051 19214
rect 14549 19211 14615 19214
rect 10869 19140 10935 19141
rect 10869 19138 10916 19140
rect 10824 19136 10916 19138
rect 10824 19080 10874 19136
rect 10824 19078 10916 19080
rect 10869 19076 10916 19078
rect 10980 19076 10986 19140
rect 10869 19075 10935 19076
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 0 18730 800 18760
rect 1301 18730 1367 18733
rect 0 18728 1367 18730
rect 0 18672 1306 18728
rect 1362 18672 1367 18728
rect 0 18670 1367 18672
rect 0 18640 800 18670
rect 1301 18667 1367 18670
rect 18321 18730 18387 18733
rect 20110 18730 20116 18732
rect 18321 18728 20116 18730
rect 18321 18672 18326 18728
rect 18382 18672 20116 18728
rect 18321 18670 20116 18672
rect 18321 18667 18387 18670
rect 20110 18668 20116 18670
rect 20180 18668 20186 18732
rect 24669 18730 24735 18733
rect 26200 18730 27000 18760
rect 24669 18728 27000 18730
rect 24669 18672 24674 18728
rect 24730 18672 27000 18728
rect 24669 18670 27000 18672
rect 24669 18667 24735 18670
rect 26200 18640 27000 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 11053 18186 11119 18189
rect 13813 18186 13879 18189
rect 11053 18184 13879 18186
rect 11053 18128 11058 18184
rect 11114 18128 13818 18184
rect 13874 18128 13879 18184
rect 11053 18126 13879 18128
rect 11053 18123 11119 18126
rect 13813 18123 13879 18126
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 12709 17916 12775 17917
rect 12709 17914 12756 17916
rect 12664 17912 12756 17914
rect 12664 17856 12714 17912
rect 12664 17854 12756 17856
rect 12709 17852 12756 17854
rect 12820 17852 12826 17916
rect 23381 17914 23447 17917
rect 26200 17914 27000 17944
rect 23381 17912 27000 17914
rect 23381 17856 23386 17912
rect 23442 17856 27000 17912
rect 23381 17854 27000 17856
rect 12709 17851 12775 17852
rect 23381 17851 23447 17854
rect 26200 17824 27000 17854
rect 16205 17644 16271 17645
rect 16205 17642 16252 17644
rect 16160 17640 16252 17642
rect 16160 17584 16210 17640
rect 16160 17582 16252 17584
rect 16205 17580 16252 17582
rect 16316 17580 16322 17644
rect 17861 17642 17927 17645
rect 19558 17642 19564 17644
rect 17861 17640 19564 17642
rect 17861 17584 17866 17640
rect 17922 17584 19564 17640
rect 17861 17582 19564 17584
rect 16205 17579 16271 17580
rect 17861 17579 17927 17582
rect 19558 17580 19564 17582
rect 19628 17580 19634 17644
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 24761 17098 24827 17101
rect 26200 17098 27000 17128
rect 24761 17096 27000 17098
rect 24761 17040 24766 17096
rect 24822 17040 27000 17096
rect 24761 17038 27000 17040
rect 24761 17035 24827 17038
rect 26200 17008 27000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 2497 16554 2563 16557
rect 4061 16554 4127 16557
rect 9489 16554 9555 16557
rect 2497 16552 9555 16554
rect 2497 16496 2502 16552
rect 2558 16496 4066 16552
rect 4122 16496 9494 16552
rect 9550 16496 9555 16552
rect 2497 16494 9555 16496
rect 2497 16491 2563 16494
rect 4061 16491 4127 16494
rect 9489 16491 9555 16494
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 16246 16220 16252 16284
rect 16316 16282 16322 16284
rect 16389 16282 16455 16285
rect 16316 16280 16455 16282
rect 16316 16224 16394 16280
rect 16450 16224 16455 16280
rect 16316 16222 16455 16224
rect 16316 16220 16322 16222
rect 16389 16219 16455 16222
rect 24669 16282 24735 16285
rect 26200 16282 27000 16312
rect 24669 16280 27000 16282
rect 24669 16224 24674 16280
rect 24730 16224 27000 16280
rect 24669 16222 27000 16224
rect 24669 16219 24735 16222
rect 26200 16192 27000 16222
rect 14181 16148 14247 16149
rect 14181 16146 14228 16148
rect 14136 16144 14228 16146
rect 14136 16088 14186 16144
rect 14136 16086 14228 16088
rect 14181 16084 14228 16086
rect 14292 16084 14298 16148
rect 14181 16083 14247 16084
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 24945 15466 25011 15469
rect 26200 15466 27000 15496
rect 24945 15464 27000 15466
rect 24945 15408 24950 15464
rect 25006 15408 27000 15464
rect 24945 15406 27000 15408
rect 24945 15403 25011 15406
rect 26200 15376 27000 15406
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 25129 14650 25195 14653
rect 26200 14650 27000 14680
rect 25129 14648 27000 14650
rect 25129 14592 25134 14648
rect 25190 14592 27000 14648
rect 25129 14590 27000 14592
rect 25129 14587 25195 14590
rect 26200 14560 27000 14590
rect 18597 14516 18663 14517
rect 18597 14514 18644 14516
rect 18552 14512 18644 14514
rect 18552 14456 18602 14512
rect 18552 14454 18644 14456
rect 18597 14452 18644 14454
rect 18708 14452 18714 14516
rect 18597 14451 18663 14452
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 0 13834 800 13864
rect 1301 13834 1367 13837
rect 0 13832 1367 13834
rect 0 13776 1306 13832
rect 1362 13776 1367 13832
rect 0 13774 1367 13776
rect 0 13744 800 13774
rect 1301 13771 1367 13774
rect 24761 13834 24827 13837
rect 26200 13834 27000 13864
rect 24761 13832 27000 13834
rect 24761 13776 24766 13832
rect 24822 13776 27000 13832
rect 24761 13774 27000 13776
rect 24761 13771 24827 13774
rect 26200 13744 27000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 25681 13018 25747 13021
rect 26200 13018 27000 13048
rect 25681 13016 27000 13018
rect 25681 12960 25686 13016
rect 25742 12960 27000 13016
rect 25681 12958 27000 12960
rect 25681 12955 25747 12958
rect 26200 12928 27000 12958
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 25129 12202 25195 12205
rect 26200 12202 27000 12232
rect 25129 12200 27000 12202
rect 25129 12144 25134 12200
rect 25190 12144 27000 12200
rect 25129 12142 27000 12144
rect 25129 12139 25195 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 17493 11932 17559 11933
rect 17493 11930 17540 11932
rect 17448 11928 17540 11930
rect 17448 11872 17498 11928
rect 17448 11870 17540 11872
rect 17493 11868 17540 11870
rect 17604 11868 17610 11932
rect 17493 11867 17559 11868
rect 3877 11658 3943 11661
rect 1902 11656 3943 11658
rect 1902 11600 3882 11656
rect 3938 11600 3943 11656
rect 1902 11598 3943 11600
rect 0 11386 800 11416
rect 1902 11386 1962 11598
rect 3877 11595 3943 11598
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 0 11326 1962 11386
rect 24761 11386 24827 11389
rect 26200 11386 27000 11416
rect 24761 11384 27000 11386
rect 24761 11328 24766 11384
rect 24822 11328 27000 11384
rect 24761 11326 27000 11328
rect 0 11296 800 11326
rect 24761 11323 24827 11326
rect 26200 11296 27000 11326
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 24669 10570 24735 10573
rect 26200 10570 27000 10600
rect 24669 10568 27000 10570
rect 24669 10512 24674 10568
rect 24730 10512 27000 10568
rect 24669 10510 27000 10512
rect 24669 10507 24735 10510
rect 26200 10480 27000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 24853 9754 24919 9757
rect 26200 9754 27000 9784
rect 24853 9752 27000 9754
rect 24853 9696 24858 9752
rect 24914 9696 27000 9752
rect 24853 9694 27000 9696
rect 24853 9691 24919 9694
rect 26200 9664 27000 9694
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 0 8938 800 8968
rect 3049 8938 3115 8941
rect 0 8936 3115 8938
rect 0 8880 3054 8936
rect 3110 8880 3115 8936
rect 0 8878 3115 8880
rect 0 8848 800 8878
rect 3049 8875 3115 8878
rect 25129 8938 25195 8941
rect 26200 8938 27000 8968
rect 25129 8936 27000 8938
rect 25129 8880 25134 8936
rect 25190 8880 27000 8936
rect 25129 8878 27000 8880
rect 25129 8875 25195 8878
rect 26200 8848 27000 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 25129 8122 25195 8125
rect 26200 8122 27000 8152
rect 25129 8120 27000 8122
rect 25129 8064 25134 8120
rect 25190 8064 27000 8120
rect 25129 8062 27000 8064
rect 25129 8059 25195 8062
rect 26200 8032 27000 8062
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 25129 7306 25195 7309
rect 26200 7306 27000 7336
rect 25129 7304 27000 7306
rect 25129 7248 25134 7304
rect 25190 7248 27000 7304
rect 25129 7246 27000 7248
rect 25129 7243 25195 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 3049 6490 3115 6493
rect 0 6488 3115 6490
rect 0 6432 3054 6488
rect 3110 6432 3115 6488
rect 0 6430 3115 6432
rect 0 6400 800 6430
rect 3049 6427 3115 6430
rect 24945 6490 25011 6493
rect 26200 6490 27000 6520
rect 24945 6488 27000 6490
rect 24945 6432 24950 6488
rect 25006 6432 27000 6488
rect 24945 6430 27000 6432
rect 24945 6427 25011 6430
rect 26200 6400 27000 6430
rect 5901 6354 5967 6357
rect 10910 6354 10916 6356
rect 5901 6352 10916 6354
rect 5901 6296 5906 6352
rect 5962 6296 10916 6352
rect 5901 6294 10916 6296
rect 5901 6291 5967 6294
rect 10910 6292 10916 6294
rect 10980 6292 10986 6356
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 7005 5674 7071 5677
rect 12198 5674 12204 5676
rect 7005 5672 12204 5674
rect 7005 5616 7010 5672
rect 7066 5616 12204 5672
rect 7005 5614 12204 5616
rect 7005 5611 7071 5614
rect 12198 5612 12204 5614
rect 12268 5612 12274 5676
rect 24761 5674 24827 5677
rect 26200 5674 27000 5704
rect 24761 5672 27000 5674
rect 24761 5616 24766 5672
rect 24822 5616 27000 5672
rect 24761 5614 27000 5616
rect 24761 5611 24827 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 23381 4858 23447 4861
rect 26200 4858 27000 4888
rect 23381 4856 27000 4858
rect 23381 4800 23386 4856
rect 23442 4800 27000 4856
rect 23381 4798 27000 4800
rect 23381 4795 23447 4798
rect 26200 4768 27000 4798
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 0 4042 800 4072
rect 3141 4042 3207 4045
rect 0 4040 3207 4042
rect 0 3984 3146 4040
rect 3202 3984 3207 4040
rect 0 3982 3207 3984
rect 0 3952 800 3982
rect 3141 3979 3207 3982
rect 20161 4042 20227 4045
rect 22093 4042 22159 4045
rect 20161 4040 22159 4042
rect 20161 3984 20166 4040
rect 20222 3984 22098 4040
rect 22154 3984 22159 4040
rect 20161 3982 22159 3984
rect 20161 3979 20227 3982
rect 22093 3979 22159 3982
rect 22369 4042 22435 4045
rect 26200 4042 27000 4072
rect 22369 4040 27000 4042
rect 22369 3984 22374 4040
rect 22430 3984 27000 4040
rect 22369 3982 27000 3984
rect 22369 3979 22435 3982
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 16297 3634 16363 3637
rect 23933 3634 23999 3637
rect 16297 3632 23999 3634
rect 16297 3576 16302 3632
rect 16358 3576 23938 3632
rect 23994 3576 23999 3632
rect 16297 3574 23999 3576
rect 16297 3571 16363 3574
rect 23933 3571 23999 3574
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 22553 3226 22619 3229
rect 26200 3226 27000 3256
rect 22553 3224 27000 3226
rect 22553 3168 22558 3224
rect 22614 3168 27000 3224
rect 22553 3166 27000 3168
rect 22553 3163 22619 3166
rect 26200 3136 27000 3166
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 22185 2410 22251 2413
rect 26200 2410 27000 2440
rect 22185 2408 27000 2410
rect 22185 2352 22190 2408
rect 22246 2352 27000 2408
rect 22185 2350 27000 2352
rect 22185 2347 22251 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1594 800 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 800 1534
rect 2865 1531 2931 1534
rect 25313 1594 25379 1597
rect 26200 1594 27000 1624
rect 25313 1592 27000 1594
rect 25313 1536 25318 1592
rect 25374 1536 27000 1592
rect 25313 1534 27000 1536
rect 25313 1531 25379 1534
rect 26200 1504 27000 1534
rect 24945 778 25011 781
rect 26200 778 27000 808
rect 24945 776 27000 778
rect 24945 720 24950 776
rect 25006 720 27000 776
rect 24945 718 27000 720
rect 24945 715 25011 718
rect 26200 688 27000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 17172 53892 17236 53956
rect 22692 53952 22756 53956
rect 22692 53896 22742 53952
rect 22742 53896 22756 53952
rect 22692 53892 22756 53896
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 14596 52940 14660 53004
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 14044 52592 14108 52596
rect 14044 52536 14058 52592
rect 14058 52536 14108 52592
rect 14044 52532 14108 52536
rect 16436 52592 16500 52596
rect 16436 52536 16450 52592
rect 16450 52536 16500 52592
rect 16436 52532 16500 52536
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 18828 47696 18892 47700
rect 18828 47640 18842 47696
rect 18842 47640 18892 47696
rect 18828 47636 18892 47640
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 19196 47092 19260 47156
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 21956 46608 22020 46612
rect 21956 46552 21970 46608
rect 21970 46552 22020 46608
rect 21956 46548 22020 46552
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 23612 45596 23676 45660
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 12388 44508 12452 44572
rect 9628 44236 9692 44300
rect 20668 44236 20732 44300
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 21588 43072 21652 43076
rect 21588 43016 21638 43072
rect 21638 43016 21652 43072
rect 21588 43012 21652 43016
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 9260 42468 9324 42532
rect 10548 42468 10612 42532
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 11652 41244 11716 41308
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 22508 40564 22572 40628
rect 15884 40488 15948 40492
rect 15884 40432 15898 40488
rect 15898 40432 15948 40488
rect 15884 40428 15948 40432
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 18828 38796 18892 38860
rect 16068 38720 16132 38724
rect 16068 38664 16082 38720
rect 16082 38664 16132 38720
rect 16068 38660 16132 38664
rect 17356 38660 17420 38724
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 9812 38116 9876 38180
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 20300 38116 20364 38180
rect 12756 37844 12820 37908
rect 10548 37708 10612 37772
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 19196 37300 19260 37364
rect 20484 37360 20548 37364
rect 20484 37304 20498 37360
rect 20498 37304 20548 37360
rect 20484 37300 20548 37304
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 11652 36212 11716 36276
rect 23612 36212 23676 36276
rect 9260 35940 9324 36004
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 12756 35804 12820 35868
rect 13492 35864 13556 35868
rect 13492 35808 13506 35864
rect 13506 35808 13556 35864
rect 13492 35804 13556 35808
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 22508 34912 22572 34916
rect 22508 34856 22522 34912
rect 22522 34856 22572 34912
rect 22508 34852 22572 34856
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 15148 34444 15212 34508
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 12020 33688 12084 33692
rect 12020 33632 12070 33688
rect 12070 33632 12084 33688
rect 12020 33628 12084 33632
rect 13860 33492 13924 33556
rect 17540 33356 17604 33420
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 22692 32540 22756 32604
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 20116 31180 20180 31244
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 12572 30968 12636 30972
rect 12572 30912 12622 30968
rect 12622 30912 12636 30968
rect 12572 30908 12636 30912
rect 20300 30908 20364 30972
rect 13492 30560 13556 30564
rect 13492 30504 13542 30560
rect 13542 30504 13556 30560
rect 13492 30500 13556 30504
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 14044 30364 14108 30428
rect 14596 30228 14660 30292
rect 20668 30228 20732 30292
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 20484 29276 20548 29340
rect 16252 29004 16316 29068
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 21588 28460 21652 28524
rect 14228 28324 14292 28388
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 15884 28248 15948 28252
rect 15884 28192 15934 28248
rect 15934 28192 15948 28248
rect 15884 28188 15948 28192
rect 19932 28188 19996 28252
rect 21956 28188 22020 28252
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 17172 27432 17236 27436
rect 17172 27376 17222 27432
rect 17222 27376 17236 27432
rect 17172 27372 17236 27376
rect 14964 27236 15028 27300
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 15148 26284 15212 26348
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 16068 25664 16132 25668
rect 16068 25608 16118 25664
rect 16118 25608 16132 25664
rect 16068 25604 16132 25608
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 18644 24788 18708 24852
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 12204 24032 12268 24036
rect 12204 23976 12218 24032
rect 12218 23976 12268 24032
rect 12204 23972 12268 23976
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 18644 23700 18708 23764
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 17724 23292 17788 23356
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 15148 22748 15212 22812
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 12388 22204 12452 22268
rect 12756 22204 12820 22268
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 19932 21176 19996 21180
rect 19932 21120 19982 21176
rect 19982 21120 19996 21176
rect 19932 21116 19996 21120
rect 16068 20768 16132 20772
rect 16068 20712 16082 20768
rect 16082 20712 16132 20768
rect 16068 20708 16132 20712
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 17356 20632 17420 20636
rect 17356 20576 17370 20632
rect 17370 20576 17420 20632
rect 17356 20572 17420 20576
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 18828 19892 18892 19956
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 14964 19348 15028 19412
rect 17540 19348 17604 19412
rect 12572 19212 12636 19276
rect 10916 19136 10980 19140
rect 10916 19080 10930 19136
rect 10930 19080 10980 19136
rect 10916 19076 10980 19080
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 20116 18668 20180 18732
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 12756 17912 12820 17916
rect 12756 17856 12770 17912
rect 12770 17856 12820 17912
rect 12756 17852 12820 17856
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 16252 16220 16316 16284
rect 14228 16144 14292 16148
rect 14228 16088 14242 16144
rect 14242 16088 14292 16144
rect 14228 16084 14292 16088
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 18644 14512 18708 14516
rect 18644 14456 18658 14512
rect 18658 14456 18708 14512
rect 18644 14452 18708 14456
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 19564 13500 19628 13564
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 17540 11928 17604 11932
rect 17540 11872 17554 11928
rect 17554 11872 17604 11928
rect 17540 11868 17604 11872
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 10916 6292 10980 6356
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 12204 5612 12268 5676
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 15700 2680 15764 2684
rect 15700 2624 15714 2680
rect 15714 2624 15764 2680
rect 15700 2620 15764 2624
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 12944 53888 13264 54448
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17171 53956 17237 53957
rect 17171 53892 17172 53956
rect 17236 53892 17237 53956
rect 17171 53891 17237 53892
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 14595 53004 14661 53005
rect 14595 52940 14596 53004
rect 14660 52940 14661 53004
rect 14595 52939 14661 52940
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 14043 52596 14109 52597
rect 14043 52532 14044 52596
rect 14108 52532 14109 52596
rect 14043 52531 14109 52532
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12387 44572 12453 44573
rect 12387 44508 12388 44572
rect 12452 44508 12453 44572
rect 12387 44507 12453 44508
rect 9627 44300 9693 44301
rect 9627 44236 9628 44300
rect 9692 44236 9693 44300
rect 9627 44235 9693 44236
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 9259 42532 9325 42533
rect 9259 42468 9260 42532
rect 9324 42468 9325 42532
rect 9259 42467 9325 42468
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 9262 36005 9322 42467
rect 9630 38670 9690 44235
rect 10547 42532 10613 42533
rect 10547 42468 10548 42532
rect 10612 42468 10613 42532
rect 10547 42467 10613 42468
rect 9630 38610 9874 38670
rect 9814 38181 9874 38610
rect 9811 38180 9877 38181
rect 9811 38116 9812 38180
rect 9876 38116 9877 38180
rect 9811 38115 9877 38116
rect 10550 37773 10610 42467
rect 12390 41430 12450 44507
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12390 41370 12818 41430
rect 11651 41308 11717 41309
rect 11651 41244 11652 41308
rect 11716 41244 11717 41308
rect 11651 41243 11717 41244
rect 10547 37772 10613 37773
rect 10547 37708 10548 37772
rect 10612 37708 10613 37772
rect 10547 37707 10613 37708
rect 11654 36277 11714 41243
rect 12758 37909 12818 41370
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12755 37908 12821 37909
rect 12755 37844 12756 37908
rect 12820 37844 12821 37908
rect 12755 37843 12821 37844
rect 11651 36276 11717 36277
rect 11651 36212 11652 36276
rect 11716 36212 11717 36276
rect 11651 36211 11717 36212
rect 9259 36004 9325 36005
rect 9259 35940 9260 36004
rect 9324 35940 9325 36004
rect 9259 35939 9325 35940
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 12758 35869 12818 37843
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12755 35868 12821 35869
rect 12755 35804 12756 35868
rect 12820 35804 12821 35868
rect 12755 35803 12821 35804
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 12571 30972 12637 30973
rect 12571 30908 12572 30972
rect 12636 30908 12637 30972
rect 12571 30907 12637 30908
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 13862 30701 13922 33491
rect 14414 31925 14474 52531
rect 14595 40764 14661 40765
rect 14595 40700 14596 40764
rect 14660 40700 14661 40764
rect 14595 40699 14661 40700
rect 14411 31924 14477 31925
rect 14411 31860 14412 31924
rect 14476 31860 14477 31924
rect 14411 31859 14477 31860
rect 13859 30700 13925 30701
rect 13859 30636 13860 30700
rect 13924 30636 13925 30700
rect 13859 30635 13925 30636
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12755 29476 12821 29477
rect 12755 29412 12756 29476
rect 12820 29412 12821 29476
rect 12755 29411 12821 29412
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 12203 24036 12269 24037
rect 12203 23972 12204 24036
rect 12268 23972 12269 24036
rect 12203 23971 12269 23972
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 10915 19140 10981 19141
rect 10915 19076 10916 19140
rect 10980 19076 10981 19140
rect 10915 19075 10981 19076
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 10918 6357 10978 19075
rect 10915 6356 10981 6357
rect 10915 6292 10916 6356
rect 10980 6292 10981 6356
rect 10915 6291 10981 6292
rect 12206 5677 12266 23971
rect 12387 22268 12453 22269
rect 12387 22204 12388 22268
rect 12452 22204 12453 22268
rect 12387 22203 12453 22204
rect 12390 21450 12450 22203
rect 12574 22110 12634 30907
rect 12758 22269 12818 35803
rect 12944 35392 13264 36416
rect 13491 35868 13557 35869
rect 13491 35804 13492 35868
rect 13556 35804 13557 35868
rect 13491 35803 13557 35804
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 13494 30565 13554 35803
rect 13491 30564 13557 30565
rect 13491 30500 13492 30564
rect 13556 30500 13557 30564
rect 13491 30499 13557 30500
rect 14046 30429 14106 52531
rect 14043 30428 14109 30429
rect 14043 30364 14044 30428
rect 14108 30364 14109 30428
rect 14043 30363 14109 30364
rect 14598 30293 14658 52939
rect 16435 52596 16501 52597
rect 16435 52532 16436 52596
rect 16500 52532 16501 52596
rect 16435 52531 16501 52532
rect 15883 40492 15949 40493
rect 15883 40428 15884 40492
rect 15948 40428 15949 40492
rect 15883 40427 15949 40428
rect 14595 30292 14661 30293
rect 14595 30228 14596 30292
rect 14660 30228 14661 30292
rect 14595 30227 14661 30228
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 14227 28388 14293 28389
rect 14227 28324 14228 28388
rect 14292 28324 14293 28388
rect 14227 28323 14293 28324
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 13491 23492 13557 23493
rect 13491 23428 13492 23492
rect 13556 23428 13557 23492
rect 13491 23427 13557 23428
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12755 22676 12821 22677
rect 12755 22612 12756 22676
rect 12820 22612 12821 22676
rect 12755 22611 12821 22612
rect 12944 22336 13264 23360
rect 13494 22541 13554 23427
rect 13491 22540 13557 22541
rect 13491 22476 13492 22540
rect 13556 22476 13557 22540
rect 13491 22475 13557 22476
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12755 22268 12821 22269
rect 12755 22204 12756 22268
rect 12820 22204 12821 22268
rect 12755 22203 12821 22204
rect 12574 22050 12818 22110
rect 12390 21390 12634 21450
rect 12574 19277 12634 21390
rect 12571 19276 12637 19277
rect 12571 19212 12572 19276
rect 12636 19212 12637 19276
rect 12571 19211 12637 19212
rect 12758 17917 12818 22050
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12755 17916 12821 17917
rect 12755 17852 12756 17916
rect 12820 17852 12821 17916
rect 12755 17851 12821 17852
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 14230 16149 14290 28323
rect 15886 28253 15946 40427
rect 16067 38724 16133 38725
rect 16067 38660 16068 38724
rect 16132 38660 16133 38724
rect 16067 38659 16133 38660
rect 15883 28252 15949 28253
rect 15883 28188 15884 28252
rect 15948 28188 15949 28252
rect 15883 28187 15949 28188
rect 14963 27300 15029 27301
rect 14963 27236 14964 27300
rect 15028 27236 15029 27300
rect 14963 27235 15029 27236
rect 14966 19413 15026 27235
rect 15147 26348 15213 26349
rect 15147 26284 15148 26348
rect 15212 26284 15213 26348
rect 15147 26283 15213 26284
rect 15150 22813 15210 26283
rect 15147 22812 15213 22813
rect 15147 22748 15148 22812
rect 15212 22748 15213 22812
rect 15147 22747 15213 22748
rect 16070 20773 16130 38659
rect 16438 31770 16498 52531
rect 16254 31710 16498 31770
rect 16254 29069 16314 31710
rect 16251 29068 16317 29069
rect 16251 29004 16252 29068
rect 16316 29004 16317 29068
rect 16251 29003 16317 29004
rect 16067 20772 16133 20773
rect 16067 20708 16068 20772
rect 16132 20708 16133 20772
rect 16067 20707 16133 20708
rect 14963 19412 15029 19413
rect 14963 19348 14964 19412
rect 15028 19348 15029 19412
rect 14963 19347 15029 19348
rect 16254 16285 16314 29003
rect 17174 27437 17234 53891
rect 17944 53344 18264 54368
rect 22691 53956 22757 53957
rect 22691 53892 22692 53956
rect 22756 53892 22757 53956
rect 22691 53891 22757 53892
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 18827 47700 18893 47701
rect 18827 47636 18828 47700
rect 18892 47636 18893 47700
rect 18827 47635 18893 47636
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 19379 44300 19445 44301
rect 19379 44236 19380 44300
rect 19444 44236 19445 44300
rect 19379 44235 19445 44236
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17355 38724 17421 38725
rect 17355 38660 17356 38724
rect 17420 38660 17421 38724
rect 17355 38659 17421 38660
rect 17171 27436 17237 27437
rect 17171 27372 17172 27436
rect 17236 27372 17237 27436
rect 17171 27371 17237 27372
rect 17358 20637 17418 38659
rect 17944 38112 18264 39136
rect 18830 38861 18890 47635
rect 19195 47156 19261 47157
rect 19195 47092 19196 47156
rect 19260 47092 19261 47156
rect 19195 47091 19261 47092
rect 18827 38860 18893 38861
rect 18827 38796 18828 38860
rect 18892 38796 18893 38860
rect 18827 38795 18893 38796
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 18643 24852 18709 24853
rect 18643 24788 18644 24852
rect 18708 24788 18709 24852
rect 18643 24787 18709 24788
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 18646 23765 18706 24787
rect 18643 23764 18709 23765
rect 18643 23700 18644 23764
rect 18708 23700 18709 23764
rect 18643 23699 18709 23700
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17723 22268 17789 22269
rect 17723 22204 17724 22268
rect 17788 22204 17789 22268
rect 17723 22203 17789 22204
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17539 19412 17605 19413
rect 17539 19348 17540 19412
rect 17604 19348 17605 19412
rect 17539 19347 17605 19348
rect 16251 16284 16317 16285
rect 16251 16220 16252 16284
rect 16316 16220 16317 16284
rect 16251 16219 16317 16220
rect 14227 16148 14293 16149
rect 14227 16084 14228 16148
rect 14292 16084 14293 16148
rect 14227 16083 14293 16084
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 17542 11933 17602 19347
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 18646 14517 18706 23699
rect 18830 19957 18890 38795
rect 19198 37365 19258 47091
rect 21955 46612 22021 46613
rect 21955 46548 21956 46612
rect 22020 46548 22021 46612
rect 21955 46547 22021 46548
rect 20667 44300 20733 44301
rect 20667 44236 20668 44300
rect 20732 44236 20733 44300
rect 20667 44235 20733 44236
rect 20299 38180 20365 38181
rect 20299 38116 20300 38180
rect 20364 38116 20365 38180
rect 20299 38115 20365 38116
rect 19195 37364 19261 37365
rect 19195 37300 19196 37364
rect 19260 37300 19261 37364
rect 19195 37299 19261 37300
rect 20115 31244 20181 31245
rect 20115 31180 20116 31244
rect 20180 31180 20181 31244
rect 20115 31179 20181 31180
rect 19931 28252 19997 28253
rect 19931 28188 19932 28252
rect 19996 28188 19997 28252
rect 19931 28187 19997 28188
rect 19934 21181 19994 28187
rect 19931 21180 19997 21181
rect 19931 21116 19932 21180
rect 19996 21116 19997 21180
rect 19931 21115 19997 21116
rect 18827 19956 18893 19957
rect 18827 19892 18828 19956
rect 18892 19892 18893 19956
rect 18827 19891 18893 19892
rect 20118 18733 20178 31179
rect 20302 30973 20362 38115
rect 20483 37364 20549 37365
rect 20483 37300 20484 37364
rect 20548 37300 20549 37364
rect 20483 37299 20549 37300
rect 20299 30972 20365 30973
rect 20299 30908 20300 30972
rect 20364 30908 20365 30972
rect 20299 30907 20365 30908
rect 20486 29341 20546 37299
rect 20670 30293 20730 44235
rect 21587 43076 21653 43077
rect 21587 43012 21588 43076
rect 21652 43012 21653 43076
rect 21587 43011 21653 43012
rect 20667 30292 20733 30293
rect 20667 30228 20668 30292
rect 20732 30228 20733 30292
rect 20667 30227 20733 30228
rect 20483 29340 20549 29341
rect 20483 29276 20484 29340
rect 20548 29276 20549 29340
rect 20483 29275 20549 29276
rect 21590 28525 21650 43011
rect 21587 28524 21653 28525
rect 21587 28460 21588 28524
rect 21652 28460 21653 28524
rect 21587 28459 21653 28460
rect 21958 28253 22018 46547
rect 22507 40628 22573 40629
rect 22507 40564 22508 40628
rect 22572 40564 22573 40628
rect 22507 40563 22573 40564
rect 22510 34917 22570 40563
rect 22507 34916 22573 34917
rect 22507 34852 22508 34916
rect 22572 34852 22573 34916
rect 22507 34851 22573 34852
rect 22694 32605 22754 53891
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 23611 45660 23677 45661
rect 23611 45596 23612 45660
rect 23676 45596 23677 45660
rect 23611 45595 23677 45596
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 23614 36277 23674 45595
rect 23611 36276 23677 36277
rect 23611 36212 23612 36276
rect 23676 36212 23677 36276
rect 23611 36211 23677 36212
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22507 35188 22573 35189
rect 22507 35124 22508 35188
rect 22572 35124 22573 35188
rect 22507 35123 22573 35124
rect 22323 31788 22389 31789
rect 22323 31724 22324 31788
rect 22388 31724 22389 31788
rect 22323 31723 22389 31724
rect 22510 29749 22570 35123
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22691 32604 22757 32605
rect 22691 32540 22692 32604
rect 22756 32540 22757 32604
rect 22691 32539 22757 32540
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22507 29748 22573 29749
rect 22507 29684 22508 29748
rect 22572 29684 22573 29748
rect 22507 29683 22573 29684
rect 22944 28864 23264 29888
rect 23427 29476 23493 29477
rect 23427 29412 23428 29476
rect 23492 29412 23493 29476
rect 23427 29411 23493 29412
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 21955 28252 22021 28253
rect 21955 28188 21956 28252
rect 22020 28188 22021 28252
rect 21955 28187 22021 28188
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 23430 26213 23490 29411
rect 23427 26212 23493 26213
rect 23427 26148 23428 26212
rect 23492 26148 23493 26212
rect 23427 26147 23493 26148
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 20851 24580 20917 24581
rect 20851 24516 20852 24580
rect 20916 24516 20917 24580
rect 20851 24515 20917 24516
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 20115 18732 20181 18733
rect 20115 18668 20116 18732
rect 20180 18668 20181 18732
rect 20115 18667 20181 18668
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 18643 14516 18709 14517
rect 18643 14452 18644 14516
rect 18708 14452 18709 14516
rect 18643 14451 18709 14452
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 19566 13565 19626 17579
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 19563 13564 19629 13565
rect 19563 13500 19564 13564
rect 19628 13500 19629 13564
rect 19563 13499 19629 13500
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17539 11932 17605 11933
rect 17539 11868 17540 11932
rect 17604 11868 17605 11932
rect 17539 11867 17605 11868
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12203 5676 12269 5677
rect 12203 5612 12204 5676
rect 12268 5612 12269 5676
rect 12203 5611 12269 5612
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 16803 3500 16869 3501
rect 16803 3436 16804 3500
rect 16868 3436 16869 3500
rect 16803 3435 16869 3436
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 15699 2684 15765 2685
rect 15699 2620 15700 2684
rect 15764 2620 15765 2684
rect 15699 2619 15765 2620
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _109_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _111_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23184 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _112_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23736 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1676037725
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1676037725
transform 1 0 24656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 16008 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 23184 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 20700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 21160 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 21160 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1676037725
transform 1 0 24656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform 1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1676037725
transform 1 0 21896 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 23184 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1676037725
transform 1 0 23736 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform 1 0 24564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1676037725
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 25024 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform -1 0 23000 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22172 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 14076 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 13616 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 15824 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 15272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 17112 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 18400 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 19504 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 20608 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 19596 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 20332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 18676 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 20792 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1676037725
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform 1 0 21068 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1676037725
transform 1 0 20240 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1676037725
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1676037725
transform 1 0 3128 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform 1 0 4876 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform 1 0 4140 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform 1 0 12696 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 4692 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1676037725
transform 1 0 4968 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1676037725
transform 1 0 6532 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1676037725
transform 1 0 6808 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1676037725
transform 1 0 6624 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1676037725
transform 1 0 6532 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1676037725
transform 1 0 7268 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _179_
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1676037725
transform 1 0 7636 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1676037725
transform 1 0 7912 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1676037725
transform 1 0 8832 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1676037725
transform 1 0 6808 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1676037725
transform 1 0 9108 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1676037725
transform 1 0 8372 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1676037725
transform 1 0 10396 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1676037725
transform 1 0 9200 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1676037725
transform 1 0 11408 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1676037725
transform 1 0 10856 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1676037725
transform 1 0 11408 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1676037725
transform 1 0 9016 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1676037725
transform 1 0 9292 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1676037725
transform 1 0 12236 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1676037725
transform 1 0 10212 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1676037725
transform 1 0 11684 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1676037725
transform 1 0 12604 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1676037725
transform 1 0 12328 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1676037725
transform 1 0 2392 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1676037725
transform 1 0 2024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1676037725
transform 1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1676037725
transform 1 0 2024 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1676037725
transform 1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1676037725
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1676037725
transform 1 0 2024 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11960 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 11224 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1676037725
transform 1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1676037725
transform 1 0 17388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1676037725
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1676037725
transform 1 0 16100 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1676037725
transform 1 0 17204 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1676037725
transform 1 0 17112 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1676037725
transform 1 0 18952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1676037725
transform 1 0 18124 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1676037725
transform 1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1676037725
transform 1 0 20700 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1676037725
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A
timestamp 1676037725
transform 1 0 3680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A
timestamp 1676037725
transform 1 0 5428 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1676037725
transform 1 0 3772 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1676037725
transform 1 0 5244 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1676037725
transform 1 0 5520 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1676037725
transform 1 0 7084 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1676037725
transform 1 0 7176 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1676037725
transform 1 0 6348 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1676037725
transform 1 0 8464 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1676037725
transform 1 0 9384 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1676037725
transform 1 0 9660 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1676037725
transform 1 0 10212 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1676037725
transform 1 0 11960 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1676037725
transform 1 0 11040 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1676037725
transform 1 0 12052 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 9384 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11868 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 7728 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11960 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 10028 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12972 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 7820 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 13524 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 13800 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 12420 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 12604 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__S
timestamp 1676037725
transform 1 0 11040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 12144 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16008 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 14628 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 12420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 11040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16192 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 12604 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 12972 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 10028 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 8556 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 13156 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 15272 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 13616 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 11776 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 12052 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 10028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 10396 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 3956 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 5704 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 2576 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6624 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 4324 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 5980 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 16652 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 12328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform 1 0 9200 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 17112 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 21528 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform 1 0 17480 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform 1 0 20332 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 10304 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform 1 0 10672 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 13156 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 21068 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform 1 0 18492 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1676037725
transform 1 0 2024 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform 1 0 2024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform 1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform 1 0 25208 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform 1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform 1 0 24748 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform 1 0 24472 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform 1 0 24748 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform 1 0 24564 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform 1 0 24564 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform 1 0 25392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform 1 0 25208 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform 1 0 25392 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform 1 0 24748 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 24748 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 24748 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 25392 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform 1 0 23552 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform 1 0 25392 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform 1 0 25208 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform 1 0 24748 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform 1 0 24748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform 1 0 24748 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform 1 0 24748 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform 1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform 1 0 4600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform 1 0 7176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform 1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform 1 0 2208 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform 1 0 9016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 10580 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform 1 0 9200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform 1 0 3036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform 1 0 5796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform 1 0 16284 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform 1 0 18860 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform 1 0 17204 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform 1 0 18860 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform 1 0 18676 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform 1 0 19688 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform 1 0 19320 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform 1 0 19504 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform 1 0 21436 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform 1 0 20700 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform 1 0 13156 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform 1 0 20792 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform 1 0 21160 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform 1 0 20976 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform 1 0 23276 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform 1 0 22264 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1676037725
transform 1 0 22540 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1676037725
transform 1 0 24380 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1676037725
transform 1 0 14812 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1676037725
transform 1 0 14904 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1676037725
transform 1 0 14444 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1676037725
transform 1 0 16100 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1676037725
transform 1 0 16100 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1676037725
transform 1 0 16376 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1676037725
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1676037725
transform 1 0 2024 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1676037725
transform 1 0 2024 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1676037725
transform 1 0 2024 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1676037725
transform 1 0 2024 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1676037725
transform 1 0 2116 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1676037725
transform 1 0 25392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1676037725
transform 1 0 24656 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1676037725
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1676037725
transform 1 0 24656 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1676037725
transform 1 0 24656 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1676037725
transform 1 0 25208 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1676037725
transform 1 0 24472 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1676037725
transform 1 0 24564 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1676037725
transform 1 0 2116 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1676037725
transform 1 0 5060 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16100 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18492 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21896 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 17940 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20884 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25116 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25116 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18216 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 15824 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17112 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16100 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 14904 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17940 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20424 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20792 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25392 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24748 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25392 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23920 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25208 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24656 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 23736 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21344 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20332 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20424 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 17664 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 17112 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 15640 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14904 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12420 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11592 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13248 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14352 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14720 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13156 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11776 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10304 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9752 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8556 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8372 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8464 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10304 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8372 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13524 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23736 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22908 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20240 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 8832 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 12236 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15180 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 14168 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14260 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12972 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10580 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8648 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 7268 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8648 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 7544 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8464 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 7084 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10304 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10856 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10120 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8096 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 5980 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6900 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 7912 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9292 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12788 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 17848 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 12328 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 11592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18860 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20056 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 20424 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 16836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19688 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23000 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 19872 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17480 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18676 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21436 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 18124 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 16468 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16744 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17940 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 13064 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18584 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18768 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 17204 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20516 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20700 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 19688 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15732 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17296 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 18032 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18768 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 13064 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_45.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20424 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 23276 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 22816 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 22632 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21896 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 22264 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 22264 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 21252 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 21436 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21620 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 23920 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24104 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 19412 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 23184 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23000 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 20608 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 21252 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21620 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 22080 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21896 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 18584 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 20608 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20700 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 20976 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 20792 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 15732 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19320 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 20240 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 19044 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19044 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 17848 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 13800 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17664 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 17204 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 12328 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15640 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 14168 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 11592 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13616 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 10028 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16100 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 12696 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17848 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 11040 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16100 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15088 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 8832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 8556 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12420 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12236 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 7268 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15272 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12880 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12512 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 6900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16008 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17204 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17296 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18308 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 23276 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 23092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21068 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18308 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 18124 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 14536 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 15548 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 8832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 9016 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 12144 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 12328 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 10580 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 10764 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 8464 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 8464 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 12420 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 7084 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12512 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 7268 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 7452 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15732 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14352 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 9108 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13984 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 12512 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 4600 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 7452 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_44.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_52.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4048 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9752 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 5704 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9936 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 8004 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11040 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6624 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 5336 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9752 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 5796 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11684 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 8740 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__256 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 11316 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9936 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 8280 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 7084 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15640 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15272 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 14260 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 11408 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 10120 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__257
timestamp 1676037725
transform 1 0 13248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10488 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14444 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14352 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12972 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10396 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12328 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11776 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 8740 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__258
timestamp 1676037725
transform 1 0 11868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 8924 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 6256 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4232 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13524 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__259
timestamp 1676037725
transform 1 0 9844 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9476 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 6808 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4048 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3680 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 4232 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 3036 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 2944 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 2760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 4232 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 3956 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 4508 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 3404 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3956 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 3680 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 9016 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9844 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8464 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 10488 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 8004 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 9936 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 17480 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 17848 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 20516 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 9108 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 10212 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 9292 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 11960 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 19412 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18
timestamp 1676037725
transform 1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35
timestamp 1676037725
transform 1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1676037725
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1676037725
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1676037725
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1676037725
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1676037725
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1676037725
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp 1676037725
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_264
timestamp 1676037725
transform 1 0 25392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_5
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1676037725
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_33
timestamp 1676037725
transform 1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_37
timestamp 1676037725
transform 1 0 4508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_40
timestamp 1676037725
transform 1 0 4784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_59
timestamp 1676037725
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_66
timestamp 1676037725
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1676037725
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1676037725
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1676037725
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1676037725
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1676037725
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1676037725
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_207 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1676037725
transform 1 0 23460 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_10
timestamp 1676037725
transform 1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_16
timestamp 1676037725
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_25
timestamp 1676037725
transform 1 0 3404 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_37
timestamp 1676037725
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_47
timestamp 1676037725
transform 1 0 5428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_51
timestamp 1676037725
transform 1 0 5796 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1676037725
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_63
timestamp 1676037725
transform 1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_68
timestamp 1676037725
transform 1 0 7360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_73
timestamp 1676037725
transform 1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_79
timestamp 1676037725
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_91
timestamp 1676037725
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_99
timestamp 1676037725
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_105
timestamp 1676037725
transform 1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1676037725
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1676037725
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1676037725
transform 1 0 14812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1676037725
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1676037725
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_235
timestamp 1676037725
transform 1 0 22724 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1676037725
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_261
timestamp 1676037725
transform 1 0 25116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_8
timestamp 1676037725
transform 1 0 1840 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_12
timestamp 1676037725
transform 1 0 2208 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_24
timestamp 1676037725
transform 1 0 3312 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_36
timestamp 1676037725
transform 1 0 4416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 1676037725
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_59
timestamp 1676037725
transform 1 0 6532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_71
timestamp 1676037725
transform 1 0 7636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_83
timestamp 1676037725
transform 1 0 8740 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_95
timestamp 1676037725
transform 1 0 9844 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_98
timestamp 1676037725
transform 1 0 10120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1676037725
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp 1676037725
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_151
timestamp 1676037725
transform 1 0 14996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_159
timestamp 1676037725
transform 1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1676037725
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1676037725
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_263
timestamp 1676037725
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_5
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_17
timestamp 1676037725
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1676037725
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1676037725
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1676037725
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_235
timestamp 1676037725
transform 1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1676037725
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_259
timestamp 1676037725
transform 1 0 24932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1676037725
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1676037725
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1676037725
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1676037725
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1676037725
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1676037725
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_227
timestamp 1676037725
transform 1 0 21988 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1676037725
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_185
timestamp 1676037725
transform 1 0 18124 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1676037725
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_243
timestamp 1676037725
transform 1 0 23460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_247
timestamp 1676037725
transform 1 0 23828 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_203
timestamp 1676037725
transform 1 0 19780 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp 1676037725
transform 1 0 20516 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1676037725
transform 1 0 18492 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_195
timestamp 1676037725
transform 1 0 19044 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_203
timestamp 1676037725
transform 1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_55
timestamp 1676037725
transform 1 0 6164 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_59
timestamp 1676037725
transform 1 0 6532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_71
timestamp 1676037725
transform 1 0 7636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_205
timestamp 1676037725
transform 1 0 19964 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_211
timestamp 1676037725
transform 1 0 20516 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_220
timestamp 1676037725
transform 1 0 21344 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_232
timestamp 1676037725
transform 1 0 22448 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_71
timestamp 1676037725
transform 1 0 7636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_83
timestamp 1676037725
transform 1 0 8740 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_95
timestamp 1676037725
transform 1 0 9844 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1676037725
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_199
timestamp 1676037725
transform 1 0 19412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_211
timestamp 1676037725
transform 1 0 20516 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 1676037725
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_225
timestamp 1676037725
transform 1 0 21804 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_237
timestamp 1676037725
transform 1 0 22908 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1676037725
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_68
timestamp 1676037725
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_80
timestamp 1676037725
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_92
timestamp 1676037725
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1676037725
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_175
timestamp 1676037725
transform 1 0 17204 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_198
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_210
timestamp 1676037725
transform 1 0 20424 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_233
timestamp 1676037725
transform 1 0 22540 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_238
timestamp 1676037725
transform 1 0 23000 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_246
timestamp 1676037725
transform 1 0 23736 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1676037725
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1676037725
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_150
timestamp 1676037725
transform 1 0 14904 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_162
timestamp 1676037725
transform 1 0 16008 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_168
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_173
timestamp 1676037725
transform 1 0 17020 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_185
timestamp 1676037725
transform 1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1676037725
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1676037725
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_222
timestamp 1676037725
transform 1 0 21528 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_226
timestamp 1676037725
transform 1 0 21896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1676037725
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_259
timestamp 1676037725
transform 1 0 24932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1676037725
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_122
timestamp 1676037725
transform 1 0 12328 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_134
timestamp 1676037725
transform 1 0 13432 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_146
timestamp 1676037725
transform 1 0 14536 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_150
timestamp 1676037725
transform 1 0 14904 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1676037725
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1676037725
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_189
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_195
timestamp 1676037725
transform 1 0 19044 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_205
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_212
timestamp 1676037725
transform 1 0 20608 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_243
timestamp 1676037725
transform 1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_247
timestamp 1676037725
transform 1 0 23828 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1676037725
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_155
timestamp 1676037725
transform 1 0 15364 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_204
timestamp 1676037725
transform 1 0 19872 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_212
timestamp 1676037725
transform 1 0 20608 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_217
timestamp 1676037725
transform 1 0 21068 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_229
timestamp 1676037725
transform 1 0 22172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_241
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1676037725
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1676037725
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_160
timestamp 1676037725
transform 1 0 15824 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1676037725
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1676037725
transform 1 0 17204 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_179
timestamp 1676037725
transform 1 0 17572 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1676037725
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp 1676037725
transform 1 0 20056 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1676037725
transform 1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1676037725
transform 1 0 21160 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_245
timestamp 1676037725
transform 1 0 23644 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1676037725
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_137
timestamp 1676037725
transform 1 0 13708 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1676037725
transform 1 0 15272 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_173
timestamp 1676037725
transform 1 0 17020 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_199
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_207
timestamp 1676037725
transform 1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_226
timestamp 1676037725
transform 1 0 21896 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_238
timestamp 1676037725
transform 1 0 23000 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1676037725
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_265
timestamp 1676037725
transform 1 0 25484 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_86
timestamp 1676037725
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_115
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_127
timestamp 1676037725
transform 1 0 12788 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_135
timestamp 1676037725
transform 1 0 13524 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1676037725
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_148
timestamp 1676037725
transform 1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1676037725
transform 1 0 15088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_158
timestamp 1676037725
transform 1 0 15640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_162
timestamp 1676037725
transform 1 0 16008 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_192
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_196
timestamp 1676037725
transform 1 0 19136 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_245
timestamp 1676037725
transform 1 0 23644 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_264
timestamp 1676037725
transform 1 0 25392 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_61
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1676037725
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_87
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_120
timestamp 1676037725
transform 1 0 12144 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1676037725
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1676037725
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1676037725
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1676037725
transform 1 0 16376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_170
timestamp 1676037725
transform 1 0 16744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_174
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_180
timestamp 1676037725
transform 1 0 17664 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1676037725
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1676037725
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_212
timestamp 1676037725
transform 1 0 20608 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_215
timestamp 1676037725
transform 1 0 20884 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_221
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_224
timestamp 1676037725
transform 1 0 21712 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_232
timestamp 1676037725
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_95
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_99
timestamp 1676037725
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_130
timestamp 1676037725
transform 1 0 13064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_138
timestamp 1676037725
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_142
timestamp 1676037725
transform 1 0 14168 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_154
timestamp 1676037725
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1676037725
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_194
timestamp 1676037725
transform 1 0 18952 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_213
timestamp 1676037725
transform 1 0 20700 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1676037725
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_227
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_235
timestamp 1676037725
transform 1 0 22724 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_241
timestamp 1676037725
transform 1 0 23276 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_247
timestamp 1676037725
transform 1 0 23828 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1676037725
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1676037725
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_120
timestamp 1676037725
transform 1 0 12144 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_124
timestamp 1676037725
transform 1 0 12512 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_127
timestamp 1676037725
transform 1 0 12788 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_143
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_179
timestamp 1676037725
transform 1 0 17572 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_187
timestamp 1676037725
transform 1 0 18308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1676037725
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_202
timestamp 1676037725
transform 1 0 19688 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_207
timestamp 1676037725
transform 1 0 20148 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_235
timestamp 1676037725
transform 1 0 22724 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_239
timestamp 1676037725
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_115
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1676037725
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1676037725
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_151
timestamp 1676037725
transform 1 0 14996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1676037725
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1676037725
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1676037725
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_178
timestamp 1676037725
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_182
timestamp 1676037725
transform 1 0 17848 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1676037725
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_204
timestamp 1676037725
transform 1 0 19872 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_216
timestamp 1676037725
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_229
timestamp 1676037725
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_233
timestamp 1676037725
transform 1 0 22540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_245
timestamp 1676037725
transform 1 0 23644 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8004 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1676037725
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_105
timestamp 1676037725
transform 1 0 10764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_129
timestamp 1676037725
transform 1 0 12972 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1676037725
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_152
timestamp 1676037725
transform 1 0 15088 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_164
timestamp 1676037725
transform 1 0 16192 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_185
timestamp 1676037725
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_208
timestamp 1676037725
transform 1 0 20240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1676037725
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1676037725
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_223
timestamp 1676037725
transform 1 0 21620 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_228
timestamp 1676037725
transform 1 0 22080 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_11
timestamp 1676037725
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_18
timestamp 1676037725
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_30
timestamp 1676037725
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_42
timestamp 1676037725
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_80
timestamp 1676037725
transform 1 0 8464 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_84
timestamp 1676037725
transform 1 0 8832 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_94
timestamp 1676037725
transform 1 0 9752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1676037725
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_124
timestamp 1676037725
transform 1 0 12512 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_128
timestamp 1676037725
transform 1 0 12880 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_131
timestamp 1676037725
transform 1 0 13156 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1676037725
transform 1 0 13892 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_145
timestamp 1676037725
transform 1 0 14444 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_157
timestamp 1676037725
transform 1 0 15548 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_164
timestamp 1676037725
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_171
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1676037725
transform 1 0 17572 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_191
timestamp 1676037725
transform 1 0 18676 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_195
timestamp 1676037725
transform 1 0 19044 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_213
timestamp 1676037725
transform 1 0 20700 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1676037725
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_243
timestamp 1676037725
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1676037725
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_45
timestamp 1676037725
transform 1 0 5244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_66
timestamp 1676037725
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_70
timestamp 1676037725
transform 1 0 7544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_96
timestamp 1676037725
transform 1 0 9936 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_111
timestamp 1676037725
transform 1 0 11316 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_115
timestamp 1676037725
transform 1 0 11684 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1676037725
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_167
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_179
timestamp 1676037725
transform 1 0 17572 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1676037725
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_205
timestamp 1676037725
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1676037725
transform 1 0 20884 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_223
timestamp 1676037725
transform 1 0 21620 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_244
timestamp 1676037725
transform 1 0 23552 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1676037725
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_263
timestamp 1676037725
transform 1 0 25300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_82
timestamp 1676037725
transform 1 0 8648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_92
timestamp 1676037725
transform 1 0 9568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_96
timestamp 1676037725
transform 1 0 9936 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_106
timestamp 1676037725
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_152
timestamp 1676037725
transform 1 0 15088 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_160
timestamp 1676037725
transform 1 0 15824 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1676037725
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_174
timestamp 1676037725
transform 1 0 17112 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_200
timestamp 1676037725
transform 1 0 19504 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_204
timestamp 1676037725
transform 1 0 19872 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_213
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_217
timestamp 1676037725
transform 1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_221
timestamp 1676037725
transform 1 0 21436 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_231
timestamp 1676037725
transform 1 0 22356 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_239
timestamp 1676037725
transform 1 0 23092 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_247
timestamp 1676037725
transform 1 0 23828 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1676037725
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_78
timestamp 1676037725
transform 1 0 8280 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_96
timestamp 1676037725
transform 1 0 9936 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_113
timestamp 1676037725
transform 1 0 11500 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_120
timestamp 1676037725
transform 1 0 12144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_124
timestamp 1676037725
transform 1 0 12512 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1676037725
transform 1 0 12788 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_160
timestamp 1676037725
transform 1 0 15824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_173
timestamp 1676037725
transform 1 0 17020 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_203
timestamp 1676037725
transform 1 0 19780 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_224
timestamp 1676037725
transform 1 0 21712 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_248
timestamp 1676037725
transform 1 0 23920 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_259
timestamp 1676037725
transform 1 0 24932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_265
timestamp 1676037725
transform 1 0 25484 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_65
timestamp 1676037725
transform 1 0 7084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_76
timestamp 1676037725
transform 1 0 8096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1676037725
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_95
timestamp 1676037725
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1676037725
transform 1 0 10212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_124
timestamp 1676037725
transform 1 0 12512 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_132
timestamp 1676037725
transform 1 0 13248 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_141
timestamp 1676037725
transform 1 0 14076 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_152
timestamp 1676037725
transform 1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_156
timestamp 1676037725
transform 1 0 15456 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1676037725
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_176
timestamp 1676037725
transform 1 0 17296 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_189
timestamp 1676037725
transform 1 0 18492 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_213
timestamp 1676037725
transform 1 0 20700 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_217
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 20148 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_244
timestamp 1676037725
transform 1 0 23552 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_89
timestamp 1676037725
transform 1 0 9292 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_92
timestamp 1676037725
transform 1 0 9568 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_152
timestamp 1676037725
transform 1 0 15088 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_185
timestamp 1676037725
transform 1 0 18124 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_191
timestamp 1676037725
transform 1 0 18676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_204
timestamp 1676037725
transform 1 0 19872 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_208
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_220
timestamp 1676037725
transform 1 0 21344 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_224
timestamp 1676037725
transform 1 0 21712 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_255
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_263
timestamp 1676037725
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_9
timestamp 1676037725
transform 1 0 1932 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_13
timestamp 1676037725
transform 1 0 2300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_25
timestamp 1676037725
transform 1 0 3404 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_33
timestamp 1676037725
transform 1 0 4140 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_37
timestamp 1676037725
transform 1 0 4508 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1676037725
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_92
timestamp 1676037725
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_104
timestamp 1676037725
transform 1 0 10672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_124
timestamp 1676037725
transform 1 0 12512 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_130
timestamp 1676037725
transform 1 0 13064 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_133
timestamp 1676037725
transform 1 0 13340 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_148
timestamp 1676037725
transform 1 0 14720 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1676037725
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1676037725
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_187
timestamp 1676037725
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_195
timestamp 1676037725
transform 1 0 19044 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_208
timestamp 1676037725
transform 1 0 20240 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_212
timestamp 1676037725
transform 1 0 20608 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_247
timestamp 1676037725
transform 1 0 23828 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_251
timestamp 1676037725
transform 1 0 24196 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_263
timestamp 1676037725
transform 1 0 25300 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_46
timestamp 1676037725
transform 1 0 5336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_70
timestamp 1676037725
transform 1 0 7544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_74
timestamp 1676037725
transform 1 0 7912 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_78
timestamp 1676037725
transform 1 0 8280 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_114
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_124
timestamp 1676037725
transform 1 0 12512 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_136
timestamp 1676037725
transform 1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_152
timestamp 1676037725
transform 1 0 15088 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_156
timestamp 1676037725
transform 1 0 15456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_168
timestamp 1676037725
transform 1 0 16560 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_178
timestamp 1676037725
transform 1 0 17480 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_184
timestamp 1676037725
transform 1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_188
timestamp 1676037725
transform 1 0 18400 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_199
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_207
timestamp 1676037725
transform 1 0 20148 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_210
timestamp 1676037725
transform 1 0 20424 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_222
timestamp 1676037725
transform 1 0 21528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1676037725
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_79
timestamp 1676037725
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_92
timestamp 1676037725
transform 1 0 9568 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_128
timestamp 1676037725
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_139
timestamp 1676037725
transform 1 0 13892 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1676037725
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1676037725
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_177
timestamp 1676037725
transform 1 0 17388 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_183
timestamp 1676037725
transform 1 0 17940 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_190
timestamp 1676037725
transform 1 0 18584 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_203
timestamp 1676037725
transform 1 0 19780 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_215
timestamp 1676037725
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_244
timestamp 1676037725
transform 1 0 23552 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1676037725
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_9
timestamp 1676037725
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_13
timestamp 1676037725
transform 1 0 2300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_17
timestamp 1676037725
transform 1 0 2668 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_35
timestamp 1676037725
transform 1 0 4324 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_59
timestamp 1676037725
transform 1 0 6532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_71
timestamp 1676037725
transform 1 0 7636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_93
timestamp 1676037725
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_115
timestamp 1676037725
transform 1 0 11684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_119
timestamp 1676037725
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_131
timestamp 1676037725
transform 1 0 13156 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_137
timestamp 1676037725
transform 1 0 13708 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_160
timestamp 1676037725
transform 1 0 15824 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_166
timestamp 1676037725
transform 1 0 16376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_170
timestamp 1676037725
transform 1 0 16744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp 1676037725
transform 1 0 17020 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_184
timestamp 1676037725
transform 1 0 18032 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_190
timestamp 1676037725
transform 1 0 18584 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_203
timestamp 1676037725
transform 1 0 19780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_224
timestamp 1676037725
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_228
timestamp 1676037725
transform 1 0 22080 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_33
timestamp 1676037725
transform 1 0 4140 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1676037725
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_74
timestamp 1676037725
transform 1 0 7912 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_87
timestamp 1676037725
transform 1 0 9108 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_100
timestamp 1676037725
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_124
timestamp 1676037725
transform 1 0 12512 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_132
timestamp 1676037725
transform 1 0 13248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_144
timestamp 1676037725
transform 1 0 14352 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_148
timestamp 1676037725
transform 1 0 14720 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_158
timestamp 1676037725
transform 1 0 15640 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1676037725
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_174
timestamp 1676037725
transform 1 0 17112 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_183
timestamp 1676037725
transform 1 0 17940 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_192
timestamp 1676037725
transform 1 0 18768 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_204
timestamp 1676037725
transform 1 0 19872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_208
timestamp 1676037725
transform 1 0 20240 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_211
timestamp 1676037725
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1676037725
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1676037725
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_262
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_37
timestamp 1676037725
transform 1 0 4508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_49
timestamp 1676037725
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_61
timestamp 1676037725
transform 1 0 6716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_73
timestamp 1676037725
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1676037725
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_105
timestamp 1676037725
transform 1 0 10764 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_110
timestamp 1676037725
transform 1 0 11224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1676037725
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_129
timestamp 1676037725
transform 1 0 12972 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1676037725
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_163
timestamp 1676037725
transform 1 0 16100 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_169
timestamp 1676037725
transform 1 0 16652 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1676037725
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 1676037725
transform 1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_223
timestamp 1676037725
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_259
timestamp 1676037725
transform 1 0 24932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_265
timestamp 1676037725
transform 1 0 24932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_263
timestamp 1676037725
transform 1 0 25300 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_9
timestamp 1676037725
transform 1 0 1932 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_13
timestamp 1676037725
transform 1 0 2300 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_25
timestamp 1676037725
transform 1 0 3404 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_37
timestamp 1676037725
transform 1 0 4508 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_61
timestamp 1676037725
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_71
timestamp 1676037725
transform 1 0 7636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_86
timestamp 1676037725
transform 1 0 9016 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_90
timestamp 1676037725
transform 1 0 9384 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_96
timestamp 1676037725
transform 1 0 9936 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_99
timestamp 1676037725
transform 1 0 10212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_116
timestamp 1676037725
transform 1 0 11776 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_127
timestamp 1676037725
transform 1 0 12788 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_131
timestamp 1676037725
transform 1 0 13156 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_142
timestamp 1676037725
transform 1 0 14168 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_157
timestamp 1676037725
transform 1 0 15548 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1676037725
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_177
timestamp 1676037725
transform 1 0 17388 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_180
timestamp 1676037725
transform 1 0 17664 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_206
timestamp 1676037725
transform 1 0 20056 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_210
timestamp 1676037725
transform 1 0 20424 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_248
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_254
timestamp 1676037725
transform 1 0 24472 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1676037725
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_263
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_9
timestamp 1676037725
transform 1 0 1932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_13
timestamp 1676037725
transform 1 0 2300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_17
timestamp 1676037725
transform 1 0 2668 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1676037725
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_36
timestamp 1676037725
transform 1 0 4416 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_47
timestamp 1676037725
transform 1 0 5428 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_71
timestamp 1676037725
transform 1 0 7636 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_75
timestamp 1676037725
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_93
timestamp 1676037725
transform 1 0 9660 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_107
timestamp 1676037725
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_120
timestamp 1676037725
transform 1 0 12144 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_127
timestamp 1676037725
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_163
timestamp 1676037725
transform 1 0 16100 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_187
timestamp 1676037725
transform 1 0 18308 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_191
timestamp 1676037725
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_219
timestamp 1676037725
transform 1 0 21252 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_223
timestamp 1676037725
transform 1 0 21620 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_230
timestamp 1676037725
transform 1 0 22356 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_21
timestamp 1676037725
transform 1 0 3036 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_33
timestamp 1676037725
transform 1 0 4140 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_59
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_91
timestamp 1676037725
transform 1 0 9476 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_98
timestamp 1676037725
transform 1 0 10120 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_102
timestamp 1676037725
transform 1 0 10488 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1676037725
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_115
timestamp 1676037725
transform 1 0 11684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1676037725
transform 1 0 11960 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_126
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_140
timestamp 1676037725
transform 1 0 13984 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_152
timestamp 1676037725
transform 1 0 15088 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1676037725
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_176
timestamp 1676037725
transform 1 0 17296 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1676037725
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_215
timestamp 1676037725
transform 1 0 20884 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_219
timestamp 1676037725
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_257
timestamp 1676037725
transform 1 0 24748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1676037725
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_13
timestamp 1676037725
transform 1 0 2300 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_18
timestamp 1676037725
transform 1 0 2760 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_51
timestamp 1676037725
transform 1 0 5796 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_58
timestamp 1676037725
transform 1 0 6440 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_74
timestamp 1676037725
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 1676037725
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_99
timestamp 1676037725
transform 1 0 10212 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_103
timestamp 1676037725
transform 1 0 10580 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_114
timestamp 1676037725
transform 1 0 11592 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_127
timestamp 1676037725
transform 1 0 12788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_134
timestamp 1676037725
transform 1 0 13432 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_146
timestamp 1676037725
transform 1 0 14536 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_158
timestamp 1676037725
transform 1 0 15640 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_175
timestamp 1676037725
transform 1 0 17204 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_182
timestamp 1676037725
transform 1 0 17848 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_201
timestamp 1676037725
transform 1 0 19596 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_230
timestamp 1676037725
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_48
timestamp 1676037725
transform 1 0 5520 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1676037725
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_65
timestamp 1676037725
transform 1 0 7084 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_80
timestamp 1676037725
transform 1 0 8464 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_100
timestamp 1676037725
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1676037725
transform 1 0 11960 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_124
timestamp 1676037725
transform 1 0 12512 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_132
timestamp 1676037725
transform 1 0 13248 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_143
timestamp 1676037725
transform 1 0 14260 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1676037725
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1676037725
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_201
timestamp 1676037725
transform 1 0 19596 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_206
timestamp 1676037725
transform 1 0 20056 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_257
timestamp 1676037725
transform 1 0 24748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1676037725
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3404 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_34
timestamp 1676037725
transform 1 0 4232 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_46
timestamp 1676037725
transform 1 0 5336 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_58
timestamp 1676037725
transform 1 0 6440 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1676037725
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_87
timestamp 1676037725
transform 1 0 9108 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_93
timestamp 1676037725
transform 1 0 9660 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_106
timestamp 1676037725
transform 1 0 10856 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_110
timestamp 1676037725
transform 1 0 11224 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1676037725
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_147
timestamp 1676037725
transform 1 0 14628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_157
timestamp 1676037725
transform 1 0 15548 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_181
timestamp 1676037725
transform 1 0 17756 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_187
timestamp 1676037725
transform 1 0 18308 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_208
timestamp 1676037725
transform 1 0 20240 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_220
timestamp 1676037725
transform 1 0 21344 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_237
timestamp 1676037725
transform 1 0 22908 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_243
timestamp 1676037725
transform 1 0 23460 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_259
timestamp 1676037725
transform 1 0 24932 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_263
timestamp 1676037725
transform 1 0 25300 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_14
timestamp 1676037725
transform 1 0 2392 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_20
timestamp 1676037725
transform 1 0 2944 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_29
timestamp 1676037725
transform 1 0 3772 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_78
timestamp 1676037725
transform 1 0 8280 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_82
timestamp 1676037725
transform 1 0 8648 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_86
timestamp 1676037725
transform 1 0 9016 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_97
timestamp 1676037725
transform 1 0 10028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1676037725
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_117
timestamp 1676037725
transform 1 0 11868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_121
timestamp 1676037725
transform 1 0 12236 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_146
timestamp 1676037725
transform 1 0 14536 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_150
timestamp 1676037725
transform 1 0 14904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_154
timestamp 1676037725
transform 1 0 15272 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1676037725
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_177
timestamp 1676037725
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_200
timestamp 1676037725
transform 1 0 19504 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_213
timestamp 1676037725
transform 1 0 20700 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1676037725
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_236
timestamp 1676037725
transform 1 0 22816 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_244
timestamp 1676037725
transform 1 0 23552 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_264
timestamp 1676037725
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1676037725
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_33
timestamp 1676037725
transform 1 0 4140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_45
timestamp 1676037725
transform 1 0 5244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_57
timestamp 1676037725
transform 1 0 6348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_78
timestamp 1676037725
transform 1 0 8280 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_90
timestamp 1676037725
transform 1 0 9384 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_116
timestamp 1676037725
transform 1 0 11776 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_129
timestamp 1676037725
transform 1 0 12972 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1676037725
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_146
timestamp 1676037725
transform 1 0 14536 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_154
timestamp 1676037725
transform 1 0 15272 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_175
timestamp 1676037725
transform 1 0 17204 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_179
timestamp 1676037725
transform 1 0 17572 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_191
timestamp 1676037725
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_208
timestamp 1676037725
transform 1 0 20240 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_232
timestamp 1676037725
transform 1 0 22448 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_245
timestamp 1676037725
transform 1 0 23644 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1676037725
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_259
timestamp 1676037725
transform 1 0 24932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_263
timestamp 1676037725
transform 1 0 25300 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_24
timestamp 1676037725
transform 1 0 3312 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_49
timestamp 1676037725
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_79
timestamp 1676037725
transform 1 0 8372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_92
timestamp 1676037725
transform 1 0 9568 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_100
timestamp 1676037725
transform 1 0 10304 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_118
timestamp 1676037725
transform 1 0 11960 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_144
timestamp 1676037725
transform 1 0 14352 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_157
timestamp 1676037725
transform 1 0 15548 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1676037725
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_177
timestamp 1676037725
transform 1 0 17388 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_188
timestamp 1676037725
transform 1 0 18400 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_209
timestamp 1676037725
transform 1 0 20332 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_216
timestamp 1676037725
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_232
timestamp 1676037725
transform 1 0 22448 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_256
timestamp 1676037725
transform 1 0 24656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_264
timestamp 1676037725
transform 1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_75
timestamp 1676037725
transform 1 0 8004 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1676037725
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_129
timestamp 1676037725
transform 1 0 12972 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_149
timestamp 1676037725
transform 1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_161
timestamp 1676037725
transform 1 0 15916 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_167
timestamp 1676037725
transform 1 0 16468 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_179
timestamp 1676037725
transform 1 0 17572 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_188
timestamp 1676037725
transform 1 0 18400 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_201
timestamp 1676037725
transform 1 0 19596 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_204
timestamp 1676037725
transform 1 0 19872 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_215
timestamp 1676037725
transform 1 0 20884 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_223
timestamp 1676037725
transform 1 0 21620 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_247
timestamp 1676037725
transform 1 0 23828 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_259
timestamp 1676037725
transform 1 0 24932 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_263
timestamp 1676037725
transform 1 0 25300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_9
timestamp 1676037725
transform 1 0 1932 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_13
timestamp 1676037725
transform 1 0 2300 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_25
timestamp 1676037725
transform 1 0 3404 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_30
timestamp 1676037725
transform 1 0 3864 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_42
timestamp 1676037725
transform 1 0 4968 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1676037725
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_77
timestamp 1676037725
transform 1 0 8188 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_98
timestamp 1676037725
transform 1 0 10120 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_102
timestamp 1676037725
transform 1 0 10488 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1676037725
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_128
timestamp 1676037725
transform 1 0 12880 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_134
timestamp 1676037725
transform 1 0 13432 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_146
timestamp 1676037725
transform 1 0 14536 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_47_154
timestamp 1676037725
transform 1 0 15272 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1676037725
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_173
timestamp 1676037725
transform 1 0 17020 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_177
timestamp 1676037725
transform 1 0 17388 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_180
timestamp 1676037725
transform 1 0 17664 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_191
timestamp 1676037725
transform 1 0 18676 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_204
timestamp 1676037725
transform 1 0 19872 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_208
timestamp 1676037725
transform 1 0 20240 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_212
timestamp 1676037725
transform 1 0 20608 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_220
timestamp 1676037725
transform 1 0 21344 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_248
timestamp 1676037725
transform 1 0 23920 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_252
timestamp 1676037725
transform 1 0 24288 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_259
timestamp 1676037725
transform 1 0 24932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_263
timestamp 1676037725
transform 1 0 25300 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1676037725
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_33
timestamp 1676037725
transform 1 0 4140 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_55
timestamp 1676037725
transform 1 0 6164 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_79
timestamp 1676037725
transform 1 0 8372 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_123
timestamp 1676037725
transform 1 0 12420 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_136
timestamp 1676037725
transform 1 0 13616 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_152
timestamp 1676037725
transform 1 0 15088 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_156
timestamp 1676037725
transform 1 0 15456 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_167
timestamp 1676037725
transform 1 0 16468 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_171
timestamp 1676037725
transform 1 0 16836 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_184
timestamp 1676037725
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_219
timestamp 1676037725
transform 1 0 21252 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_223
timestamp 1676037725
transform 1 0 21620 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_235
timestamp 1676037725
transform 1 0 22724 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1676037725
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_258
timestamp 1676037725
transform 1 0 24840 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_92
timestamp 1676037725
transform 1 0 9568 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_96
timestamp 1676037725
transform 1 0 10396 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp 1676037725
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_121
timestamp 1676037725
transform 1 0 12236 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_133
timestamp 1676037725
transform 1 0 13340 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1676037725
transform 1 0 14536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_159
timestamp 1676037725
transform 1 0 15732 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_165
timestamp 1676037725
transform 1 0 16284 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_180
timestamp 1676037725
transform 1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_186
timestamp 1676037725
transform 1 0 18216 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_198
timestamp 1676037725
transform 1 0 19320 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_204
timestamp 1676037725
transform 1 0 19872 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_215
timestamp 1676037725
transform 1 0 20884 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_219
timestamp 1676037725
transform 1 0 21252 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_236
timestamp 1676037725
transform 1 0 22816 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_246
timestamp 1676037725
transform 1 0 23736 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_251
timestamp 1676037725
transform 1 0 24196 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_259
timestamp 1676037725
transform 1 0 24932 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_33
timestamp 1676037725
transform 1 0 4140 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_55
timestamp 1676037725
transform 1 0 6164 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_71
timestamp 1676037725
transform 1 0 7636 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1676037725
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_89
timestamp 1676037725
transform 1 0 9292 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_100
timestamp 1676037725
transform 1 0 10304 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_134
timestamp 1676037725
transform 1 0 13432 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1676037725
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_147
timestamp 1676037725
transform 1 0 14628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1676037725
transform 1 0 16560 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_181
timestamp 1676037725
transform 1 0 17756 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1676037725
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_210
timestamp 1676037725
transform 1 0 20424 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_214
timestamp 1676037725
transform 1 0 20792 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_218
timestamp 1676037725
transform 1 0 21160 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_231
timestamp 1676037725
transform 1 0 22356 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1676037725
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1676037725
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_93
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_99
timestamp 1676037725
transform 1 0 10212 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1676037725
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_118
timestamp 1676037725
transform 1 0 11960 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1676037725
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_175
timestamp 1676037725
transform 1 0 17204 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_188
timestamp 1676037725
transform 1 0 18400 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_194
timestamp 1676037725
transform 1 0 18952 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_198
timestamp 1676037725
transform 1 0 19320 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_202
timestamp 1676037725
transform 1 0 19688 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1676037725
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_237
timestamp 1676037725
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_241
timestamp 1676037725
transform 1 0 23276 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_262
timestamp 1676037725
transform 1 0 25208 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_52
timestamp 1676037725
transform 1 0 5888 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_64
timestamp 1676037725
transform 1 0 6992 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_72
timestamp 1676037725
transform 1 0 7728 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1676037725
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1676037725
transform 1 0 9476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_112
timestamp 1676037725
transform 1 0 11408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_116
timestamp 1676037725
transform 1 0 11776 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_122
timestamp 1676037725
transform 1 0 12328 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_125
timestamp 1676037725
transform 1 0 12604 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_136
timestamp 1676037725
transform 1 0 13616 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_159
timestamp 1676037725
transform 1 0 15732 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_162
timestamp 1676037725
transform 1 0 16008 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_184
timestamp 1676037725
transform 1 0 18032 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_188
timestamp 1676037725
transform 1 0 18400 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_208
timestamp 1676037725
transform 1 0 20240 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_212
timestamp 1676037725
transform 1 0 20608 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_224
timestamp 1676037725
transform 1 0 21712 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_236
timestamp 1676037725
transform 1 0 22816 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_240
timestamp 1676037725
transform 1 0 23184 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_244
timestamp 1676037725
transform 1 0 23552 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1676037725
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_259
timestamp 1676037725
transform 1 0 24932 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_264
timestamp 1676037725
transform 1 0 25392 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_21
timestamp 1676037725
transform 1 0 3036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1676037725
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1676037725
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1676037725
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_67
timestamp 1676037725
transform 1 0 7268 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_78
timestamp 1676037725
transform 1 0 8280 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_91
timestamp 1676037725
transform 1 0 9476 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_103
timestamp 1676037725
transform 1 0 10580 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_148
timestamp 1676037725
transform 1 0 14720 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_152
timestamp 1676037725
transform 1 0 15088 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1676037725
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_172
timestamp 1676037725
transform 1 0 16928 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_183
timestamp 1676037725
transform 1 0 17940 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1676037725
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_209
timestamp 1676037725
transform 1 0 20332 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_215
timestamp 1676037725
transform 1 0 20884 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_249
timestamp 1676037725
transform 1 0 24012 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1676037725
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_260
timestamp 1676037725
transform 1 0 25024 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_75
timestamp 1676037725
transform 1 0 8004 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_79
timestamp 1676037725
transform 1 0 8372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_89
timestamp 1676037725
transform 1 0 9292 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_110
timestamp 1676037725
transform 1 0 11224 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_114
timestamp 1676037725
transform 1 0 11592 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_126
timestamp 1676037725
transform 1 0 12696 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_152
timestamp 1676037725
transform 1 0 15088 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_164
timestamp 1676037725
transform 1 0 16192 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_175
timestamp 1676037725
transform 1 0 17204 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_185
timestamp 1676037725
transform 1 0 17848 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_209
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_208
timestamp 1676037725
transform 1 0 20240 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_221
timestamp 1676037725
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_225
timestamp 1676037725
transform 1 0 21804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_235
timestamp 1676037725
transform 1 0 22724 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_247
timestamp 1676037725
transform 1 0 23828 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_259
timestamp 1676037725
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_264
timestamp 1676037725
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_35
timestamp 1676037725
transform 1 0 4324 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_40
timestamp 1676037725
transform 1 0 4784 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_66
timestamp 1676037725
transform 1 0 7176 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_91
timestamp 1676037725
transform 1 0 9476 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_98
timestamp 1676037725
transform 1 0 10120 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_102
timestamp 1676037725
transform 1 0 10488 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1676037725
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_116
timestamp 1676037725
transform 1 0 11776 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_127
timestamp 1676037725
transform 1 0 12788 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_134
timestamp 1676037725
transform 1 0 13432 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_180
timestamp 1676037725
transform 1 0 17664 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1676037725
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_205
timestamp 1676037725
transform 1 0 19964 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_209
timestamp 1676037725
transform 1 0 20332 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1676037725
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_227
timestamp 1676037725
transform 1 0 21988 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_232
timestamp 1676037725
transform 1 0 22448 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_239
timestamp 1676037725
transform 1 0 23092 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_243
timestamp 1676037725
transform 1 0 23460 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_255
timestamp 1676037725
transform 1 0 24564 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_259
timestamp 1676037725
transform 1 0 24932 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_264
timestamp 1676037725
transform 1 0 25392 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_78
timestamp 1676037725
transform 1 0 8280 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_89
timestamp 1676037725
transform 1 0 9292 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_99
timestamp 1676037725
transform 1 0 10212 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_107
timestamp 1676037725
transform 1 0 10948 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_118
timestamp 1676037725
transform 1 0 11960 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_130
timestamp 1676037725
transform 1 0 13064 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1676037725
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_152
timestamp 1676037725
transform 1 0 15088 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_158
timestamp 1676037725
transform 1 0 15640 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_161
timestamp 1676037725
transform 1 0 15916 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_172
timestamp 1676037725
transform 1 0 16928 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_178
timestamp 1676037725
transform 1 0 17480 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_190
timestamp 1676037725
transform 1 0 18584 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_201
timestamp 1676037725
transform 1 0 19596 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_212
timestamp 1676037725
transform 1 0 20608 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_225
timestamp 1676037725
transform 1 0 21804 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_232
timestamp 1676037725
transform 1 0 22448 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_238
timestamp 1676037725
transform 1 0 23000 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1676037725
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_259
timestamp 1676037725
transform 1 0 24932 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1676037725
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_8
timestamp 1676037725
transform 1 0 1840 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_12
timestamp 1676037725
transform 1 0 2208 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_24
timestamp 1676037725
transform 1 0 3312 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_36
timestamp 1676037725
transform 1 0 4416 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_44
timestamp 1676037725
transform 1 0 5152 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1676037725
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_67
timestamp 1676037725
transform 1 0 7268 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_79
timestamp 1676037725
transform 1 0 8372 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_91
timestamp 1676037725
transform 1 0 9476 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_97
timestamp 1676037725
transform 1 0 10028 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1676037725
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_121
timestamp 1676037725
transform 1 0 12236 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_126
timestamp 1676037725
transform 1 0 12696 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1676037725
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_204
timestamp 1676037725
transform 1 0 19872 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_217
timestamp 1676037725
transform 1 0 21068 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1676037725
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_230
timestamp 1676037725
transform 1 0 22264 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_237
timestamp 1676037725
transform 1 0 22172 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_232
timestamp 1676037725
transform 1 0 22448 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_240
timestamp 1676037725
transform 1 0 23184 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1676037725
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_47
timestamp 1676037725
transform 1 0 5428 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_68
timestamp 1676037725
transform 1 0 7360 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_72
timestamp 1676037725
transform 1 0 7728 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1676037725
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_96
timestamp 1676037725
transform 1 0 9936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_100
timestamp 1676037725
transform 1 0 10304 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_125
timestamp 1676037725
transform 1 0 12604 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1676037725
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_143
timestamp 1676037725
transform 1 0 14260 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_155
timestamp 1676037725
transform 1 0 15364 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_181
timestamp 1676037725
transform 1 0 17756 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_185
timestamp 1676037725
transform 1 0 18124 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 1676037725
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_208
timestamp 1676037725
transform 1 0 20240 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_214
timestamp 1676037725
transform 1 0 20792 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_226
timestamp 1676037725
transform 1 0 21896 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_239
timestamp 1676037725
transform 1 0 23092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_258
timestamp 1676037725
transform 1 0 24840 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_80
timestamp 1676037725
transform 1 0 8464 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_104
timestamp 1676037725
transform 1 0 10672 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1676037725
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_135
timestamp 1676037725
transform 1 0 13524 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_139
timestamp 1676037725
transform 1 0 13892 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_151
timestamp 1676037725
transform 1 0 14996 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1676037725
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1676037725
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_236
timestamp 1676037725
transform 1 0 22816 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_256
timestamp 1676037725
transform 1 0 24656 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_260
timestamp 1676037725
transform 1 0 25024 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1676037725
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_74
timestamp 1676037725
transform 1 0 7912 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_78
timestamp 1676037725
transform 1 0 8280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_98
timestamp 1676037725
transform 1 0 10120 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_110
timestamp 1676037725
transform 1 0 11224 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_122
timestamp 1676037725
transform 1 0 12328 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_128
timestamp 1676037725
transform 1 0 12880 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1676037725
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_175
timestamp 1676037725
transform 1 0 17204 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_179
timestamp 1676037725
transform 1 0 17572 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_191
timestamp 1676037725
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_219
timestamp 1676037725
transform 1 0 21252 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_223
timestamp 1676037725
transform 1 0 21620 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_229
timestamp 1676037725
transform 1 0 22172 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1676037725
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_255
timestamp 1676037725
transform 1 0 24564 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_264
timestamp 1676037725
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_33
timestamp 1676037725
transform 1 0 4140 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1676037725
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_59
timestamp 1676037725
transform 1 0 6532 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_71
timestamp 1676037725
transform 1 0 7636 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_75
timestamp 1676037725
transform 1 0 8004 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_96
timestamp 1676037725
transform 1 0 9936 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_100
timestamp 1676037725
transform 1 0 10304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_135
timestamp 1676037725
transform 1 0 13524 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_139
timestamp 1676037725
transform 1 0 13892 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_148
timestamp 1676037725
transform 1 0 14720 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_160
timestamp 1676037725
transform 1 0 15824 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_177
timestamp 1676037725
transform 1 0 17388 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_199
timestamp 1676037725
transform 1 0 19412 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_212
timestamp 1676037725
transform 1 0 20608 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_216
timestamp 1676037725
transform 1 0 20976 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_231
timestamp 1676037725
transform 1 0 22356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_235
timestamp 1676037725
transform 1 0 22724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_260
timestamp 1676037725
transform 1 0 25024 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_8
timestamp 1676037725
transform 1 0 1840 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_12
timestamp 1676037725
transform 1 0 2208 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1676037725
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1676037725
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_96
timestamp 1676037725
transform 1 0 9936 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_108
timestamp 1676037725
transform 1 0 11040 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_124
timestamp 1676037725
transform 1 0 12512 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_135
timestamp 1676037725
transform 1 0 13524 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_152
timestamp 1676037725
transform 1 0 15088 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_158
timestamp 1676037725
transform 1 0 15640 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_161
timestamp 1676037725
transform 1 0 15916 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_172
timestamp 1676037725
transform 1 0 16928 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_179
timestamp 1676037725
transform 1 0 17572 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_191
timestamp 1676037725
transform 1 0 18676 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_208
timestamp 1676037725
transform 1 0 20240 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_223
timestamp 1676037725
transform 1 0 21620 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_235
timestamp 1676037725
transform 1 0 22724 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1676037725
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_259
timestamp 1676037725
transform 1 0 24932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1676037725
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_51
timestamp 1676037725
transform 1 0 5796 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_78
timestamp 1676037725
transform 1 0 8280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_84
timestamp 1676037725
transform 1 0 8832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_95
timestamp 1676037725
transform 1 0 9844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1676037725
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_115
timestamp 1676037725
transform 1 0 11684 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_129
timestamp 1676037725
transform 1 0 12972 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_142
timestamp 1676037725
transform 1 0 14168 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_155
timestamp 1676037725
transform 1 0 15364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_171
timestamp 1676037725
transform 1 0 16836 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_182
timestamp 1676037725
transform 1 0 17848 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_194
timestamp 1676037725
transform 1 0 18952 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_202
timestamp 1676037725
transform 1 0 19688 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1676037725
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1676037725
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_233
timestamp 1676037725
transform 1 0 22540 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_256
timestamp 1676037725
transform 1 0 24656 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_260
timestamp 1676037725
transform 1 0 25024 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1676037725
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_61
timestamp 1676037725
transform 1 0 6716 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1676037725
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_98
timestamp 1676037725
transform 1 0 10120 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_102
timestamp 1676037725
transform 1 0 10488 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_119
timestamp 1676037725
transform 1 0 12052 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_126
timestamp 1676037725
transform 1 0 12696 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1676037725
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_148
timestamp 1676037725
transform 1 0 14720 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_159
timestamp 1676037725
transform 1 0 15732 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_172
timestamp 1676037725
transform 1 0 16928 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_185
timestamp 1676037725
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_192
timestamp 1676037725
transform 1 0 18768 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_210
timestamp 1676037725
transform 1 0 20424 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_214
timestamp 1676037725
transform 1 0 20792 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_219
timestamp 1676037725
transform 1 0 21252 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_232
timestamp 1676037725
transform 1 0 22448 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_244
timestamp 1676037725
transform 1 0 23552 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_258
timestamp 1676037725
transform 1 0 24840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_264
timestamp 1676037725
transform 1 0 25392 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1676037725
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_82
timestamp 1676037725
transform 1 0 8648 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_88
timestamp 1676037725
transform 1 0 9200 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_93
timestamp 1676037725
transform 1 0 9752 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_106
timestamp 1676037725
transform 1 0 10856 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_118
timestamp 1676037725
transform 1 0 11960 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_131
timestamp 1676037725
transform 1 0 13156 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_138
timestamp 1676037725
transform 1 0 13800 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_142
timestamp 1676037725
transform 1 0 14168 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_147
timestamp 1676037725
transform 1 0 14628 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_160
timestamp 1676037725
transform 1 0 15824 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_180
timestamp 1676037725
transform 1 0 17664 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_184
timestamp 1676037725
transform 1 0 18032 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_192
timestamp 1676037725
transform 1 0 18768 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_203
timestamp 1676037725
transform 1 0 19780 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_207
timestamp 1676037725
transform 1 0 20148 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_236
timestamp 1676037725
transform 1 0 22816 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_242
timestamp 1676037725
transform 1 0 23368 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1676037725
transform 1 0 25024 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_8
timestamp 1676037725
transform 1 0 1840 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_12
timestamp 1676037725
transform 1 0 2208 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1676037725
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_67
timestamp 1676037725
transform 1 0 7268 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_71
timestamp 1676037725
transform 1 0 7636 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1676037725
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_110
timestamp 1676037725
transform 1 0 11224 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_116
timestamp 1676037725
transform 1 0 11776 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_126
timestamp 1676037725
transform 1 0 12696 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_152
timestamp 1676037725
transform 1 0 15088 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_160
timestamp 1676037725
transform 1 0 15824 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_181
timestamp 1676037725
transform 1 0 17756 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1676037725
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_208
timestamp 1676037725
transform 1 0 20240 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_236
timestamp 1676037725
transform 1 0 22816 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_249
timestamp 1676037725
transform 1 0 24012 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1676037725
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1676037725
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1676037725
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_65
timestamp 1676037725
transform 1 0 7084 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_69
timestamp 1676037725
transform 1 0 7636 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_79
timestamp 1676037725
transform 1 0 8188 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_84
timestamp 1676037725
transform 1 0 8832 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_96
timestamp 1676037725
transform 1 0 9936 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_100
timestamp 1676037725
transform 1 0 10304 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_110
timestamp 1676037725
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_115
timestamp 1676037725
transform 1 0 11684 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_139
timestamp 1676037725
transform 1 0 13892 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_146
timestamp 1676037725
transform 1 0 14536 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_159
timestamp 1676037725
transform 1 0 15732 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_163
timestamp 1676037725
transform 1 0 16100 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_174
timestamp 1676037725
transform 1 0 17112 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_182
timestamp 1676037725
transform 1 0 17848 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_192
timestamp 1676037725
transform 1 0 18768 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_218
timestamp 1676037725
transform 1 0 21160 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_248
timestamp 1676037725
transform 1 0 23920 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_252
timestamp 1676037725
transform 1 0 24288 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_257
timestamp 1676037725
transform 1 0 24748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_264
timestamp 1676037725
transform 1 0 25392 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_61
timestamp 1676037725
transform 1 0 6716 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_90
timestamp 1676037725
transform 1 0 9384 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_103
timestamp 1676037725
transform 1 0 10580 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_127
timestamp 1676037725
transform 1 0 12788 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_131
timestamp 1676037725
transform 1 0 13156 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_137
timestamp 1676037725
transform 1 0 13708 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_166
timestamp 1676037725
transform 1 0 16376 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_178
timestamp 1676037725
transform 1 0 17480 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_190
timestamp 1676037725
transform 1 0 18584 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_194
timestamp 1676037725
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_208
timestamp 1676037725
transform 1 0 20240 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_212
timestamp 1676037725
transform 1 0 20608 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_218
timestamp 1676037725
transform 1 0 21160 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_228
timestamp 1676037725
transform 1 0 22080 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_232
timestamp 1676037725
transform 1 0 22448 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_243
timestamp 1676037725
transform 1 0 23460 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1676037725
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1676037725
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_65
timestamp 1676037725
transform 1 0 7084 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_76
timestamp 1676037725
transform 1 0 8096 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_103
timestamp 1676037725
transform 1 0 10580 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_110
timestamp 1676037725
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_148
timestamp 1676037725
transform 1 0 14720 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_152
timestamp 1676037725
transform 1 0 15088 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_156
timestamp 1676037725
transform 1 0 15456 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_166
timestamp 1676037725
transform 1 0 16376 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_185
timestamp 1676037725
transform 1 0 18124 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_195
timestamp 1676037725
transform 1 0 19044 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_212
timestamp 1676037725
transform 1 0 20608 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_218
timestamp 1676037725
transform 1 0 21160 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_229
timestamp 1676037725
transform 1 0 22172 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_232
timestamp 1676037725
transform 1 0 22448 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_240
timestamp 1676037725
transform 1 0 23184 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1676037725
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_75
timestamp 1676037725
transform 1 0 8004 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_79
timestamp 1676037725
transform 1 0 8372 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_105
timestamp 1676037725
transform 1 0 10764 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_134
timestamp 1676037725
transform 1 0 13432 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_138
timestamp 1676037725
transform 1 0 13800 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_162
timestamp 1676037725
transform 1 0 16008 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_168
timestamp 1676037725
transform 1 0 16560 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_178
timestamp 1676037725
transform 1 0 17480 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_190
timestamp 1676037725
transform 1 0 18584 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_205
timestamp 1676037725
transform 1 0 19964 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_210
timestamp 1676037725
transform 1 0 20424 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_214
timestamp 1676037725
transform 1 0 20792 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_224
timestamp 1676037725
transform 1 0 21712 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_230
timestamp 1676037725
transform 1 0 22264 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_241
timestamp 1676037725
transform 1 0 23276 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_247
timestamp 1676037725
transform 1 0 23828 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_259
timestamp 1676037725
transform 1 0 24932 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_264
timestamp 1676037725
transform 1 0 25392 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_8
timestamp 1676037725
transform 1 0 1840 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_12
timestamp 1676037725
transform 1 0 2208 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_20
timestamp 1676037725
transform 1 0 2944 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_26
timestamp 1676037725
transform 1 0 3496 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_30
timestamp 1676037725
transform 1 0 3864 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_42
timestamp 1676037725
transform 1 0 4968 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_54
timestamp 1676037725
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_109
timestamp 1676037725
transform 1 0 11132 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_124
timestamp 1676037725
transform 1 0 12512 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_156
timestamp 1676037725
transform 1 0 15456 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_160
timestamp 1676037725
transform 1 0 15824 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_191
timestamp 1676037725
transform 1 0 18676 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_197
timestamp 1676037725
transform 1 0 19228 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_208
timestamp 1676037725
transform 1 0 20240 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_212
timestamp 1676037725
transform 1 0 20608 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1676037725
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_230
timestamp 1676037725
transform 1 0 22264 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_236
timestamp 1676037725
transform 1 0 22816 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_257
timestamp 1676037725
transform 1 0 24748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1676037725
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1676037725
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_46
timestamp 1676037725
transform 1 0 5336 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_50
timestamp 1676037725
transform 1 0 5704 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_72
timestamp 1676037725
transform 1 0 7728 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_76
timestamp 1676037725
transform 1 0 8096 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_100
timestamp 1676037725
transform 1 0 10304 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_113
timestamp 1676037725
transform 1 0 11500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_117
timestamp 1676037725
transform 1 0 11868 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_129
timestamp 1676037725
transform 1 0 12972 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13432 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_161
timestamp 1676037725
transform 1 0 15916 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_173
timestamp 1676037725
transform 1 0 17020 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 1676037725
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_219
timestamp 1676037725
transform 1 0 21252 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_232
timestamp 1676037725
transform 1 0 22448 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1676037725
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1676037725
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_259
timestamp 1676037725
transform 1 0 24932 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1676037725
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_31
timestamp 1676037725
transform 1 0 3956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_37
timestamp 1676037725
transform 1 0 4508 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_45
timestamp 1676037725
transform 1 0 5244 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_49
timestamp 1676037725
transform 1 0 5612 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1676037725
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_63
timestamp 1676037725
transform 1 0 6900 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_67
timestamp 1676037725
transform 1 0 7268 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_89
timestamp 1676037725
transform 1 0 9292 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_102
timestamp 1676037725
transform 1 0 10488 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_106
timestamp 1676037725
transform 1 0 10856 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_138
timestamp 1676037725
transform 1 0 13800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_145
timestamp 1676037725
transform 1 0 14444 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_153
timestamp 1676037725
transform 1 0 15180 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_164
timestamp 1676037725
transform 1 0 16192 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_180
timestamp 1676037725
transform 1 0 17664 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_188
timestamp 1676037725
transform 1 0 18400 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_191
timestamp 1676037725
transform 1 0 18676 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_204
timestamp 1676037725
transform 1 0 19872 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_217
timestamp 1676037725
transform 1 0 21068 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_221
timestamp 1676037725
transform 1 0 21436 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_238
timestamp 1676037725
transform 1 0 23000 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_242
timestamp 1676037725
transform 1 0 23368 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_263
timestamp 1676037725
transform 1 0 25300 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_37
timestamp 1676037725
transform 1 0 4508 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_43
timestamp 1676037725
transform 1 0 5060 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_47
timestamp 1676037725
transform 1 0 5428 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_59
timestamp 1676037725
transform 1 0 6532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_71
timestamp 1676037725
transform 1 0 7636 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_79
timestamp 1676037725
transform 1 0 8372 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_87
timestamp 1676037725
transform 1 0 9108 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_91
timestamp 1676037725
transform 1 0 9476 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_101
timestamp 1676037725
transform 1 0 10396 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_125
timestamp 1676037725
transform 1 0 12604 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_129
timestamp 1676037725
transform 1 0 12972 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_137
timestamp 1676037725
transform 1 0 13708 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_145
timestamp 1676037725
transform 1 0 14444 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_169
timestamp 1676037725
transform 1 0 16652 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_173
timestamp 1676037725
transform 1 0 17020 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_183
timestamp 1676037725
transform 1 0 17940 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_187
timestamp 1676037725
transform 1 0 18308 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_191
timestamp 1676037725
transform 1 0 18676 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_220
timestamp 1676037725
transform 1 0 21344 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_224
timestamp 1676037725
transform 1 0 21712 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_234
timestamp 1676037725
transform 1 0 22632 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1676037725
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_255
timestamp 1676037725
transform 1 0 24564 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_265
timestamp 1676037725
transform 1 0 25484 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_9
timestamp 1676037725
transform 1 0 1932 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_13
timestamp 1676037725
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_25
timestamp 1676037725
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_37
timestamp 1676037725
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1676037725
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_75
timestamp 1676037725
transform 1 0 8004 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_83
timestamp 1676037725
transform 1 0 8740 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_96
timestamp 1676037725
transform 1 0 9936 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_100
timestamp 1676037725
transform 1 0 10304 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_110
timestamp 1676037725
transform 1 0 8280 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_102
timestamp 1676037725
transform 1 0 10488 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_106
timestamp 1676037725
transform 1 0 10856 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_121
timestamp 1676037725
transform 1 0 12236 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_143
timestamp 1676037725
transform 1 0 14260 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_156
timestamp 1676037725
transform 1 0 15456 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_160
timestamp 1676037725
transform 1 0 15824 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_171
timestamp 1676037725
transform 1 0 16836 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_182
timestamp 1676037725
transform 1 0 17848 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_186
timestamp 1676037725
transform 1 0 18216 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_207
timestamp 1676037725
transform 1 0 20148 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_211
timestamp 1676037725
transform 1 0 20516 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_219
timestamp 1676037725
transform 1 0 21252 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_236
timestamp 1676037725
transform 1 0 22816 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1676037725
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_8
timestamp 1676037725
transform 1 0 1840 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_12
timestamp 1676037725
transform 1 0 2208 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_24
timestamp 1676037725
transform 1 0 3312 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_59
timestamp 1676037725
transform 1 0 6532 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_64
timestamp 1676037725
transform 1 0 6992 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_68
timestamp 1676037725
transform 1 0 7360 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_76
timestamp 1676037725
transform 1 0 8096 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_82
timestamp 1676037725
transform 1 0 8648 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_108
timestamp 1676037725
transform 1 0 11040 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_116
timestamp 1676037725
transform 1 0 11776 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_120
timestamp 1676037725
transform 1 0 12144 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_132
timestamp 1676037725
transform 1 0 13248 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14260 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_181
timestamp 1676037725
transform 1 0 17756 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_184
timestamp 1676037725
transform 1 0 18032 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_221
timestamp 1676037725
transform 1 0 21436 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_225
timestamp 1676037725
transform 1 0 21804 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_236
timestamp 1676037725
transform 1 0 22816 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_248
timestamp 1676037725
transform 1 0 23920 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_261
timestamp 1676037725
transform 1 0 25116 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_54
timestamp 1676037725
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_63
timestamp 1676037725
transform 1 0 6900 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_71
timestamp 1676037725
transform 1 0 7636 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_78
timestamp 1676037725
transform 1 0 8280 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_88
timestamp 1676037725
transform 1 0 9200 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_92
timestamp 1676037725
transform 1 0 9568 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_104
timestamp 1676037725
transform 1 0 10672 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_110
timestamp 1676037725
transform 1 0 11224 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_115
timestamp 1676037725
transform 1 0 11684 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_126
timestamp 1676037725
transform 1 0 12696 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_130
timestamp 1676037725
transform 1 0 13064 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_151
timestamp 1676037725
transform 1 0 14996 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_155
timestamp 1676037725
transform 1 0 15364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_191
timestamp 1676037725
transform 1 0 18676 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_195
timestamp 1676037725
transform 1 0 19044 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_199
timestamp 1676037725
transform 1 0 19412 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_220
timestamp 1676037725
transform 1 0 21344 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_229
timestamp 1676037725
transform 1 0 22172 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_250
timestamp 1676037725
transform 1 0 24104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1676037725
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1676037725
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_59
timestamp 1676037725
transform 1 0 6532 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_67
timestamp 1676037725
transform 1 0 7268 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_75
timestamp 1676037725
transform 1 0 8004 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_79
timestamp 1676037725
transform 1 0 8372 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_91
timestamp 1676037725
transform 1 0 9476 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_95
timestamp 1676037725
transform 1 0 9844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_107
timestamp 1676037725
transform 1 0 10948 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_110
timestamp 1676037725
transform 1 0 11224 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_116
timestamp 1676037725
transform 1 0 11776 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_120
timestamp 1676037725
transform 1 0 12144 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_125
timestamp 1676037725
transform 1 0 12604 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_138
timestamp 1676037725
transform 1 0 13800 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_149
timestamp 1676037725
transform 1 0 14812 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_172
timestamp 1676037725
transform 1 0 16928 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_176
timestamp 1676037725
transform 1 0 17296 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_188
timestamp 1676037725
transform 1 0 18400 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_220
timestamp 1676037725
transform 1 0 21344 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_224
timestamp 1676037725
transform 1 0 21712 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_250
timestamp 1676037725
transform 1 0 24104 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_255
timestamp 1676037725
transform 1 0 24564 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_263
timestamp 1676037725
transform 1 0 25300 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_5
timestamp 1676037725
transform 1 0 1564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_17
timestamp 1676037725
transform 1 0 2668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_29
timestamp 1676037725
transform 1 0 3772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_41
timestamp 1676037725
transform 1 0 4876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_53
timestamp 1676037725
transform 1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_86
timestamp 1676037725
transform 1 0 9016 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_108
timestamp 1676037725
transform 1 0 11040 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_121
timestamp 1676037725
transform 1 0 12236 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_133
timestamp 1676037725
transform 1 0 13340 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_141
timestamp 1676037725
transform 1 0 14076 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_164
timestamp 1676037725
transform 1 0 16192 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_187
timestamp 1676037725
transform 1 0 18308 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_208
timestamp 1676037725
transform 1 0 20240 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_212
timestamp 1676037725
transform 1 0 20608 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_215
timestamp 1676037725
transform 1 0 20884 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_247
timestamp 1676037725
transform 1 0 23828 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_251
timestamp 1676037725
transform 1 0 24196 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_264
timestamp 1676037725
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1676037725
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_73
timestamp 1676037725
transform 1 0 7820 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_78
timestamp 1676037725
transform 1 0 8280 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1676037725
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_90
timestamp 1676037725
transform 1 0 9384 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_96
timestamp 1676037725
transform 1 0 9936 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_100
timestamp 1676037725
transform 1 0 10304 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_113
timestamp 1676037725
transform 1 0 11500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_138
timestamp 1676037725
transform 1 0 13800 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_143
timestamp 1676037725
transform 1 0 14260 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_155
timestamp 1676037725
transform 1 0 15364 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_163
timestamp 1676037725
transform 1 0 16100 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_168
timestamp 1676037725
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_180
timestamp 1676037725
transform 1 0 17664 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_188
timestamp 1676037725
transform 1 0 18400 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_193
timestamp 1676037725
transform 1 0 18860 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_200
timestamp 1676037725
transform 1 0 19504 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_211
timestamp 1676037725
transform 1 0 20516 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_224
timestamp 1676037725
transform 1 0 21712 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_236
timestamp 1676037725
transform 1 0 22816 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_250
timestamp 1676037725
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_255
timestamp 1676037725
transform 1 0 24564 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_263
timestamp 1676037725
transform 1 0 25300 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_65
timestamp 1676037725
transform 1 0 7084 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_109
timestamp 1676037725
transform 1 0 11132 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_121
timestamp 1676037725
transform 1 0 12236 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_142
timestamp 1676037725
transform 1 0 14168 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1676037725
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_191
timestamp 1676037725
transform 1 0 18676 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_215
timestamp 1676037725
transform 1 0 20884 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_219
timestamp 1676037725
transform 1 0 21252 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 20424 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_228
timestamp 1676037725
transform 1 0 22080 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_239
timestamp 1676037725
transform 1 0 23092 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_251
timestamp 1676037725
transform 1 0 24196 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1676037725
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_119
timestamp 1676037725
transform 1 0 12052 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_123
timestamp 1676037725
transform 1 0 12420 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1676037725
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1676037725
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_144
timestamp 1676037725
transform 1 0 14352 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_156
timestamp 1676037725
transform 1 0 15456 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_178
timestamp 1676037725
transform 1 0 17480 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_182
timestamp 1676037725
transform 1 0 17848 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1676037725
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_199
timestamp 1676037725
transform 1 0 19412 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_211
timestamp 1676037725
transform 1 0 20516 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_225
timestamp 1676037725
transform 1 0 21804 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_236
timestamp 1676037725
transform 1 0 22816 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_248
timestamp 1676037725
transform 1 0 23920 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_259
timestamp 1676037725
transform 1 0 24932 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_264
timestamp 1676037725
transform 1 0 25392 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1676037725
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1676037725
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1676037725
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1676037725
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1676037725
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_90
timestamp 1676037725
transform 1 0 9384 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_102
timestamp 1676037725
transform 1 0 10488 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_110
timestamp 1676037725
transform 1 0 11224 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_180
timestamp 1676037725
transform 1 0 17664 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_197
timestamp 1676037725
transform 1 0 19228 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_209
timestamp 1676037725
transform 1 0 20332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_221
timestamp 1676037725
transform 1 0 21436 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_253
timestamp 1676037725
transform 1 0 24380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1676037725
transform 1 0 24932 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_263
timestamp 1676037725
transform 1 0 25300 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_9
timestamp 1676037725
transform 1 0 1932 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_13
timestamp 1676037725
transform 1 0 2300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_25
timestamp 1676037725
transform 1 0 3404 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1676037725
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_182
timestamp 1676037725
transform 1 0 17848 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_194
timestamp 1676037725
transform 1 0 18952 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_241
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_259
timestamp 1676037725
transform 1 0 24932 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1676037725
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1676037725
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_129
timestamp 1676037725
transform 1 0 12972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_141
timestamp 1676037725
transform 1 0 14076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_153
timestamp 1676037725
transform 1 0 15180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_165
timestamp 1676037725
transform 1 0 16284 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1676037725
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_35
timestamp 1676037725
transform 1 0 4324 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_86_59
timestamp 1676037725
transform 1 0 6532 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_63
timestamp 1676037725
transform 1 0 6900 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_75
timestamp 1676037725
transform 1 0 8004 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_113
timestamp 1676037725
transform 1 0 11500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_117
timestamp 1676037725
transform 1 0 11868 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_129
timestamp 1676037725
transform 1 0 12972 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_137
timestamp 1676037725
transform 1 0 13708 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_259
timestamp 1676037725
transform 1 0 24932 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1676037725
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_87_25
timestamp 1676037725
transform 1 0 3404 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_87_54
timestamp 1676037725
transform 1 0 6072 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_59
timestamp 1676037725
transform 1 0 6532 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_71
timestamp 1676037725
transform 1 0 7636 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_83
timestamp 1676037725
transform 1 0 8740 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_90
timestamp 1676037725
transform 1 0 9384 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_102
timestamp 1676037725
transform 1 0 10488 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_110
timestamp 1676037725
transform 1 0 11224 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1676037725
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_88_3
timestamp 1676037725
transform 1 0 24840 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1676037725
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_5
timestamp 1676037725
transform 1 0 1564 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_9
timestamp 1676037725
transform 1 0 1932 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1676037725
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_45
timestamp 1676037725
transform 1 0 5244 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_57
timestamp 1676037725
transform 1 0 6348 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_61
timestamp 1676037725
transform 1 0 6716 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1676037725
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1676037725
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_91
timestamp 1676037725
transform 1 0 9476 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_103
timestamp 1676037725
transform 1 0 10580 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_115
timestamp 1676037725
transform 1 0 11684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_127
timestamp 1676037725
transform 1 0 12788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1676037725
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_261
timestamp 1676037725
transform 1 0 25116 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_11
timestamp 1676037725
transform 1 0 2116 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_29
timestamp 1676037725
transform 1 0 3772 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_49
timestamp 1676037725
transform 1 0 5612 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1676037725
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_65
timestamp 1676037725
transform 1 0 7084 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_79
timestamp 1676037725
transform 1 0 8372 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_87
timestamp 1676037725
transform 1 0 9108 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_255
timestamp 1676037725
transform 1 0 24564 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_258
timestamp 1676037725
transform 1 0 24840 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1676037725
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_9
timestamp 1676037725
transform 1 0 1932 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_26
timestamp 1676037725
transform 1 0 3496 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_31
timestamp 1676037725
transform 1 0 3956 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_43
timestamp 1676037725
transform 1 0 5060 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_61
timestamp 1676037725
transform 1 0 6716 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1676037725
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_97
timestamp 1676037725
transform 1 0 10028 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_102
timestamp 1676037725
transform 1 0 10488 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_114
timestamp 1676037725
transform 1 0 11592 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_126
timestamp 1676037725
transform 1 0 12696 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_138
timestamp 1676037725
transform 1 0 13800 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_250
timestamp 1676037725
transform 1 0 24104 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_255
timestamp 1676037725
transform 1 0 24564 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_258
timestamp 1676037725
transform 1 0 24840 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1676037725
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_15
timestamp 1676037725
transform 1 0 2484 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_34
timestamp 1676037725
transform 1 0 4232 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_54
timestamp 1676037725
transform 1 0 6072 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_61
timestamp 1676037725
transform 1 0 6716 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_66
timestamp 1676037725
transform 1 0 7176 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_72
timestamp 1676037725
transform 1 0 7728 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_89
timestamp 1676037725
transform 1 0 9292 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_91_109
timestamp 1676037725
transform 1 0 11132 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_118
timestamp 1676037725
transform 1 0 11960 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_133
timestamp 1676037725
transform 1 0 13340 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_145
timestamp 1676037725
transform 1 0 14444 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_157
timestamp 1676037725
transform 1 0 15548 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_165
timestamp 1676037725
transform 1 0 16284 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_261
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_9
timestamp 1676037725
transform 1 0 1932 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_26
timestamp 1676037725
transform 1 0 3496 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_45
timestamp 1676037725
transform 1 0 5244 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_62
timestamp 1676037725
transform 1 0 6808 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1676037725
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_97
timestamp 1676037725
transform 1 0 10028 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_92_121
timestamp 1676037725
transform 1 0 12236 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_128
timestamp 1676037725
transform 1 0 12880 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_132
timestamp 1676037725
transform 1 0 13248 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_92_137
timestamp 1676037725
transform 1 0 13708 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_143
timestamp 1676037725
transform 1 0 14260 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_155
timestamp 1676037725
transform 1 0 15364 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_167
timestamp 1676037725
transform 1 0 16468 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_179
timestamp 1676037725
transform 1 0 17572 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_191
timestamp 1676037725
transform 1 0 18676 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_227
timestamp 1676037725
transform 1 0 21988 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_258
timestamp 1676037725
transform 1 0 24840 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1676037725
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_8
timestamp 1676037725
transform 1 0 1840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_12
timestamp 1676037725
transform 1 0 2208 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_34
timestamp 1676037725
transform 1 0 4232 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1676037725
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_73
timestamp 1676037725
transform 1 0 7820 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_90
timestamp 1676037725
transform 1 0 9384 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1676037725
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_133
timestamp 1676037725
transform 1 0 13340 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_141
timestamp 1676037725
transform 1 0 14076 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_148
timestamp 1676037725
transform 1 0 14720 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_152
timestamp 1676037725
transform 1 0 15088 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_160
timestamp 1676037725
transform 1 0 15824 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_164
timestamp 1676037725
transform 1 0 16192 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_177
timestamp 1676037725
transform 1 0 17388 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_189
timestamp 1676037725
transform 1 0 18492 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_196
timestamp 1676037725
transform 1 0 19136 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_204
timestamp 1676037725
transform 1 0 19872 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_208
timestamp 1676037725
transform 1 0 20240 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_212
timestamp 1676037725
transform 1 0 20608 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_220
timestamp 1676037725
transform 1 0 21344 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_93_227
timestamp 1676037725
transform 1 0 21988 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_93_232
timestamp 1676037725
transform 1 0 22448 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_235
timestamp 1676037725
transform 1 0 22724 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_239
timestamp 1676037725
transform 1 0 23092 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_244
timestamp 1676037725
transform 1 0 23552 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_251
timestamp 1676037725
transform 1 0 24196 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_255
timestamp 1676037725
transform 1 0 24564 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_258
timestamp 1676037725
transform 1 0 24840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_242
timestamp 1676037725
transform 1 0 23368 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_93_264
timestamp 1676037725
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_9
timestamp 1676037725
transform 1 0 1932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1676037725
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_31
timestamp 1676037725
transform 1 0 3956 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_43
timestamp 1676037725
transform 1 0 5060 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_62
timestamp 1676037725
transform 1 0 6808 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_82
timestamp 1676037725
transform 1 0 8648 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_117
timestamp 1676037725
transform 1 0 11868 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_94_137
timestamp 1676037725
transform 1 0 13708 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_147
timestamp 1676037725
transform 1 0 14628 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_151
timestamp 1676037725
transform 1 0 14996 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_94_161
timestamp 1676037725
transform 1 0 15916 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_167
timestamp 1676037725
transform 1 0 16468 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_173
timestamp 1676037725
transform 1 0 17020 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_180
timestamp 1676037725
transform 1 0 17664 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_184
timestamp 1676037725
transform 1 0 18032 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_189
timestamp 1676037725
transform 1 0 18492 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1676037725
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_203
timestamp 1676037725
transform 1 0 19780 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_211
timestamp 1676037725
transform 1 0 20516 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_215
timestamp 1676037725
transform 1 0 20884 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_228
timestamp 1676037725
transform 1 0 22080 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_235
timestamp 1676037725
transform 1 0 22724 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_242
timestamp 1676037725
transform 1 0 23368 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1676037725
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_94_257
timestamp 1676037725
transform 1 0 24748 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_264
timestamp 1676037725
transform 1 0 25392 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1676037725
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1676037725
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_118
timestamp 1676037725
transform 1 0 11960 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_138
timestamp 1676037725
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_143
timestamp 1676037725
transform 1 0 14260 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_147
timestamp 1676037725
transform 1 0 14628 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_153
timestamp 1676037725
transform 1 0 15180 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_161
timestamp 1676037725
transform 1 0 15916 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_165
timestamp 1676037725
transform 1 0 16284 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_175
timestamp 1676037725
transform 1 0 17204 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_183
timestamp 1676037725
transform 1 0 17940 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_191
timestamp 1676037725
transform 1 0 18676 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_195
timestamp 1676037725
transform 1 0 19044 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_203
timestamp 1676037725
transform 1 0 19780 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_211
timestamp 1676037725
transform 1 0 20516 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_219
timestamp 1676037725
transform 1 0 21252 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1676037725
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_231
timestamp 1676037725
transform 1 0 22356 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_239
timestamp 1676037725
transform 1 0 23092 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_243
timestamp 1676037725
transform 1 0 23460 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1676037725
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_255
timestamp 1676037725
transform 1 0 24564 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_264
timestamp 1676037725
transform 1 0 25392 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform -1 0 1840 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 25116 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 25116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 25116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 25116 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 25116 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 24472 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 25116 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 25116 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform 1 0 23184 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1676037725
transform 1 0 24472 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1676037725
transform 1 0 24472 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 24472 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1676037725
transform 1 0 23184 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1676037725
transform 1 0 24472 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1676037725
transform 1 0 25116 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 25116 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 25116 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 23920 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 23828 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 25116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 25116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1676037725
transform 1 0 25116 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1676037725
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1676037725
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 7636 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1676037725
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1676037725
transform 1 0 7544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1676037725
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1676037725
transform 1 0 9016 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1676037725
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1676037725
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1676037725
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1676037725
transform 1 0 10304 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1676037725
transform 1 0 10948 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 11684 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1676037725
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1676037725
transform 1 0 3220 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1676037725
transform 1 0 2392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1676037725
transform 1 0 4692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1676037725
transform 1 0 5060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 11684 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1676037725
transform 1 0 16652 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1676037725
transform 1 0 17572 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 17388 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 18308 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 18124 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1676037725
transform 1 0 19412 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 19412 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1676037725
transform 1 0 20148 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1676037725
transform 1 0 20148 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1676037725
transform 1 0 13340 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1676037725
transform 1 0 20332 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 20884 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 21068 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 21988 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1676037725
transform 1 0 21804 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1676037725
transform 1 0 22448 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input81
timestamp 1676037725
transform 1 0 22724 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1676037725
transform 1 0 23092 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 23276 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 23920 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1676037725
transform 1 0 13708 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1676037725
transform 1 0 14260 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform 1 0 14444 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input88
timestamp 1676037725
transform 1 0 14812 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input89
timestamp 1676037725
transform 1 0 15548 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1676037725
transform 1 0 15548 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform 1 0 15916 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1676037725
transform 1 0 16836 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 1564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform 1 0 1564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform 1 0 1564 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform 1 0 1564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1676037725
transform 1 0 1564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input98
timestamp 1676037725
transform -1 0 25392 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1676037725
transform 1 0 25024 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input100
timestamp 1676037725
transform 1 0 25024 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1676037725
transform 1 0 25024 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1676037725
transform 1 0 25024 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input103 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24840 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1676037725
transform 1 0 25024 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input105
timestamp 1676037725
transform 1 0 23736 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1676037725
transform 1 0 23736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input107
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1676037725
transform 1 0 1564 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input109
timestamp 1676037725
transform 1 0 3956 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input110
timestamp 1676037725
transform 1 0 3956 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__conb_1  left_tile_210
timestamp 1676037725
transform 1 0 25116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output111 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18216 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 1564 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 22632 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 23920 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 23920 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 23920 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 20056 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 22080 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 23920 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 23920 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 22632 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 22080 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 23920 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 22632 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 23920 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 17572 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1676037725
transform 1 0 19412 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1676037725
transform 1 0 21252 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1676037725
transform 1 0 12420 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1676037725
transform 1 0 20516 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1676037725
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1676037725
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1676037725
transform 1 0 22356 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1676037725
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1676037725
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1676037725
transform 1 0 20792 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1676037725
transform 1 0 17480 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1676037725
transform 1 0 13524 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1676037725
transform 1 0 14260 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1676037725
transform 1 0 14628 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1676037725
transform 1 0 14996 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1676037725
transform 1 0 16836 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1676037725
transform 1 0 1932 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1676037725
transform 1 0 2024 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1676037725
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1676037725
transform 1 0 4600 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1676037725
transform 1 0 5336 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1676037725
transform 1 0 5336 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1676037725
transform 1 0 7176 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1676037725
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1676037725
transform 1 0 7820 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1676037725
transform 1 0 7176 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1676037725
transform 1 0 2024 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1676037725
transform 1 0 7912 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1676037725
transform 1 0 9660 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1676037725
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1676037725
transform 1 0 9752 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1676037725
transform 1 0 10764 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1676037725
transform 1 0 10396 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1676037725
transform 1 0 9752 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1676037725
transform 1 0 11868 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1676037725
transform 1 0 12328 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1676037725
transform 1 0 2300 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1676037725
transform 1 0 2024 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1676037725
transform 1 0 2760 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1676037725
transform 1 0 2024 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1676037725
transform 1 0 4140 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1676037725
transform 1 0 2760 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1676037725
transform 1 0 4600 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1676037725
transform 1 0 5244 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1676037725
transform 1 0 1564 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1676037725
transform 1 0 1564 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1676037725
transform 1 0 1564 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16192 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16468 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19872 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18768 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15364 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 15916 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17572 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20608 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21896 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22816 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16192 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14444 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14076 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 12880 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15916 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18032 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15364 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17572 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22172 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 25300 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23460 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22908 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23552 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23460 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22080 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22264 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22816 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform -1 0 25392 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23460 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22264 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19504 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19504 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19504 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18308 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18400 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19044 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 16836 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15640 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 15088 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14352 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 13616 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12880 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12052 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 11684 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10396 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9568 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10580 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12512 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12696 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9936 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8280 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7728 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6532 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6164 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6532 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6440 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6808 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7636 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11500 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15364 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15916 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19872 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21712 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20884 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform -1 0 21528 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18216 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3956 0 -1 50048
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9200 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 10212 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11868 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13156 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 12328 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12328 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10948 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 8924 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8464 0 -1 40256
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6808 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 5428 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6532 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 5520 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 4232 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6532 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6164 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 5244 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7544 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9384 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 8832 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8096 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6072 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 3956 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6164 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 5888 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10764 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14812 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 15916 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18032 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 11960 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15364 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1__260
timestamp 1676037725
transform 1 0 13892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 13524 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19044 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1__211
timestamp 1676037725
transform 1 0 17664 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17204 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1__226
timestamp 1676037725
transform -1 0 16928 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18952 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19596 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20240 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1__214
timestamp 1676037725
transform 1 0 21988 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17848 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20608 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18032 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3__216
timestamp 1676037725
transform 1 0 17020 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3_
timestamp 1676037725
transform 1 0 16836 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18032 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17112 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_2_
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3_
timestamp 1676037725
transform 1 0 13432 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3__261
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17204 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14720 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17572 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20700 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_2_
timestamp 1676037725
transform 1 0 17572 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19596 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1__262
timestamp 1676037725
transform 1 0 20700 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19504 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19872 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20056 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21528 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1__263
timestamp 1676037725
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22080 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23184 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16100 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19964 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18124 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1__264
timestamp 1676037725
transform 1 0 16928 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15640 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15548 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17940 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19780 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12788 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1__212
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l3_in_0_
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13064 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20332 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20792 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1_
timestamp 1676037725
transform 1 0 21068 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1__213
timestamp 1676037725
transform 1 0 22632 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18308 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1__215
timestamp 1676037725
transform 1 0 14352 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14996 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11224 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10396 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20976 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21896 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_0.mux_l2_in_1__217
timestamp 1676037725
transform 1 0 20884 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22908 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22264 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21252 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20240 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_2.mux_l2_in_1__223
timestamp 1676037725
transform 1 0 23828 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22632 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_2.mux_l2_in_1__238
timestamp 1676037725
transform 1 0 23368 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform -1 0 24840 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23184 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_4.mux_l2_in_1__234
timestamp 1676037725
transform 1 0 21988 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19780 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22264 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23644 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20240 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_6.mux_l2_in_1__243
timestamp 1676037725
transform 1 0 22448 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23184 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform -1 0 24104 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20884 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18952 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21804 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 21620 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_8.mux_l2_in_1__244
timestamp 1676037725
transform 1 0 21988 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22448 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20884 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19780 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20240 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_10.mux_l2_in_1__218
timestamp 1676037725
transform 1 0 17296 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 16100 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20608 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22172 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19688 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_12.mux_l2_in_1__219
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17020 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_14.mux_l2_in_1__220
timestamp 1676037725
transform 1 0 16836 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18216 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14352 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_16.mux_l2_in_1__221
timestamp 1676037725
transform 1 0 14260 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16652 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20056 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16192 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_18.mux_l2_in_1__222
timestamp 1676037725
transform 1 0 13524 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12880 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16100 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14628 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13340 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_20.mux_l2_in_1__224
timestamp 1676037725
transform 1 0 13156 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11960 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12604 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_22.mux_l2_in_1__225
timestamp 1676037725
transform 1 0 11684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12604 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17572 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15088 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12604 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_24.mux_l1_in_1__226
timestamp 1676037725
transform 1 0 13156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_26.mux_l1_in_1__227
timestamp 1676037725
transform 1 0 11960 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_1_
timestamp 1676037725
transform 1 0 11408 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14720 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 9200 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_28.mux_l1_in_1__228
timestamp 1676037725
transform 1 0 9384 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12144 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_1_
timestamp 1676037725
transform 1 0 8740 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_30.mux_l1_in_1__229
timestamp 1676037725
transform 1 0 8648 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16008 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11408 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_32.mux_l1_in_1__230
timestamp 1676037725
transform 1 0 8004 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_1_
timestamp 1676037725
transform 1 0 7636 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15456 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_34.mux_l1_in_1__231
timestamp 1676037725
transform 1 0 10028 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_1_
timestamp 1676037725
transform 1 0 8832 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10764 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11408 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_36.mux_l2_in_1__232
timestamp 1676037725
transform -1 0 6072 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_1_
timestamp 1676037725
transform -1 0 7360 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 8188 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14628 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12236 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_38.mux_l2_in_0__233
timestamp 1676037725
transform 1 0 14720 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform -1 0 15088 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14168 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l2_in_0_
timestamp 1676037725
transform -1 0 17664 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_40.mux_l2_in_0__235
timestamp 1676037725
transform 1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16192 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_44.mux_l2_in_0__236
timestamp 1676037725
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18400 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20424 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17480 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20056 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_46.mux_l2_in_0__237
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_48.mux_l2_in_0__238
timestamp 1676037725
transform 1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23184 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_50.mux_l1_in_1__239
timestamp 1676037725
transform 1 0 20424 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19228 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23000 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform -1 0 20240 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_52.mux_l2_in_0__240
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21068 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22724 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17756 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_54.mux_l2_in_0__241
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21528 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17296 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_56.mux_l2_in_0__242
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9108 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17112 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14904 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 10028 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_0.mux_l1_in_3__245
timestamp 1676037725
transform 1 0 9384 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform -1 0 12512 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10672 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11592 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 12696 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15364 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_2.mux_l2_in_1__248
timestamp 1676037725
transform 1 0 14168 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_2.mux_l2_in_1__263
timestamp 1676037725
transform 1 0 12236 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12696 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_2_
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 10396 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_4.mux_l2_in_1__252
timestamp 1676037725
transform 1 0 11684 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10672 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9200 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14260 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_6.mux_l1_in_3__255
timestamp 1676037725
transform 1 0 9844 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_3_
timestamp 1676037725
transform 1 0 8648 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9752 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9292 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7268 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9108 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17296 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_2_
timestamp 1676037725
transform 1 0 12788 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_10.mux_l1_in_3__246
timestamp 1676037725
transform 1 0 7912 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9200 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9108 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8004 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 16376 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 7452 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_12.mux_l2_in_1__247
timestamp 1676037725
transform 1 0 6900 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7636 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7728 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14536 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18308 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_2_
timestamp 1676037725
transform 1 0 9476 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_20.mux_l2_in_1__249
timestamp 1676037725
transform 1 0 9752 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9384 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9016 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12328 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12880 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_28.mux_l2_in_1__250
timestamp 1676037725
transform 1 0 5336 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_1_
timestamp 1676037725
transform 1 0 4968 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l3_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11408 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11868 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_36.mux_l2_in_1__251
timestamp 1676037725
transform 1 0 9108 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_1_
timestamp 1676037725
transform -1 0 8648 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7176 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_44.mux_l1_in_1__253
timestamp 1676037725
transform 1 0 10948 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19136 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_52.mux_l2_in_1__254
timestamp 1676037725
transform 1 0 14444 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 55360 800 55480 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1490 56200 1546 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1674 0 1730 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 66 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 67 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 68 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 69 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 70 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 71 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 72 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 73 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 74 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 75 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 76 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 77 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 chany_bottom_in[20]
port 78 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 chany_bottom_in[21]
port 79 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 chany_bottom_in[22]
port 80 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_in[23]
port 81 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 chany_bottom_in[24]
port 82 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_in[25]
port 83 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 chany_bottom_in[26]
port 84 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 chany_bottom_in[27]
port 85 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 chany_bottom_in[28]
port 86 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 chany_bottom_in[29]
port 87 nsew signal input
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 88 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 89 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 90 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 91 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 92 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 93 nsew signal input
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 94 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 95 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 96 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 97 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 98 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 99 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 100 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 101 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 102 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 103 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 104 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 105 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 106 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 107 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 chany_bottom_out[20]
port 108 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 chany_bottom_out[21]
port 109 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 chany_bottom_out[22]
port 110 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 chany_bottom_out[23]
port 111 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 chany_bottom_out[24]
port 112 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 chany_bottom_out[25]
port 113 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 chany_bottom_out[26]
port 114 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 chany_bottom_out[27]
port 115 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 chany_bottom_out[28]
port 116 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 chany_bottom_out[29]
port 117 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 118 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 119 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 120 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 121 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 122 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 123 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 124 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 125 nsew signal tristate
flabel metal2 s 12898 56200 12954 57000 0 FreeSans 224 90 0 0 chany_top_in_0[0]
port 126 nsew signal input
flabel metal2 s 16578 56200 16634 57000 0 FreeSans 224 90 0 0 chany_top_in_0[10]
port 127 nsew signal input
flabel metal2 s 16946 56200 17002 57000 0 FreeSans 224 90 0 0 chany_top_in_0[11]
port 128 nsew signal input
flabel metal2 s 17314 56200 17370 57000 0 FreeSans 224 90 0 0 chany_top_in_0[12]
port 129 nsew signal input
flabel metal2 s 17682 56200 17738 57000 0 FreeSans 224 90 0 0 chany_top_in_0[13]
port 130 nsew signal input
flabel metal2 s 18050 56200 18106 57000 0 FreeSans 224 90 0 0 chany_top_in_0[14]
port 131 nsew signal input
flabel metal2 s 18418 56200 18474 57000 0 FreeSans 224 90 0 0 chany_top_in_0[15]
port 132 nsew signal input
flabel metal2 s 18786 56200 18842 57000 0 FreeSans 224 90 0 0 chany_top_in_0[16]
port 133 nsew signal input
flabel metal2 s 19154 56200 19210 57000 0 FreeSans 224 90 0 0 chany_top_in_0[17]
port 134 nsew signal input
flabel metal2 s 19522 56200 19578 57000 0 FreeSans 224 90 0 0 chany_top_in_0[18]
port 135 nsew signal input
flabel metal2 s 19890 56200 19946 57000 0 FreeSans 224 90 0 0 chany_top_in_0[19]
port 136 nsew signal input
flabel metal2 s 13266 56200 13322 57000 0 FreeSans 224 90 0 0 chany_top_in_0[1]
port 137 nsew signal input
flabel metal2 s 20258 56200 20314 57000 0 FreeSans 224 90 0 0 chany_top_in_0[20]
port 138 nsew signal input
flabel metal2 s 20626 56200 20682 57000 0 FreeSans 224 90 0 0 chany_top_in_0[21]
port 139 nsew signal input
flabel metal2 s 20994 56200 21050 57000 0 FreeSans 224 90 0 0 chany_top_in_0[22]
port 140 nsew signal input
flabel metal2 s 21362 56200 21418 57000 0 FreeSans 224 90 0 0 chany_top_in_0[23]
port 141 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 chany_top_in_0[24]
port 142 nsew signal input
flabel metal2 s 22098 56200 22154 57000 0 FreeSans 224 90 0 0 chany_top_in_0[25]
port 143 nsew signal input
flabel metal2 s 22466 56200 22522 57000 0 FreeSans 224 90 0 0 chany_top_in_0[26]
port 144 nsew signal input
flabel metal2 s 22834 56200 22890 57000 0 FreeSans 224 90 0 0 chany_top_in_0[27]
port 145 nsew signal input
flabel metal2 s 23202 56200 23258 57000 0 FreeSans 224 90 0 0 chany_top_in_0[28]
port 146 nsew signal input
flabel metal2 s 23570 56200 23626 57000 0 FreeSans 224 90 0 0 chany_top_in_0[29]
port 147 nsew signal input
flabel metal2 s 13634 56200 13690 57000 0 FreeSans 224 90 0 0 chany_top_in_0[2]
port 148 nsew signal input
flabel metal2 s 14002 56200 14058 57000 0 FreeSans 224 90 0 0 chany_top_in_0[3]
port 149 nsew signal input
flabel metal2 s 14370 56200 14426 57000 0 FreeSans 224 90 0 0 chany_top_in_0[4]
port 150 nsew signal input
flabel metal2 s 14738 56200 14794 57000 0 FreeSans 224 90 0 0 chany_top_in_0[5]
port 151 nsew signal input
flabel metal2 s 15106 56200 15162 57000 0 FreeSans 224 90 0 0 chany_top_in_0[6]
port 152 nsew signal input
flabel metal2 s 15474 56200 15530 57000 0 FreeSans 224 90 0 0 chany_top_in_0[7]
port 153 nsew signal input
flabel metal2 s 15842 56200 15898 57000 0 FreeSans 224 90 0 0 chany_top_in_0[8]
port 154 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 chany_top_in_0[9]
port 155 nsew signal input
flabel metal2 s 1858 56200 1914 57000 0 FreeSans 224 90 0 0 chany_top_out_0[0]
port 156 nsew signal tristate
flabel metal2 s 5538 56200 5594 57000 0 FreeSans 224 90 0 0 chany_top_out_0[10]
port 157 nsew signal tristate
flabel metal2 s 5906 56200 5962 57000 0 FreeSans 224 90 0 0 chany_top_out_0[11]
port 158 nsew signal tristate
flabel metal2 s 6274 56200 6330 57000 0 FreeSans 224 90 0 0 chany_top_out_0[12]
port 159 nsew signal tristate
flabel metal2 s 6642 56200 6698 57000 0 FreeSans 224 90 0 0 chany_top_out_0[13]
port 160 nsew signal tristate
flabel metal2 s 7010 56200 7066 57000 0 FreeSans 224 90 0 0 chany_top_out_0[14]
port 161 nsew signal tristate
flabel metal2 s 7378 56200 7434 57000 0 FreeSans 224 90 0 0 chany_top_out_0[15]
port 162 nsew signal tristate
flabel metal2 s 7746 56200 7802 57000 0 FreeSans 224 90 0 0 chany_top_out_0[16]
port 163 nsew signal tristate
flabel metal2 s 8114 56200 8170 57000 0 FreeSans 224 90 0 0 chany_top_out_0[17]
port 164 nsew signal tristate
flabel metal2 s 8482 56200 8538 57000 0 FreeSans 224 90 0 0 chany_top_out_0[18]
port 165 nsew signal tristate
flabel metal2 s 8850 56200 8906 57000 0 FreeSans 224 90 0 0 chany_top_out_0[19]
port 166 nsew signal tristate
flabel metal2 s 2226 56200 2282 57000 0 FreeSans 224 90 0 0 chany_top_out_0[1]
port 167 nsew signal tristate
flabel metal2 s 9218 56200 9274 57000 0 FreeSans 224 90 0 0 chany_top_out_0[20]
port 168 nsew signal tristate
flabel metal2 s 9586 56200 9642 57000 0 FreeSans 224 90 0 0 chany_top_out_0[21]
port 169 nsew signal tristate
flabel metal2 s 9954 56200 10010 57000 0 FreeSans 224 90 0 0 chany_top_out_0[22]
port 170 nsew signal tristate
flabel metal2 s 10322 56200 10378 57000 0 FreeSans 224 90 0 0 chany_top_out_0[23]
port 171 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 chany_top_out_0[24]
port 172 nsew signal tristate
flabel metal2 s 11058 56200 11114 57000 0 FreeSans 224 90 0 0 chany_top_out_0[25]
port 173 nsew signal tristate
flabel metal2 s 11426 56200 11482 57000 0 FreeSans 224 90 0 0 chany_top_out_0[26]
port 174 nsew signal tristate
flabel metal2 s 11794 56200 11850 57000 0 FreeSans 224 90 0 0 chany_top_out_0[27]
port 175 nsew signal tristate
flabel metal2 s 12162 56200 12218 57000 0 FreeSans 224 90 0 0 chany_top_out_0[28]
port 176 nsew signal tristate
flabel metal2 s 12530 56200 12586 57000 0 FreeSans 224 90 0 0 chany_top_out_0[29]
port 177 nsew signal tristate
flabel metal2 s 2594 56200 2650 57000 0 FreeSans 224 90 0 0 chany_top_out_0[2]
port 178 nsew signal tristate
flabel metal2 s 2962 56200 3018 57000 0 FreeSans 224 90 0 0 chany_top_out_0[3]
port 179 nsew signal tristate
flabel metal2 s 3330 56200 3386 57000 0 FreeSans 224 90 0 0 chany_top_out_0[4]
port 180 nsew signal tristate
flabel metal2 s 3698 56200 3754 57000 0 FreeSans 224 90 0 0 chany_top_out_0[5]
port 181 nsew signal tristate
flabel metal2 s 4066 56200 4122 57000 0 FreeSans 224 90 0 0 chany_top_out_0[6]
port 182 nsew signal tristate
flabel metal2 s 4434 56200 4490 57000 0 FreeSans 224 90 0 0 chany_top_out_0[7]
port 183 nsew signal tristate
flabel metal2 s 4802 56200 4858 57000 0 FreeSans 224 90 0 0 chany_top_out_0[8]
port 184 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 chany_top_out_0[9]
port 185 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal3 s 0 35776 800 35896 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal3 s 0 38224 800 38344 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal3 s 0 25984 800 26104 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal3 s 0 43120 800 43240 0 FreeSans 480 0 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 prog_reset
port 200 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 reset
port 201 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 202 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 203 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 204 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 205 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 206 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 207 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 208 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 209 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 210 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 211 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 212 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 213 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 test_enable
port 214 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal input
flabel metal3 s 0 48016 800 48136 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal input
flabel metal3 s 0 50464 800 50584 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal input
flabel metal3 s 0 52912 800 53032 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal2 6026 24276 6026 24276 0 cby_0__1_.cby_0__1_.ccff_tail
rlabel metal2 6210 25092 6210 25092 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 4508 23018 4508 23018 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 4232 19482 4232 19482 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 3450 20978 3450 20978 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 7498 19720 7498 19720 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 7636 7786 7636 7786 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 11684 18598 11684 18598 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal2 8326 20060 8326 20060 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal2 9430 16388 9430 16388 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 16192 12274 16192 12274 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 13570 18836 13570 18836 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 10810 14246 10810 14246 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 6900 17102 6900 17102 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal1 15410 12274 15410 12274 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal1 12788 15334 12788 15334 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal2 8418 16354 8418 16354 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 14536 19890 14536 19890 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal1 12098 21454 12098 21454 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 8878 21590 8878 21590 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal1 12926 14586 12926 14586 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7912 21658 7912 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 7084 21658 7084 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 14306 16830 14306 16830 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14030 18938 14030 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12742 23222 12742 23222 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11684 19482 11684 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11362 16218 11362 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 11730 20230 11730 20230 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 8786 20876 8786 20876 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 9200 21658 9200 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9476 20570 9476 20570 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15226 15334 15226 15334 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9798 17306 9798 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 8234 17850 8234 17850 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 14674 15946 14674 15946 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13478 20060 13478 20060 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13846 18394 13846 18394 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11454 21896 11454 21896 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 11730 16048 11730 16048 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11454 16558 11454 16558 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10350 16218 10350 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 11270 17306 11270 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10534 16456 10534 16456 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15042 13158 15042 13158 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7084 17578 7084 17578 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 6302 18598 6302 18598 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13616 13226 13616 13226 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14398 18734 14398 18734 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12742 17034 12742 17034 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9338 19482 9338 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 12374 14688 12374 14688 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10580 16150 10580 16150 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7912 17714 7912 17714 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 9154 16456 9154 16456 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8142 16218 8142 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 12190 16660 12190 16660 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 6256 22746 6256 22746 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 4784 22406 4784 22406 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 11914 18326 11914 18326 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14076 20026 14076 20026 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12052 21658 12052 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 10442 19584 10442 19584 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11638 18122 11638 18122 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10810 21658 10810 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7590 21114 7590 21114 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8004 22746 8004 22746 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8234 21386 8234 21386 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 4278 24956 4278 24956 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 3036 25806 3036 25806 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal2 3450 26894 3450 26894 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel via1 3795 28186 3795 28186 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 4324 20502 4324 20502 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 2254 20876 2254 20876 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 3036 23290 3036 23290 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 3565 27098 3565 27098 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 5796 20230 5796 20230 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal2 3634 20400 3634 20400 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 2254 23052 2254 23052 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 4071 25126 4071 25126 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 3542 20910 3542 20910 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 3036 21114 3036 21114 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 4301 23086 4301 23086 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal3 1740 55420 1740 55420 0 ccff_head
rlabel metal1 2484 3910 2484 3910 0 ccff_head_0
rlabel metal1 19274 6188 19274 6188 0 ccff_tail
rlabel metal1 1794 49266 1794 49266 0 ccff_tail_0
rlabel metal2 25346 24871 25346 24871 0 chanx_right_in[0]
rlabel via2 25346 34187 25346 34187 0 chanx_right_in[10]
rlabel via2 25346 35037 25346 35037 0 chanx_right_in[11]
rlabel metal1 25116 36142 25116 36142 0 chanx_right_in[12]
rlabel metal2 25346 36703 25346 36703 0 chanx_right_in[13]
rlabel metal2 25346 37349 25346 37349 0 chanx_right_in[14]
rlabel metal2 25346 38607 25346 38607 0 chanx_right_in[15]
rlabel metal1 24794 38930 24794 38930 0 chanx_right_in[16]
rlabel metal1 25070 40494 25070 40494 0 chanx_right_in[17]
rlabel metal2 25346 40919 25346 40919 0 chanx_right_in[18]
rlabel via2 25346 41565 25346 41565 0 chanx_right_in[19]
rlabel metal2 25530 26163 25530 26163 0 chanx_right_in[1]
rlabel metal1 24702 42534 24702 42534 0 chanx_right_in[20]
rlabel metal1 25438 43622 25438 43622 0 chanx_right_in[21]
rlabel metal2 25530 44353 25530 44353 0 chanx_right_in[22]
rlabel metal3 25584 44812 25584 44812 0 chanx_right_in[23]
rlabel metal1 24748 45798 24748 45798 0 chanx_right_in[24]
rlabel metal1 24840 46954 24840 46954 0 chanx_right_in[25]
rlabel metal1 25668 48518 25668 48518 0 chanx_right_in[26]
rlabel via2 25346 48093 25346 48093 0 chanx_right_in[27]
rlabel metal2 25346 49045 25346 49045 0 chanx_right_in[28]
rlabel metal2 25346 49759 25346 49759 0 chanx_right_in[29]
rlabel metal2 24150 28407 24150 28407 0 chanx_right_in[2]
rlabel metal1 24058 28492 24058 28492 0 chanx_right_in[3]
rlabel via2 25530 29291 25530 29291 0 chanx_right_in[4]
rlabel metal2 25346 29869 25346 29869 0 chanx_right_in[5]
rlabel metal2 25346 31127 25346 31127 0 chanx_right_in[6]
rlabel via2 25346 31773 25346 31773 0 chanx_right_in[7]
rlabel metal2 25346 32725 25346 32725 0 chanx_right_in[8]
rlabel metal1 24840 32538 24840 32538 0 chanx_right_in[9]
rlabel metal3 25676 9724 25676 9724 0 chanx_right_out[10]
rlabel metal2 24702 10013 24702 10013 0 chanx_right_out[11]
rlabel metal2 24794 10965 24794 10965 0 chanx_right_out[12]
rlabel metal2 25162 11985 25162 11985 0 chanx_right_out[13]
rlabel metal3 26044 12988 26044 12988 0 chanx_right_out[14]
rlabel metal2 24794 13277 24794 13277 0 chanx_right_out[15]
rlabel metal2 25162 14297 25162 14297 0 chanx_right_out[16]
rlabel metal3 25676 15436 25676 15436 0 chanx_right_out[17]
rlabel metal2 24702 15589 24702 15589 0 chanx_right_out[18]
rlabel metal3 25584 17068 25584 17068 0 chanx_right_out[19]
rlabel metal3 24296 2380 24296 2380 0 chanx_right_out[1]
rlabel metal1 23368 18190 23368 18190 0 chanx_right_out[20]
rlabel metal2 24702 17901 24702 17901 0 chanx_right_out[21]
rlabel metal2 24794 18853 24794 18853 0 chanx_right_out[22]
rlabel metal1 24426 19890 24426 19890 0 chanx_right_out[23]
rlabel metal1 23368 20502 23368 20502 0 chanx_right_out[24]
rlabel metal1 24380 20978 24380 20978 0 chanx_right_out[25]
rlabel metal1 23874 20366 23874 20366 0 chanx_right_out[26]
rlabel metal2 23874 23341 23874 23341 0 chanx_right_out[27]
rlabel metal1 24426 24242 24426 24242 0 chanx_right_out[28]
rlabel metal2 25162 25517 25162 25517 0 chanx_right_out[29]
rlabel metal2 22494 5236 22494 5236 0 chanx_right_out[2]
rlabel metal1 19228 5270 19228 5270 0 chanx_right_out[3]
rlabel metal3 24894 4828 24894 4828 0 chanx_right_out[4]
rlabel metal2 24794 5389 24794 5389 0 chanx_right_out[5]
rlabel metal3 25676 6460 25676 6460 0 chanx_right_out[6]
rlabel metal3 25768 7276 25768 7276 0 chanx_right_out[7]
rlabel metal2 25162 7769 25162 7769 0 chanx_right_out[8]
rlabel metal2 25162 8721 25162 8721 0 chanx_right_out[9]
rlabel metal1 1840 3502 1840 3502 0 chany_bottom_in[0]
rlabel metal1 5198 3026 5198 3026 0 chany_bottom_in[10]
rlabel metal1 5934 2346 5934 2346 0 chany_bottom_in[11]
rlabel metal2 6118 2132 6118 2132 0 chany_bottom_in[12]
rlabel metal2 6486 1792 6486 1792 0 chany_bottom_in[13]
rlabel metal2 6854 1894 6854 1894 0 chany_bottom_in[14]
rlabel metal2 7222 1588 7222 1588 0 chany_bottom_in[15]
rlabel metal1 7636 2414 7636 2414 0 chany_bottom_in[16]
rlabel metal1 7820 3366 7820 3366 0 chany_bottom_in[17]
rlabel metal1 7912 3026 7912 3026 0 chany_bottom_in[18]
rlabel metal2 8694 2064 8694 2064 0 chany_bottom_in[19]
rlabel metal1 1978 3026 1978 3026 0 chany_bottom_in[1]
rlabel metal2 9062 1860 9062 1860 0 chany_bottom_in[20]
rlabel metal1 9292 3502 9292 3502 0 chany_bottom_in[21]
rlabel metal1 9844 3502 9844 3502 0 chany_bottom_in[22]
rlabel metal1 9890 2414 9890 2414 0 chany_bottom_in[23]
rlabel metal1 10442 2958 10442 2958 0 chany_bottom_in[24]
rlabel metal1 10948 3502 10948 3502 0 chany_bottom_in[25]
rlabel metal1 11500 3026 11500 3026 0 chany_bottom_in[26]
rlabel metal1 11684 4046 11684 4046 0 chany_bottom_in[27]
rlabel metal1 11914 2448 11914 2448 0 chany_bottom_in[28]
rlabel metal1 10350 2380 10350 2380 0 chany_bottom_in[29]
rlabel metal1 2024 2414 2024 2414 0 chany_bottom_in[2]
rlabel metal1 2668 3026 2668 3026 0 chany_bottom_in[3]
rlabel metal1 3312 2958 3312 2958 0 chany_bottom_in[4]
rlabel metal1 2438 2380 2438 2380 0 chany_bottom_in[5]
rlabel metal1 3542 2414 3542 2414 0 chany_bottom_in[6]
rlabel metal1 4140 2414 4140 2414 0 chany_bottom_in[7]
rlabel metal1 4692 2414 4692 2414 0 chany_bottom_in[8]
rlabel metal1 4922 3366 4922 3366 0 chany_bottom_in[9]
rlabel metal2 12742 2166 12742 2166 0 chany_bottom_out[0]
rlabel metal2 16422 2404 16422 2404 0 chany_bottom_out[10]
rlabel metal2 16790 1792 16790 1792 0 chany_bottom_out[11]
rlabel metal2 17158 1826 17158 1826 0 chany_bottom_out[12]
rlabel metal2 17526 2404 17526 2404 0 chany_bottom_out[13]
rlabel metal2 17894 2166 17894 2166 0 chany_bottom_out[14]
rlabel metal2 18262 959 18262 959 0 chany_bottom_out[15]
rlabel metal2 18630 1928 18630 1928 0 chany_bottom_out[16]
rlabel metal2 18998 2098 18998 2098 0 chany_bottom_out[17]
rlabel metal2 19366 2948 19366 2948 0 chany_bottom_out[18]
rlabel metal2 19734 2676 19734 2676 0 chany_bottom_out[19]
rlabel metal2 13110 823 13110 823 0 chany_bottom_out[1]
rlabel metal2 20102 2404 20102 2404 0 chany_bottom_out[20]
rlabel metal2 20470 1775 20470 1775 0 chany_bottom_out[21]
rlabel metal2 20838 1792 20838 1792 0 chany_bottom_out[22]
rlabel metal2 21206 2370 21206 2370 0 chany_bottom_out[23]
rlabel metal2 21574 3254 21574 3254 0 chany_bottom_out[24]
rlabel metal2 21942 3492 21942 3492 0 chany_bottom_out[25]
rlabel metal1 22448 7310 22448 7310 0 chany_bottom_out[26]
rlabel metal2 22678 3560 22678 3560 0 chany_bottom_out[27]
rlabel metal2 23046 1639 23046 1639 0 chany_bottom_out[28]
rlabel metal2 23414 1826 23414 1826 0 chany_bottom_out[29]
rlabel metal2 13478 2370 13478 2370 0 chany_bottom_out[2]
rlabel metal2 13846 1554 13846 1554 0 chany_bottom_out[3]
rlabel metal2 14214 1860 14214 1860 0 chany_bottom_out[4]
rlabel metal2 14582 1622 14582 1622 0 chany_bottom_out[5]
rlabel metal2 14950 2166 14950 2166 0 chany_bottom_out[6]
rlabel metal2 15318 1622 15318 1622 0 chany_bottom_out[7]
rlabel metal2 15686 1860 15686 1860 0 chany_bottom_out[8]
rlabel metal2 16054 2166 16054 2166 0 chany_bottom_out[9]
rlabel metal1 11914 54196 11914 54196 0 chany_top_in_0[0]
rlabel metal1 16652 53550 16652 53550 0 chany_top_in_0[10]
rlabel metal1 17296 54162 17296 54162 0 chany_top_in_0[11]
rlabel metal1 17480 53550 17480 53550 0 chany_top_in_0[12]
rlabel metal1 18078 54230 18078 54230 0 chany_top_in_0[13]
rlabel metal2 18262 56236 18262 56236 0 chany_top_in_0[14]
rlabel metal1 19458 54128 19458 54128 0 chany_top_in_0[15]
rlabel metal1 18952 53074 18952 53074 0 chany_top_in_0[16]
rlabel metal1 19320 53550 19320 53550 0 chany_top_in_0[17]
rlabel metal1 19872 54162 19872 54162 0 chany_top_in_0[18]
rlabel metal1 20102 53550 20102 53550 0 chany_top_in_0[19]
rlabel metal2 13294 55711 13294 55711 0 chany_top_in_0[1]
rlabel metal1 20424 53074 20424 53074 0 chany_top_in_0[20]
rlabel metal2 20654 55711 20654 55711 0 chany_top_in_0[21]
rlabel metal1 21068 53550 21068 53550 0 chany_top_in_0[22]
rlabel metal1 21712 54162 21712 54162 0 chany_top_in_0[23]
rlabel metal1 21896 53550 21896 53550 0 chany_top_in_0[24]
rlabel metal1 22218 53210 22218 53210 0 chany_top_in_0[25]
rlabel metal1 22632 54162 22632 54162 0 chany_top_in_0[26]
rlabel metal1 23092 53550 23092 53550 0 chany_top_in_0[27]
rlabel metal2 23230 55711 23230 55711 0 chany_top_in_0[28]
rlabel metal1 23874 53074 23874 53074 0 chany_top_in_0[29]
rlabel metal1 13754 53142 13754 53142 0 chany_top_in_0[2]
rlabel metal1 14168 53550 14168 53550 0 chany_top_in_0[3]
rlabel metal1 14536 53074 14536 53074 0 chany_top_in_0[4]
rlabel metal1 14674 54298 14674 54298 0 chany_top_in_0[5]
rlabel metal1 15410 54162 15410 54162 0 chany_top_in_0[6]
rlabel metal1 15594 53550 15594 53550 0 chany_top_in_0[7]
rlabel metal1 16008 53074 16008 53074 0 chany_top_in_0[8]
rlabel metal1 16721 54162 16721 54162 0 chany_top_in_0[9]
rlabel metal1 2714 52870 2714 52870 0 chany_top_out_0[0]
rlabel metal1 5566 53652 5566 53652 0 chany_top_out_0[10]
rlabel metal1 4600 54094 4600 54094 0 chany_top_out_0[11]
rlabel metal1 6072 53142 6072 53142 0 chany_top_out_0[12]
rlabel metal1 6624 52462 6624 52462 0 chany_top_out_0[13]
rlabel metal1 7314 51442 7314 51442 0 chany_top_out_0[14]
rlabel metal1 6992 53618 6992 53618 0 chany_top_out_0[15]
rlabel metal2 7774 54376 7774 54376 0 chany_top_out_0[16]
rlabel metal2 7958 56236 7958 56236 0 chany_top_out_0[17]
rlabel metal2 8510 54070 8510 54070 0 chany_top_out_0[18]
rlabel metal1 8648 53618 8648 53618 0 chany_top_out_0[19]
rlabel metal1 2852 52666 2852 52666 0 chany_top_out_0[1]
rlabel metal1 9200 53142 9200 53142 0 chany_top_out_0[20]
rlabel metal2 9752 53550 9752 53550 0 chany_top_out_0[21]
rlabel metal1 9982 54264 9982 54264 0 chany_top_out_0[22]
rlabel metal2 10350 54614 10350 54614 0 chany_top_out_0[23]
rlabel metal1 10994 52530 10994 52530 0 chany_top_out_0[24]
rlabel metal2 11086 54920 11086 54920 0 chany_top_out_0[25]
rlabel metal1 11224 54230 11224 54230 0 chany_top_out_0[26]
rlabel metal1 12098 53006 12098 53006 0 chany_top_out_0[27]
rlabel metal1 12466 53618 12466 53618 0 chany_top_out_0[28]
rlabel metal1 12696 54094 12696 54094 0 chany_top_out_0[29]
rlabel metal2 2714 52972 2714 52972 0 chany_top_out_0[2]
rlabel metal2 2990 55711 2990 55711 0 chany_top_out_0[3]
rlabel metal2 3358 54070 3358 54070 0 chany_top_out_0[4]
rlabel metal1 3496 52530 3496 52530 0 chany_top_out_0[5]
rlabel metal2 4186 52972 4186 52972 0 chany_top_out_0[6]
rlabel metal1 4232 53142 4232 53142 0 chany_top_out_0[7]
rlabel metal1 4968 51918 4968 51918 0 chany_top_out_0[8]
rlabel metal2 5382 53244 5382 53244 0 chany_top_out_0[9]
rlabel metal1 18446 41990 18446 41990 0 clknet_0_prog_clk
rlabel metal1 5474 7922 5474 7922 0 clknet_4_0_0_prog_clk
rlabel metal1 6072 41650 6072 41650 0 clknet_4_10_0_prog_clk
rlabel metal1 13202 44404 13202 44404 0 clknet_4_11_0_prog_clk
rlabel metal1 19826 35122 19826 35122 0 clknet_4_12_0_prog_clk
rlabel metal1 22172 37230 22172 37230 0 clknet_4_13_0_prog_clk
rlabel metal1 19458 42126 19458 42126 0 clknet_4_14_0_prog_clk
rlabel metal1 22908 41038 22908 41038 0 clknet_4_15_0_prog_clk
rlabel metal2 11546 11968 11546 11968 0 clknet_4_1_0_prog_clk
rlabel metal1 9016 19890 9016 19890 0 clknet_4_2_0_prog_clk
rlabel metal1 9890 20842 9890 20842 0 clknet_4_3_0_prog_clk
rlabel metal1 18630 18190 18630 18190 0 clknet_4_4_0_prog_clk
rlabel metal1 18262 11798 18262 11798 0 clknet_4_5_0_prog_clk
rlabel metal2 15410 26180 15410 26180 0 clknet_4_6_0_prog_clk
rlabel metal1 23414 21556 23414 21556 0 clknet_4_7_0_prog_clk
rlabel metal1 6854 37162 6854 37162 0 clknet_4_8_0_prog_clk
rlabel metal1 12972 31246 12972 31246 0 clknet_4_9_0_prog_clk
rlabel metal3 1004 13804 1004 13804 0 gfpga_pad_io_soc_dir[0]
rlabel metal3 1004 16252 1004 16252 0 gfpga_pad_io_soc_dir[1]
rlabel metal3 1004 18700 1004 18700 0 gfpga_pad_io_soc_dir[2]
rlabel metal3 1004 21148 1004 21148 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 1564 33490 1564 33490 0 gfpga_pad_io_soc_in[0]
rlabel metal1 1932 36142 1932 36142 0 gfpga_pad_io_soc_in[1]
rlabel metal1 1564 38318 1564 38318 0 gfpga_pad_io_soc_in[2]
rlabel metal1 1564 41106 1564 41106 0 gfpga_pad_io_soc_in[3]
rlabel metal3 1004 23596 1004 23596 0 gfpga_pad_io_soc_out[0]
rlabel metal2 2806 26163 2806 26163 0 gfpga_pad_io_soc_out[1]
rlabel metal3 1004 28492 1004 28492 0 gfpga_pad_io_soc_out[2]
rlabel metal3 1004 30940 1004 30940 0 gfpga_pad_io_soc_out[3]
rlabel metal1 1518 43282 1518 43282 0 isol_n
rlabel metal1 4130 49606 4130 49606 0 net1
rlabel metal1 23299 39066 23299 39066 0 net10
rlabel metal1 18722 41446 18722 41446 0 net100
rlabel metal1 24978 38998 24978 38998 0 net101
rlabel metal1 23046 37774 23046 37774 0 net102
rlabel metal1 22218 40630 22218 40630 0 net103
rlabel metal2 23598 38488 23598 38488 0 net104
rlabel metal1 23506 32742 23506 32742 0 net105
rlabel metal2 23506 38080 23506 38080 0 net106
rlabel metal1 9430 43214 9430 43214 0 net107
rlabel metal1 16951 42126 16951 42126 0 net108
rlabel metal1 4278 50252 4278 50252 0 net109
rlabel metal1 20424 35734 20424 35734 0 net11
rlabel metal1 9246 43418 9246 43418 0 net110
rlabel metal2 18446 7310 18446 7310 0 net111
rlabel metal1 11086 43622 11086 43622 0 net112
rlabel metal1 22678 9996 22678 9996 0 net113
rlabel metal1 23920 9554 23920 9554 0 net114
rlabel metal1 23966 10608 23966 10608 0 net115
rlabel metal1 23276 11730 23276 11730 0 net116
rlabel metal1 22494 17034 22494 17034 0 net117
rlabel metal1 23184 17034 23184 17034 0 net118
rlabel metal1 23092 13974 23092 13974 0 net119
rlabel metal2 21114 38556 21114 38556 0 net12
rlabel metal1 24518 17510 24518 17510 0 net120
rlabel metal1 23046 19754 23046 19754 0 net121
rlabel metal1 24518 21862 24518 21862 0 net122
rlabel metal1 22862 5882 22862 5882 0 net123
rlabel metal2 22172 23052 22172 23052 0 net124
rlabel metal1 23874 17170 23874 17170 0 net125
rlabel metal2 24058 21726 24058 21726 0 net126
rlabel metal1 24058 19822 24058 19822 0 net127
rlabel metal1 22356 20434 22356 20434 0 net128
rlabel metal1 22448 20910 22448 20910 0 net129
rlabel metal1 22402 39576 22402 39576 0 net13
rlabel metal1 24610 20434 24610 20434 0 net130
rlabel metal1 23092 23086 23092 23086 0 net131
rlabel metal1 23184 24174 23184 24174 0 net132
rlabel metal1 23920 25874 23920 25874 0 net133
rlabel metal2 24886 5813 24886 5813 0 net134
rlabel metal2 17802 4964 17802 4964 0 net135
rlabel metal1 23184 7854 23184 7854 0 net136
rlabel metal1 24426 7718 24426 7718 0 net137
rlabel metal1 23782 9078 23782 9078 0 net138
rlabel metal1 24426 9894 24426 9894 0 net139
rlabel metal1 18492 24786 18492 24786 0 net14
rlabel metal2 23966 5491 23966 5491 0 net140
rlabel metal2 23966 9452 23966 9452 0 net141
rlabel metal1 13064 15606 13064 15606 0 net142
rlabel metal1 16790 4114 16790 4114 0 net143
rlabel metal2 19458 6222 19458 6222 0 net144
rlabel metal1 17848 3026 17848 3026 0 net145
rlabel metal2 18722 5507 18722 5507 0 net146
rlabel metal1 17158 3638 17158 3638 0 net147
rlabel metal1 18630 2482 18630 2482 0 net148
rlabel metal1 19044 4590 19044 4590 0 net149
rlabel metal1 23046 41004 23046 41004 0 net15
rlabel metal1 21160 3502 21160 3502 0 net150
rlabel metal2 19550 6051 19550 6051 0 net151
rlabel metal1 21114 8398 21114 8398 0 net152
rlabel metal2 12650 3604 12650 3604 0 net153
rlabel metal3 21160 4012 21160 4012 0 net154
rlabel metal1 20608 13838 20608 13838 0 net155
rlabel metal1 21942 5202 21942 5202 0 net156
rlabel metal1 21574 9418 21574 9418 0 net157
rlabel metal1 21528 5678 21528 5678 0 net158
rlabel metal1 21620 11594 21620 11594 0 net159
rlabel metal2 23966 41310 23966 41310 0 net16
rlabel metal1 22080 7378 22080 7378 0 net160
rlabel metal1 20700 6290 20700 6290 0 net161
rlabel metal1 20562 7718 20562 7718 0 net162
rlabel metal1 19044 6630 19044 6630 0 net163
rlabel metal1 13524 4114 13524 4114 0 net164
rlabel metal1 12420 10506 12420 10506 0 net165
rlabel metal2 14306 4963 14306 4963 0 net166
rlabel metal2 14674 7548 14674 7548 0 net167
rlabel metal2 15134 4369 15134 4369 0 net168
rlabel metal2 16882 6154 16882 6154 0 net169
rlabel metal1 24104 36006 24104 36006 0 net17
rlabel metal1 16836 3026 16836 3026 0 net170
rlabel metal1 16560 3502 16560 3502 0 net171
rlabel metal1 2760 49810 2760 49810 0 net172
rlabel metal1 3358 53550 3358 53550 0 net173
rlabel metal1 3404 54162 3404 54162 0 net174
rlabel metal1 5612 53074 5612 53074 0 net175
rlabel metal1 5612 52462 5612 52462 0 net176
rlabel metal1 8142 44438 8142 44438 0 net177
rlabel metal2 6854 52020 6854 52020 0 net178
rlabel metal1 8372 44982 8372 44982 0 net179
rlabel metal2 24794 37485 24794 37485 0 net18
rlabel metal2 4646 48756 4646 48756 0 net180
rlabel metal1 10396 43418 10396 43418 0 net181
rlabel metal1 9200 50490 9200 50490 0 net182
rlabel metal1 2254 50218 2254 50218 0 net183
rlabel metal1 10994 44438 10994 44438 0 net184
rlabel metal1 10442 44506 10442 44506 0 net185
rlabel metal1 11454 45050 11454 45050 0 net186
rlabel metal1 9522 49878 9522 49878 0 net187
rlabel metal1 10212 50966 10212 50966 0 net188
rlabel metal1 11500 44914 11500 44914 0 net189
rlabel metal3 23575 45628 23575 45628 0 net19
rlabel metal1 10120 51578 10120 51578 0 net190
rlabel metal1 11822 52122 11822 52122 0 net191
rlabel metal2 12650 53108 12650 53108 0 net192
rlabel metal2 12374 53142 12374 53142 0 net193
rlabel metal1 2530 50932 2530 50932 0 net194
rlabel metal1 2254 51340 2254 51340 0 net195
rlabel metal1 4968 42738 4968 42738 0 net196
rlabel metal1 3726 52462 3726 52462 0 net197
rlabel metal1 4692 42262 4692 42262 0 net198
rlabel metal1 2990 53040 2990 53040 0 net199
rlabel metal1 2208 3978 2208 3978 0 net2
rlabel metal1 25392 47158 25392 47158 0 net20
rlabel metal1 5796 43962 5796 43962 0 net200
rlabel metal1 6118 51374 6118 51374 0 net201
rlabel metal2 1794 14892 1794 14892 0 net202
rlabel metal1 1794 19482 1794 19482 0 net203
rlabel metal2 1794 19754 1794 19754 0 net204
rlabel metal1 1840 21522 1840 21522 0 net205
rlabel metal1 1932 22746 1932 22746 0 net206
rlabel metal1 1932 26350 1932 26350 0 net207
rlabel metal1 1978 26010 1978 26010 0 net208
rlabel metal1 2024 28186 2024 28186 0 net209
rlabel metal3 22839 40596 22839 40596 0 net21
rlabel metal2 25346 1989 25346 1989 0 net210
rlabel metal2 17618 21182 17618 21182 0 net211
rlabel metal1 12926 28186 12926 28186 0 net212
rlabel metal2 21482 33728 21482 33728 0 net213
rlabel metal1 24978 23120 24978 23120 0 net214
rlabel metal1 14904 37842 14904 37842 0 net215
rlabel metal1 17158 21998 17158 21998 0 net216
rlabel metal2 20930 29376 20930 29376 0 net217
rlabel metal1 16928 36074 16928 36074 0 net218
rlabel metal1 17986 36890 17986 36890 0 net219
rlabel metal1 18952 42330 18952 42330 0 net22
rlabel metal1 17066 37978 17066 37978 0 net220
rlabel metal1 14536 39066 14536 39066 0 net221
rlabel metal1 13432 37230 13432 37230 0 net222
rlabel metal1 23460 39338 23460 39338 0 net223
rlabel metal1 12788 32402 12788 32402 0 net224
rlabel metal1 11270 30226 11270 30226 0 net225
rlabel metal1 13018 24242 13018 24242 0 net226
rlabel metal2 11822 25534 11822 25534 0 net227
rlabel metal2 9430 25602 9430 25602 0 net228
rlabel metal2 9154 26690 9154 26690 0 net229
rlabel metal1 19366 42534 19366 42534 0 net23
rlabel metal1 7958 24922 7958 24922 0 net230
rlabel metal1 10074 24820 10074 24820 0 net231
rlabel metal1 6394 9554 6394 9554 0 net232
rlabel metal2 14766 11458 14766 11458 0 net233
rlabel metal1 20608 32878 20608 32878 0 net234
rlabel metal2 17250 13056 17250 13056 0 net235
rlabel metal1 18768 15130 18768 15130 0 net236
rlabel metal2 20470 16830 20470 16830 0 net237
rlabel metal1 22356 15130 22356 15130 0 net238
rlabel metal1 20056 16082 20056 16082 0 net239
rlabel metal1 23092 49946 23092 49946 0 net24
rlabel metal1 21758 12206 21758 12206 0 net240
rlabel metal1 19596 10778 19596 10778 0 net241
rlabel metal1 19642 13294 19642 13294 0 net242
rlabel metal1 23184 34714 23184 34714 0 net243
rlabel metal2 22034 41344 22034 41344 0 net244
rlabel metal1 9936 37842 9936 37842 0 net245
rlabel metal1 7912 30770 7912 30770 0 net246
rlabel metal1 7406 32538 7406 32538 0 net247
rlabel metal1 13800 42194 13800 42194 0 net248
rlabel metal2 9798 33150 9798 33150 0 net249
rlabel metal1 16974 24718 16974 24718 0 net25
rlabel metal2 5382 32980 5382 32980 0 net250
rlabel metal1 8280 38318 8280 38318 0 net251
rlabel metal1 11270 37978 11270 37978 0 net252
rlabel metal1 10902 39066 10902 39066 0 net253
rlabel metal1 14582 35802 14582 35802 0 net254
rlabel metal1 9476 31450 9476 31450 0 net255
rlabel metal2 11730 23358 11730 23358 0 net256
rlabel metal1 12880 20434 12880 20434 0 net257
rlabel metal1 9430 16558 9430 16558 0 net258
rlabel metal1 9844 23834 9844 23834 0 net259
rlabel metal1 15778 31790 15778 31790 0 net26
rlabel metal2 13938 22100 13938 22100 0 net260
rlabel metal1 14076 24242 14076 24242 0 net261
rlabel metal1 20332 26962 20332 26962 0 net262
rlabel metal2 21666 25534 21666 25534 0 net263
rlabel metal2 17250 29716 17250 29716 0 net264
rlabel metal1 20102 36006 20102 36006 0 net27
rlabel metal1 19596 38182 19596 38182 0 net28
rlabel metal1 18998 35802 18998 35802 0 net29
rlabel metal1 19734 24718 19734 24718 0 net3
rlabel metal1 22770 33932 22770 33932 0 net30
rlabel metal1 25162 32776 25162 32776 0 net31
rlabel metal1 17296 32470 17296 32470 0 net32
rlabel metal1 3680 3638 3680 3638 0 net33
rlabel metal1 6578 44370 6578 44370 0 net34
rlabel metal2 5934 4743 5934 4743 0 net35
rlabel metal2 16146 3876 16146 3876 0 net36
rlabel metal1 8004 44778 8004 44778 0 net37
rlabel metal2 7038 4403 7038 4403 0 net38
rlabel metal1 9200 44370 9200 44370 0 net39
rlabel metal1 25162 34680 25162 34680 0 net4
rlabel metal1 7866 2482 7866 2482 0 net40
rlabel metal2 8234 3944 8234 3944 0 net41
rlabel metal1 7498 3162 7498 3162 0 net42
rlabel metal1 10396 42534 10396 42534 0 net43
rlabel metal1 3496 2890 3496 2890 0 net44
rlabel metal1 10396 5542 10396 5542 0 net45
rlabel metal1 9430 3706 9430 3706 0 net46
rlabel metal2 10074 4658 10074 4658 0 net47
rlabel metal1 10810 2618 10810 2618 0 net48
rlabel metal1 12742 3094 12742 3094 0 net49
rlabel metal1 25070 34918 25070 34918 0 net5
rlabel metal1 13846 6358 13846 6358 0 net50
rlabel metal1 12420 44846 12420 44846 0 net51
rlabel metal1 13984 3910 13984 3910 0 net52
rlabel metal1 13570 2278 13570 2278 0 net53
rlabel metal1 11730 2550 11730 2550 0 net54
rlabel metal1 5934 41990 5934 41990 0 net55
rlabel metal1 4094 42194 4094 42194 0 net56
rlabel metal2 3542 7548 3542 7548 0 net57
rlabel metal2 2622 4148 2622 4148 0 net58
rlabel metal1 4094 2550 4094 2550 0 net59
rlabel metal1 21528 33082 21528 33082 0 net6
rlabel metal1 6578 42194 6578 42194 0 net60
rlabel metal1 5957 2482 5957 2482 0 net61
rlabel metal2 5290 7072 5290 7072 0 net62
rlabel metal1 12236 49742 12236 49742 0 net63
rlabel metal2 16882 52122 16882 52122 0 net64
rlabel metal1 15548 43078 15548 43078 0 net65
rlabel metal1 17940 47770 17940 47770 0 net66
rlabel metal1 18170 48246 18170 48246 0 net67
rlabel metal1 18446 47702 18446 47702 0 net68
rlabel metal1 18032 43690 18032 43690 0 net69
rlabel metal2 20102 36856 20102 36856 0 net7
rlabel metal2 18630 49980 18630 49980 0 net70
rlabel metal1 16882 18394 16882 18394 0 net71
rlabel metal3 20769 44268 20769 44268 0 net72
rlabel metal1 21068 47226 21068 47226 0 net73
rlabel metal1 13616 52462 13616 52462 0 net74
rlabel metal2 20194 49436 20194 49436 0 net75
rlabel via2 21666 43061 21666 43061 0 net76
rlabel metal1 21252 43622 21252 43622 0 net77
rlabel metal1 22080 46682 22080 46682 0 net78
rlabel metal2 21390 49708 21390 49708 0 net79
rlabel metal1 25162 37162 25162 37162 0 net8
rlabel metal2 22494 50252 22494 50252 0 net80
rlabel metal1 20838 11798 20838 11798 0 net81
rlabel metal1 22448 43418 22448 43418 0 net82
rlabel metal1 22356 43826 22356 43826 0 net83
rlabel metal1 23368 46682 23368 46682 0 net84
rlabel via3 14053 52564 14053 52564 0 net85
rlabel metal3 14559 52972 14559 52972 0 net86
rlabel metal1 14766 43418 14766 43418 0 net87
rlabel metal1 13984 12410 13984 12410 0 net88
rlabel metal1 15548 53958 15548 53958 0 net89
rlabel metal1 23644 36074 23644 36074 0 net9
rlabel via3 16445 52564 16445 52564 0 net90
rlabel metal2 15962 50320 15962 50320 0 net91
rlabel via2 17526 11883 17526 11883 0 net92
rlabel metal1 2576 33286 2576 33286 0 net93
rlabel metal1 2530 36006 2530 36006 0 net94
rlabel metal1 2852 38182 2852 38182 0 net95
rlabel metal2 1610 35836 1610 35836 0 net96
rlabel metal1 2944 43146 2944 43146 0 net97
rlabel metal1 24794 3162 24794 3162 0 net98
rlabel metal1 23230 37842 23230 37842 0 net99
rlabel metal2 23782 7300 23782 7300 0 prog_clk
rlabel metal2 23598 3230 23598 3230 0 prog_reset
rlabel metal2 25070 50711 25070 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 25530 51561 25530 51561 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 24794 52309 24794 52309 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 25070 53023 25070 53023 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 24978 53975 24978 53975 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 24932 53550 24932 53550 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 25446 55420 25446 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel via2 23437 56100 23437 56100 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal3 1924 4012 1924 4012 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 1878 6460 1878 6460 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1878 8908 1878 8908 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1303 11356 1303 11356 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 19044 13838 19044 13838 0 sb_0__1_.mem_bottom_track_1.ccff_head
rlabel metal1 16100 22066 16100 22066 0 sb_0__1_.mem_bottom_track_1.ccff_tail
rlabel metal1 16928 18802 16928 18802 0 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 14398 21930 14398 21930 0 sb_0__1_.mem_bottom_track_1.mem_out\[1\]
rlabel metal1 20562 21862 20562 21862 0 sb_0__1_.mem_bottom_track_11.ccff_head
rlabel metal1 17388 25126 17388 25126 0 sb_0__1_.mem_bottom_track_11.ccff_tail
rlabel metal1 18906 34034 18906 34034 0 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
rlabel metal1 17480 26554 17480 26554 0 sb_0__1_.mem_bottom_track_11.mem_out\[1\]
rlabel metal1 20562 25840 20562 25840 0 sb_0__1_.mem_bottom_track_13.ccff_tail
rlabel metal1 20562 34442 20562 34442 0 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
rlabel metal2 21206 29172 21206 29172 0 sb_0__1_.mem_bottom_track_13.mem_out\[1\]
rlabel metal2 24702 26350 24702 26350 0 sb_0__1_.mem_bottom_track_21.ccff_tail
rlabel metal1 22356 34442 22356 34442 0 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
rlabel metal2 22678 25959 22678 25959 0 sb_0__1_.mem_bottom_track_21.mem_out\[1\]
rlabel metal1 15548 32334 15548 32334 0 sb_0__1_.mem_bottom_track_29.ccff_tail
rlabel metal1 16882 32946 16882 32946 0 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
rlabel metal1 17710 32334 17710 32334 0 sb_0__1_.mem_bottom_track_29.mem_out\[1\]
rlabel metal2 21666 20570 21666 20570 0 sb_0__1_.mem_bottom_track_3.ccff_tail
rlabel metal1 19872 27982 19872 27982 0 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 19780 20842 19780 20842 0 sb_0__1_.mem_bottom_track_3.mem_out\[1\]
rlabel metal1 15502 33898 15502 33898 0 sb_0__1_.mem_bottom_track_37.ccff_tail
rlabel metal1 18906 38794 18906 38794 0 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
rlabel metal1 14674 33286 14674 33286 0 sb_0__1_.mem_bottom_track_37.mem_out\[1\]
rlabel metal1 19734 33626 19734 33626 0 sb_0__1_.mem_bottom_track_45.ccff_tail
rlabel metal1 20325 35258 20325 35258 0 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
rlabel metal1 21436 34034 21436 34034 0 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
rlabel metal1 23138 21454 23138 21454 0 sb_0__1_.mem_bottom_track_5.ccff_tail
rlabel metal1 20424 29070 20424 29070 0 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 24656 23630 24656 23630 0 sb_0__1_.mem_bottom_track_5.mem_out\[1\]
rlabel metal1 12742 43826 12742 43826 0 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
rlabel metal2 22862 21794 22862 21794 0 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
rlabel metal1 19218 22202 19218 22202 0 sb_0__1_.mem_bottom_track_7.mem_out\[1\]
rlabel metal1 17802 38182 17802 38182 0 sb_0__1_.mem_right_track_0.ccff_head
rlabel metal1 23690 29682 23690 29682 0 sb_0__1_.mem_right_track_0.ccff_tail
rlabel metal2 21574 34238 21574 34238 0 sb_0__1_.mem_right_track_0.mem_out\[0\]
rlabel metal1 23046 31858 23046 31858 0 sb_0__1_.mem_right_track_0.mem_out\[1\]
rlabel metal1 23414 44710 23414 44710 0 sb_0__1_.mem_right_track_10.ccff_head
rlabel metal2 21206 43044 21206 43044 0 sb_0__1_.mem_right_track_10.ccff_tail
rlabel metal1 20095 42874 20095 42874 0 sb_0__1_.mem_right_track_10.mem_out\[0\]
rlabel metal1 19596 41514 19596 41514 0 sb_0__1_.mem_right_track_10.mem_out\[1\]
rlabel metal2 20102 44404 20102 44404 0 sb_0__1_.mem_right_track_12.ccff_tail
rlabel metal2 19826 44642 19826 44642 0 sb_0__1_.mem_right_track_12.mem_out\[0\]
rlabel metal1 19182 43214 19182 43214 0 sb_0__1_.mem_right_track_12.mem_out\[1\]
rlabel metal1 18722 44166 18722 44166 0 sb_0__1_.mem_right_track_14.ccff_tail
rlabel metal2 19366 46036 19366 46036 0 sb_0__1_.mem_right_track_14.mem_out\[0\]
rlabel metal1 18906 41650 18906 41650 0 sb_0__1_.mem_right_track_14.mem_out\[1\]
rlabel metal1 16928 44710 16928 44710 0 sb_0__1_.mem_right_track_16.ccff_tail
rlabel metal2 18722 47396 18722 47396 0 sb_0__1_.mem_right_track_16.mem_out\[0\]
rlabel metal1 17434 43214 17434 43214 0 sb_0__1_.mem_right_track_16.mem_out\[1\]
rlabel metal1 15502 40902 15502 40902 0 sb_0__1_.mem_right_track_18.ccff_tail
rlabel metal1 17434 47532 17434 47532 0 sb_0__1_.mem_right_track_18.mem_out\[0\]
rlabel metal2 16146 43452 16146 43452 0 sb_0__1_.mem_right_track_18.mem_out\[1\]
rlabel metal1 25438 43078 25438 43078 0 sb_0__1_.mem_right_track_2.ccff_tail
rlabel metal1 22816 41174 22816 41174 0 sb_0__1_.mem_right_track_2.mem_out\[0\]
rlabel metal1 23460 41650 23460 41650 0 sb_0__1_.mem_right_track_2.mem_out\[1\]
rlabel metal1 14168 34510 14168 34510 0 sb_0__1_.mem_right_track_20.ccff_tail
rlabel metal1 14996 43146 14996 43146 0 sb_0__1_.mem_right_track_20.mem_out\[0\]
rlabel metal2 13938 37706 13938 37706 0 sb_0__1_.mem_right_track_20.mem_out\[1\]
rlabel metal1 12811 29682 12811 29682 0 sb_0__1_.mem_right_track_22.ccff_tail
rlabel metal1 13570 35530 13570 35530 0 sb_0__1_.mem_right_track_22.mem_out\[0\]
rlabel metal1 13570 34068 13570 34068 0 sb_0__1_.mem_right_track_22.mem_out\[1\]
rlabel metal1 14352 26758 14352 26758 0 sb_0__1_.mem_right_track_24.ccff_tail
rlabel metal2 12834 27200 12834 27200 0 sb_0__1_.mem_right_track_24.mem_out\[0\]
rlabel metal2 12926 27200 12926 27200 0 sb_0__1_.mem_right_track_26.ccff_tail
rlabel metal1 14720 25806 14720 25806 0 sb_0__1_.mem_right_track_26.mem_out\[0\]
rlabel metal1 10948 27914 10948 27914 0 sb_0__1_.mem_right_track_28.ccff_tail
rlabel metal2 13662 27574 13662 27574 0 sb_0__1_.mem_right_track_28.mem_out\[0\]
rlabel metal1 9108 28594 9108 28594 0 sb_0__1_.mem_right_track_30.ccff_tail
rlabel metal1 12466 29104 12466 29104 0 sb_0__1_.mem_right_track_30.mem_out\[0\]
rlabel metal1 9016 26826 9016 26826 0 sb_0__1_.mem_right_track_32.ccff_tail
rlabel metal1 7912 27574 7912 27574 0 sb_0__1_.mem_right_track_32.mem_out\[0\]
rlabel metal2 8602 24752 8602 24752 0 sb_0__1_.mem_right_track_34.ccff_tail
rlabel metal1 14306 29172 14306 29172 0 sb_0__1_.mem_right_track_34.mem_out\[0\]
rlabel metal2 8786 12954 8786 12954 0 sb_0__1_.mem_right_track_36.ccff_tail
rlabel metal1 8142 23834 8142 23834 0 sb_0__1_.mem_right_track_36.mem_out\[0\]
rlabel metal1 7728 18190 7728 18190 0 sb_0__1_.mem_right_track_36.mem_out\[1\]
rlabel metal1 13616 11662 13616 11662 0 sb_0__1_.mem_right_track_38.ccff_tail
rlabel metal1 12834 13804 12834 13804 0 sb_0__1_.mem_right_track_38.mem_out\[0\]
rlabel metal2 23414 34816 23414 34816 0 sb_0__1_.mem_right_track_4.ccff_tail
rlabel metal1 24334 42330 24334 42330 0 sb_0__1_.mem_right_track_4.mem_out\[0\]
rlabel metal1 23782 38726 23782 38726 0 sb_0__1_.mem_right_track_4.mem_out\[1\]
rlabel metal1 16146 13498 16146 13498 0 sb_0__1_.mem_right_track_40.ccff_tail
rlabel metal2 14858 14076 14858 14076 0 sb_0__1_.mem_right_track_40.mem_out\[0\]
rlabel metal2 18630 16660 18630 16660 0 sb_0__1_.mem_right_track_44.ccff_tail
rlabel metal2 17158 16932 17158 16932 0 sb_0__1_.mem_right_track_44.mem_out\[0\]
rlabel metal2 20194 17816 20194 17816 0 sb_0__1_.mem_right_track_46.ccff_tail
rlabel metal1 19182 18360 19182 18360 0 sb_0__1_.mem_right_track_46.mem_out\[0\]
rlabel metal1 23230 17850 23230 17850 0 sb_0__1_.mem_right_track_48.ccff_tail
rlabel metal1 22310 17714 22310 17714 0 sb_0__1_.mem_right_track_48.mem_out\[0\]
rlabel metal2 21850 18122 21850 18122 0 sb_0__1_.mem_right_track_50.ccff_tail
rlabel metal1 22540 19278 22540 19278 0 sb_0__1_.mem_right_track_50.mem_out\[0\]
rlabel metal1 21804 12274 21804 12274 0 sb_0__1_.mem_right_track_52.ccff_tail
rlabel metal2 21206 15436 21206 15436 0 sb_0__1_.mem_right_track_52.mem_out\[0\]
rlabel metal2 20010 12070 20010 12070 0 sb_0__1_.mem_right_track_54.ccff_tail
rlabel metal1 18492 13362 18492 13362 0 sb_0__1_.mem_right_track_54.mem_out\[0\]
rlabel metal1 18216 12410 18216 12410 0 sb_0__1_.mem_right_track_56.mem_out\[0\]
rlabel metal1 24932 37774 24932 37774 0 sb_0__1_.mem_right_track_6.ccff_tail
rlabel metal1 22908 36822 22908 36822 0 sb_0__1_.mem_right_track_6.mem_out\[0\]
rlabel metal2 23874 38148 23874 38148 0 sb_0__1_.mem_right_track_6.mem_out\[1\]
rlabel metal1 22632 44302 22632 44302 0 sb_0__1_.mem_right_track_8.mem_out\[0\]
rlabel metal2 22586 44642 22586 44642 0 sb_0__1_.mem_right_track_8.mem_out\[1\]
rlabel metal2 12190 46444 12190 46444 0 sb_0__1_.mem_top_track_0.ccff_tail
rlabel metal1 17710 42806 17710 42806 0 sb_0__1_.mem_top_track_0.mem_out\[0\]
rlabel metal1 12466 44268 12466 44268 0 sb_0__1_.mem_top_track_0.mem_out\[1\]
rlabel metal1 7544 38386 7544 38386 0 sb_0__1_.mem_top_track_10.ccff_head
rlabel metal2 6026 36244 6026 36244 0 sb_0__1_.mem_top_track_10.ccff_tail
rlabel metal2 16790 37502 16790 37502 0 sb_0__1_.mem_top_track_10.mem_out\[0\]
rlabel metal1 9476 34034 9476 34034 0 sb_0__1_.mem_top_track_10.mem_out\[1\]
rlabel metal1 7682 32334 7682 32334 0 sb_0__1_.mem_top_track_12.ccff_tail
rlabel metal2 13754 33286 13754 33286 0 sb_0__1_.mem_top_track_12.mem_out\[0\]
rlabel metal1 8234 32946 8234 32946 0 sb_0__1_.mem_top_track_12.mem_out\[1\]
rlabel metal1 13110 44914 13110 44914 0 sb_0__1_.mem_top_track_2.ccff_tail
rlabel metal1 17434 42194 17434 42194 0 sb_0__1_.mem_top_track_2.mem_out\[0\]
rlabel metal1 14582 44302 14582 44302 0 sb_0__1_.mem_top_track_2.mem_out\[1\]
rlabel metal2 9614 35700 9614 35700 0 sb_0__1_.mem_top_track_20.ccff_tail
rlabel metal1 17020 31382 17020 31382 0 sb_0__1_.mem_top_track_20.mem_out\[0\]
rlabel metal1 10067 34374 10067 34374 0 sb_0__1_.mem_top_track_20.mem_out\[1\]
rlabel metal2 5842 38522 5842 38522 0 sb_0__1_.mem_top_track_28.ccff_tail
rlabel metal2 13570 34612 13570 34612 0 sb_0__1_.mem_top_track_28.mem_out\[0\]
rlabel metal1 7774 35258 7774 35258 0 sb_0__1_.mem_top_track_28.mem_out\[1\]
rlabel metal1 8372 42126 8372 42126 0 sb_0__1_.mem_top_track_36.ccff_tail
rlabel metal1 7452 40562 7452 40562 0 sb_0__1_.mem_top_track_36.mem_out\[0\]
rlabel metal1 6210 41480 6210 41480 0 sb_0__1_.mem_top_track_36.mem_out\[1\]
rlabel metal1 10994 41650 10994 41650 0 sb_0__1_.mem_top_track_4.ccff_tail
rlabel metal1 14122 43384 14122 43384 0 sb_0__1_.mem_top_track_4.mem_out\[0\]
rlabel metal2 12742 38828 12742 38828 0 sb_0__1_.mem_top_track_4.mem_out\[1\]
rlabel metal1 12558 42568 12558 42568 0 sb_0__1_.mem_top_track_44.ccff_tail
rlabel metal1 10994 42602 10994 42602 0 sb_0__1_.mem_top_track_44.mem_out\[0\]
rlabel metal1 16698 42534 16698 42534 0 sb_0__1_.mem_top_track_52.mem_out\[0\]
rlabel metal1 16146 38386 16146 38386 0 sb_0__1_.mem_top_track_52.mem_out\[1\]
rlabel metal1 8924 31926 8924 31926 0 sb_0__1_.mem_top_track_6.mem_out\[0\]
rlabel metal2 8602 37842 8602 37842 0 sb_0__1_.mem_top_track_6.mem_out\[1\]
rlabel metal1 18124 6766 18124 6766 0 sb_0__1_.mux_bottom_track_1.out
rlabel metal1 15732 26010 15732 26010 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17894 32198 17894 32198 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13846 21590 13846 21590 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15088 22746 15088 22746 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13708 21658 13708 21658 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15180 22406 15180 22406 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 17342 9792 17342 9792 0 sb_0__1_.mux_bottom_track_11.out
rlabel metal1 17434 28594 17434 28594 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18124 28526 18124 28526 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16882 25024 16882 25024 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14306 24650 14306 24650 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16928 24242 16928 24242 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 16790 24820 16790 24820 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16882 17170 16882 17170 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 18906 9622 18906 9622 0 sb_0__1_.mux_bottom_track_13.out
rlabel metal1 20102 29716 20102 29716 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20378 29614 20378 29614 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18814 27098 18814 27098 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20378 27744 20378 27744 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19918 26010 19918 26010 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18814 19822 18814 19822 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 20838 8534 20838 8534 0 sb_0__1_.mux_bottom_track_21.out
rlabel metal1 21850 29478 21850 29478 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21988 29614 21988 29614 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21114 26452 21114 26452 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21574 26826 21574 26826 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24932 24038 24932 24038 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 22494 16116 22494 16116 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16284 9622 16284 9622 0 sb_0__1_.mux_bottom_track_29.out
rlabel metal1 16790 32538 16790 32538 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17250 34476 17250 34476 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17434 29274 17434 29274 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16514 28526 16514 28526 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 16054 28764 16054 28764 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15732 28390 15732 28390 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 17434 12036 17434 12036 0 sb_0__1_.mux_bottom_track_3.out
rlabel metal1 19504 25330 19504 25330 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19642 25262 19642 25262 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19504 20570 19504 20570 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19366 20808 19366 20808 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19826 17612 19826 17612 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14168 10030 14168 10030 0 sb_0__1_.mux_bottom_track_37.out
rlabel metal1 16146 34646 16146 34646 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17894 34714 17894 34714 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14904 34714 14904 34714 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13478 28730 13478 28730 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13340 21998 13340 21998 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17618 9962 17618 9962 0 sb_0__1_.mux_bottom_track_45.out
rlabel metal2 21298 37468 21298 37468 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20194 31790 20194 31790 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20838 34102 20838 34102 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18860 20434 18860 20434 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20976 7854 20976 7854 0 sb_0__1_.mux_bottom_track_5.out
rlabel metal1 20102 29240 20102 29240 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22770 26350 22770 26350 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21183 24582 21183 24582 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22724 26486 22724 26486 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23000 21658 23000 21658 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 22218 21318 22218 21318 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11178 12138 11178 12138 0 sb_0__1_.mux_bottom_track_53.out
rlabel metal1 13662 38760 13662 38760 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12236 37162 12236 37162 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10902 37094 10902 37094 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19044 8534 19044 8534 0 sb_0__1_.mux_bottom_track_7.out
rlabel metal1 19458 26418 19458 26418 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20654 28968 20654 28968 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18308 24582 18308 24582 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16882 21896 16882 21896 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19734 24582 19734 24582 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18860 21862 18860 21862 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 19044 19414 19044 19414 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 22632 26962 22632 26962 0 sb_0__1_.mux_right_track_0.out
rlabel metal2 21390 32028 21390 32028 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21620 31654 21620 31654 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22678 31926 22678 31926 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23322 29240 23322 29240 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24794 28560 24794 28560 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23414 32470 23414 32470 0 sb_0__1_.mux_right_track_10.out
rlabel metal1 20838 45798 20838 45798 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20240 40154 20240 40154 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20700 38386 20700 38386 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17342 36278 17342 36278 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22034 32402 22034 32402 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23690 32538 23690 32538 0 sb_0__1_.mux_right_track_12.out
rlabel metal1 19826 45798 19826 45798 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19688 39474 19688 39474 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19228 39338 19228 39338 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19504 39270 19504 39270 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23092 33082 23092 33082 0 sb_0__1_.mux_right_track_14.out
rlabel metal1 18584 41650 18584 41650 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 18492 41446 18492 41446 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16928 37706 16928 37706 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22402 34068 22402 34068 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20102 29070 20102 29070 0 sb_0__1_.mux_right_track_16.out
rlabel metal1 17802 47430 17802 47430 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17112 40562 17112 40562 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15732 39610 15732 39610 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20286 32470 20286 32470 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21924 24106 21924 24106 0 sb_0__1_.mux_right_track_18.out
rlabel metal2 16652 41582 16652 41582 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16376 41446 16376 41446 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15640 37230 15640 37230 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 16376 34442 16376 34442 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24656 29206 24656 29206 0 sb_0__1_.mux_right_track_2.out
rlabel metal1 22816 46342 22816 46342 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22310 40562 22310 40562 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20332 37978 20332 37978 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 25070 40596 25070 40596 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24978 39474 24978 39474 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24702 33966 24702 33966 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24150 21896 24150 21896 0 sb_0__1_.mux_right_track_20.out
rlabel metal1 14260 36822 14260 36822 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14628 32946 14628 32946 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14674 32640 14674 32640 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14398 32742 14398 32742 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19964 19890 19964 19890 0 sb_0__1_.mux_right_track_22.out
rlabel metal1 13018 40630 13018 40630 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12926 33830 12926 33830 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13018 29682 13018 29682 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17572 24174 17572 24174 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 24886 19244 24886 19244 0 sb_0__1_.mux_right_track_24.out
rlabel metal1 15180 24786 15180 24786 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13938 24922 13938 24922 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18308 20910 18308 20910 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21298 18224 21298 18224 0 sb_0__1_.mux_right_track_26.out
rlabel metal1 15180 27098 15180 27098 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13570 26180 13570 26180 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18078 21522 18078 21522 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22540 17170 22540 17170 0 sb_0__1_.mux_right_track_28.out
rlabel metal1 13478 26350 13478 26350 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12558 26078 12558 26078 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13938 21454 13938 21454 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21114 19448 21114 19448 0 sb_0__1_.mux_right_track_30.out
rlabel metal2 10902 27506 10902 27506 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10672 26010 10672 26010 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16238 21454 16238 21454 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21298 16014 21298 16014 0 sb_0__1_.mux_right_track_32.out
rlabel metal1 10672 25262 10672 25262 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8050 24650 8050 24650 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15686 20468 15686 20468 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21620 15402 21620 15402 0 sb_0__1_.mux_right_track_34.out
rlabel metal2 11270 26758 11270 26758 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11178 24378 11178 24378 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17066 19822 17066 19822 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20838 10778 20838 10778 0 sb_0__1_.mux_right_track_36.out
rlabel metal1 7636 18394 7636 18394 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 8694 15504 8694 15504 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7590 12818 7590 12818 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14858 10676 14858 10676 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22218 10064 22218 10064 0 sb_0__1_.mux_right_track_38.out
rlabel metal1 14950 11798 14950 11798 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15778 11084 15778 11084 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25116 27030 25116 27030 0 sb_0__1_.mux_right_track_4.out
rlabel metal1 21988 43622 21988 43622 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22816 38250 22816 38250 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22540 34034 22540 34034 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20378 33082 20378 33082 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22402 33830 22402 33830 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23414 10676 23414 10676 0 sb_0__1_.mux_right_track_40.out
rlabel metal1 17204 12886 17204 12886 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19642 10642 19642 10642 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24012 9962 24012 9962 0 sb_0__1_.mux_right_track_44.out
rlabel metal2 18906 16354 18906 16354 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20010 12206 20010 12206 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24748 8942 24748 8942 0 sb_0__1_.mux_right_track_46.out
rlabel metal2 20562 17986 20562 17986 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22862 14518 22862 14518 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24886 9962 24886 9962 0 sb_0__1_.mux_right_track_48.out
rlabel metal2 21574 17850 21574 17850 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23414 12240 23414 12240 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23690 8942 23690 8942 0 sb_0__1_.mux_right_track_50.out
rlabel metal1 21620 25670 21620 25670 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19274 17714 19274 17714 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21298 13940 21298 13940 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23000 4658 23000 4658 0 sb_0__1_.mux_right_track_52.out
rlabel metal1 21436 12274 21436 12274 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22034 9554 22034 9554 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24012 4590 24012 4590 0 sb_0__1_.mux_right_track_54.out
rlabel metal1 18722 10574 18722 10574 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21758 9690 21758 9690 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23644 5678 23644 5678 0 sb_0__1_.mux_right_track_56.out
rlabel metal2 19918 14484 19918 14484 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20654 10030 20654 10030 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24564 26350 24564 26350 0 sb_0__1_.mux_right_track_6.out
rlabel metal1 25024 38318 25024 38318 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24702 38080 24702 38080 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 23690 34034 23690 34034 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23782 37196 23782 37196 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23690 35943 23690 35943 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23828 31450 23828 31450 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24564 34714 24564 34714 0 sb_0__1_.mux_right_track_8.out
rlabel metal1 22172 42738 22172 42738 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22218 41616 22218 41616 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21620 41514 21620 41514 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 22954 40477 22954 40477 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22724 40494 22724 40494 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal3 23276 37196 23276 37196 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11822 49402 11822 49402 0 sb_0__1_.mux_top_track_0.out
rlabel metal1 10166 43146 10166 43146 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17158 42772 17158 42772 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14950 39168 14950 39168 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11086 37706 11086 37706 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11546 44506 11546 44506 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11408 45866 11408 45866 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 10718 47668 10718 47668 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7958 44506 7958 44506 0 sb_0__1_.mux_top_track_10.out
rlabel metal1 9430 38386 9430 38386 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16836 37434 16836 37434 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12696 30906 12696 30906 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8602 33898 8602 33898 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8188 36890 8188 36890 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 9154 35462 9154 35462 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7866 44370 7866 44370 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8464 49810 8464 49810 0 sb_0__1_.mux_top_track_12.out
rlabel metal1 10856 33626 10856 33626 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11638 32742 11638 32742 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7866 32810 7866 32810 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10396 33626 10396 33626 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 7636 33082 7636 33082 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7452 43282 7452 43282 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12788 48858 12788 48858 0 sb_0__1_.mux_top_track_2.out
rlabel metal1 16376 42330 16376 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15778 41956 15778 41956 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13018 42126 13018 42126 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15318 42330 15318 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13248 42330 13248 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12788 45050 12788 45050 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8924 50286 8924 50286 0 sb_0__1_.mux_top_track_20.out
rlabel metal1 14030 35054 14030 35054 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17066 34578 17066 34578 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9706 32742 9706 32742 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 10626 36006 10626 36006 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9384 33082 9384 33082 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8832 43758 8832 43758 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 5842 47396 5842 47396 0 sb_0__1_.mux_top_track_28.out
rlabel metal1 9890 36142 9890 36142 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12834 33626 12834 33626 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8510 36346 8510 36346 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 5014 35190 5014 35190 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 5704 44370 5704 44370 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7360 46682 7360 46682 0 sb_0__1_.mux_top_track_36.out
rlabel metal1 11914 38386 11914 38386 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11040 38454 11040 38454 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8326 41990 8326 41990 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9522 41990 9522 41990 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 10902 49334 10902 49334 0 sb_0__1_.mux_top_track_4.out
rlabel metal1 14996 38318 14996 38318 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17250 38233 17250 38233 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11040 33082 11040 33082 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12696 41446 12696 41446 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10764 38522 10764 38522 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10902 41786 10902 41786 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9108 47770 9108 47770 0 sb_0__1_.mux_top_track_44.out
rlabel metal1 13708 42262 13708 42262 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11684 42194 11684 42194 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10580 47634 10580 47634 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8878 46070 8878 46070 0 sb_0__1_.mux_top_track_52.out
rlabel metal1 20286 38998 20286 38998 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17618 39066 17618 39066 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14858 36346 14858 36346 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10626 45934 10626 45934 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9200 46138 9200 46138 0 sb_0__1_.mux_top_track_6.out
rlabel metal2 10258 40052 10258 40052 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17986 38522 17986 38522 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11086 31960 11086 31960 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9200 34986 9200 34986 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8786 39610 8786 39610 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9062 35258 9062 35258 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9016 45934 9016 45934 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 1380 45594 1380 45594 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 1518 48042 1518 48042 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 2668 50354 2668 50354 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 4002 52564 4002 52564 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
