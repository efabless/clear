magic
tech sky130A
magscale 1 2
timestamp 1681684910
<< viali >>
rect 3985 54281 4019 54315
rect 14105 54281 14139 54315
rect 14565 54281 14599 54315
rect 5825 54213 5859 54247
rect 8401 54213 8435 54247
rect 10977 54213 11011 54247
rect 14289 54213 14323 54247
rect 24133 54213 24167 54247
rect 2237 54145 2271 54179
rect 4629 54145 4663 54179
rect 7389 54145 7423 54179
rect 9965 54145 9999 54179
rect 11897 54145 11931 54179
rect 12357 54145 12391 54179
rect 14841 54145 14875 54179
rect 15485 54145 15519 54179
rect 15945 54145 15979 54179
rect 16865 54145 16899 54179
rect 17969 54145 18003 54179
rect 18889 54145 18923 54179
rect 19441 54145 19475 54179
rect 20545 54145 20579 54179
rect 22017 54145 22051 54179
rect 23121 54145 23155 54179
rect 24593 54145 24627 54179
rect 3249 54077 3283 54111
rect 12817 54077 12851 54111
rect 25145 54077 25179 54111
rect 21465 54009 21499 54043
rect 25421 54009 25455 54043
rect 3801 53941 3835 53975
rect 11713 53941 11747 53975
rect 16129 53941 16163 53975
rect 17509 53941 17543 53975
rect 18613 53941 18647 53975
rect 20085 53941 20119 53975
rect 21189 53941 21223 53975
rect 22661 53941 22695 53975
rect 23765 53941 23799 53975
rect 24777 53941 24811 53975
rect 18981 53737 19015 53771
rect 18797 53669 18831 53703
rect 23857 53669 23891 53703
rect 3249 53601 3283 53635
rect 6561 53601 6595 53635
rect 8401 53601 8435 53635
rect 11069 53601 11103 53635
rect 12725 53601 12759 53635
rect 18705 53601 18739 53635
rect 25145 53601 25179 53635
rect 2237 53533 2271 53567
rect 3985 53533 4019 53567
rect 5549 53533 5583 53567
rect 7297 53533 7331 53567
rect 10609 53533 10643 53567
rect 12449 53533 12483 53567
rect 14289 53533 14323 53567
rect 15393 53533 15427 53567
rect 16589 53533 16623 53567
rect 17693 53533 17727 53567
rect 19441 53533 19475 53567
rect 20545 53533 20579 53567
rect 21649 53533 21683 53567
rect 22753 53533 22787 53567
rect 24041 53533 24075 53567
rect 24685 53533 24719 53567
rect 24869 53533 24903 53567
rect 25329 53465 25363 53499
rect 4629 53397 4663 53431
rect 14933 53397 14967 53431
rect 16037 53397 16071 53431
rect 17233 53397 17267 53431
rect 18337 53397 18371 53431
rect 20085 53397 20119 53431
rect 21189 53397 21223 53431
rect 22293 53397 22327 53431
rect 23397 53397 23431 53431
rect 11621 53193 11655 53227
rect 17417 53193 17451 53227
rect 17693 53193 17727 53227
rect 3985 53125 4019 53159
rect 5825 53125 5859 53159
rect 9137 53125 9171 53159
rect 16037 53125 16071 53159
rect 19349 53125 19383 53159
rect 1685 53057 1719 53091
rect 2973 53057 3007 53091
rect 4721 53057 4755 53091
rect 6561 53057 6595 53091
rect 7941 53057 7975 53091
rect 9781 53057 9815 53091
rect 11897 53057 11931 53091
rect 13737 53057 13771 53091
rect 14841 53057 14875 53091
rect 16865 53057 16899 53091
rect 17877 53057 17911 53091
rect 18153 53057 18187 53091
rect 20085 53057 20119 53091
rect 20729 53057 20763 53091
rect 21281 53057 21315 53091
rect 22017 53057 22051 53091
rect 22753 53057 22787 53091
rect 23489 53057 23523 53091
rect 24317 53057 24351 53091
rect 25053 53057 25087 53091
rect 10333 52989 10367 53023
rect 12357 52989 12391 53023
rect 7205 52921 7239 52955
rect 16221 52921 16255 52955
rect 21465 52921 21499 52955
rect 22201 52921 22235 52955
rect 2329 52853 2363 52887
rect 14381 52853 14415 52887
rect 15485 52853 15519 52887
rect 17049 52853 17083 52887
rect 18797 52853 18831 52887
rect 19441 52853 19475 52887
rect 22937 52853 22971 52887
rect 23673 52853 23707 52887
rect 24501 52853 24535 52887
rect 25237 52853 25271 52887
rect 12633 52649 12667 52683
rect 14841 52649 14875 52683
rect 15209 52649 15243 52683
rect 16405 52649 16439 52683
rect 17049 52649 17083 52683
rect 22385 52649 22419 52683
rect 24041 52649 24075 52683
rect 24225 52649 24259 52683
rect 24777 52649 24811 52683
rect 17785 52581 17819 52615
rect 21833 52581 21867 52615
rect 23305 52581 23339 52615
rect 25237 52581 25271 52615
rect 3249 52513 3283 52547
rect 3985 52513 4019 52547
rect 4261 52513 4295 52547
rect 7757 52513 7791 52547
rect 11253 52513 11287 52547
rect 22845 52513 22879 52547
rect 2237 52445 2271 52479
rect 5457 52445 5491 52479
rect 6561 52445 6595 52479
rect 7297 52445 7331 52479
rect 10793 52445 10827 52479
rect 12817 52445 12851 52479
rect 13645 52445 13679 52479
rect 14289 52445 14323 52479
rect 15577 52445 15611 52479
rect 16865 52445 16899 52479
rect 17601 52445 17635 52479
rect 18429 52445 18463 52479
rect 19441 52445 19475 52479
rect 20177 52445 20211 52479
rect 20913 52445 20947 52479
rect 21649 52445 21683 52479
rect 22569 52445 22603 52479
rect 23489 52445 23523 52479
rect 23765 52445 23799 52479
rect 24593 52445 24627 52479
rect 25053 52445 25087 52479
rect 13461 52377 13495 52411
rect 14473 52309 14507 52343
rect 15761 52309 15795 52343
rect 18521 52309 18555 52343
rect 19625 52309 19659 52343
rect 20361 52309 20395 52343
rect 21097 52309 21131 52343
rect 7021 52105 7055 52139
rect 11713 52105 11747 52139
rect 12357 52105 12391 52139
rect 19901 52105 19935 52139
rect 21465 52105 21499 52139
rect 6929 52037 6963 52071
rect 13829 52037 13863 52071
rect 1685 51969 1719 52003
rect 2973 51969 3007 52003
rect 4813 51969 4847 52003
rect 8033 51969 8067 52003
rect 9689 51969 9723 52003
rect 11897 51969 11931 52003
rect 12541 51969 12575 52003
rect 14657 51969 14691 52003
rect 14933 51969 14967 52003
rect 16129 51969 16163 52003
rect 16405 51969 16439 52003
rect 17601 51969 17635 52003
rect 17877 51969 17911 52003
rect 19073 51969 19107 52003
rect 19349 51969 19383 52003
rect 20545 51969 20579 52003
rect 20821 51969 20855 52003
rect 23305 51969 23339 52003
rect 23581 51969 23615 52003
rect 24133 51969 24167 52003
rect 24409 51969 24443 52003
rect 24685 51969 24719 52003
rect 25053 51969 25087 52003
rect 3341 51901 3375 51935
rect 5089 51901 5123 51935
rect 8493 51901 8527 51935
rect 10149 51901 10183 51935
rect 14013 51833 14047 51867
rect 14473 51833 14507 51867
rect 15945 51833 15979 51867
rect 17417 51833 17451 51867
rect 23949 51833 23983 51867
rect 2329 51765 2363 51799
rect 18889 51765 18923 51799
rect 20361 51765 20395 51799
rect 23121 51765 23155 51799
rect 25237 51765 25271 51799
rect 10241 51561 10275 51595
rect 2881 51425 2915 51459
rect 7573 51425 7607 51459
rect 2237 51357 2271 51391
rect 3985 51357 4019 51391
rect 5457 51357 5491 51391
rect 6193 51357 6227 51391
rect 7113 51357 7147 51391
rect 10425 51357 10459 51391
rect 24777 51357 24811 51391
rect 25053 51357 25087 51391
rect 4629 51221 4663 51255
rect 25237 51221 25271 51255
rect 1593 51017 1627 51051
rect 6929 51017 6963 51051
rect 9597 50949 9631 50983
rect 1777 50881 1811 50915
rect 2513 50881 2547 50915
rect 4261 50881 4295 50915
rect 6837 50881 6871 50915
rect 7757 50881 7791 50915
rect 9413 50881 9447 50915
rect 24777 50881 24811 50915
rect 25053 50881 25087 50915
rect 2789 50813 2823 50847
rect 4629 50813 4663 50847
rect 7481 50813 7515 50847
rect 25237 50677 25271 50711
rect 6837 50473 6871 50507
rect 9229 50473 9263 50507
rect 3249 50337 3283 50371
rect 3985 50337 4019 50371
rect 5089 50337 5123 50371
rect 2237 50269 2271 50303
rect 4261 50269 4295 50303
rect 7021 50269 7055 50303
rect 9413 50269 9447 50303
rect 25421 50133 25455 50167
rect 6561 49929 6595 49963
rect 25145 49929 25179 49963
rect 3157 49861 3191 49895
rect 4261 49861 4295 49895
rect 6377 49861 6411 49895
rect 9321 49861 9355 49895
rect 1961 49793 1995 49827
rect 3985 49793 4019 49827
rect 9137 49793 9171 49827
rect 25329 49793 25363 49827
rect 6009 49725 6043 49759
rect 11621 49385 11655 49419
rect 2053 49249 2087 49283
rect 1777 49181 1811 49215
rect 11805 49181 11839 49215
rect 24869 49181 24903 49215
rect 25329 49181 25363 49215
rect 3341 49045 3375 49079
rect 25145 49045 25179 49079
rect 12725 48841 12759 48875
rect 12909 48705 12943 48739
rect 25513 48501 25547 48535
rect 17785 48229 17819 48263
rect 24869 48093 24903 48127
rect 25329 48093 25363 48127
rect 1685 48025 1719 48059
rect 2145 48025 2179 48059
rect 1777 47957 1811 47991
rect 25145 47957 25179 47991
rect 9137 47753 9171 47787
rect 17233 47753 17267 47787
rect 17325 47753 17359 47787
rect 18429 47753 18463 47787
rect 18521 47753 18555 47787
rect 19073 47753 19107 47787
rect 9321 47617 9355 47651
rect 24777 47617 24811 47651
rect 17417 47549 17451 47583
rect 18613 47549 18647 47583
rect 24501 47549 24535 47583
rect 16865 47413 16899 47447
rect 18061 47413 18095 47447
rect 9873 47209 9907 47243
rect 15932 47209 15966 47243
rect 19349 47209 19383 47243
rect 21649 47209 21683 47243
rect 18153 47141 18187 47175
rect 25145 47141 25179 47175
rect 10241 47073 10275 47107
rect 15669 47073 15703 47107
rect 17417 47073 17451 47107
rect 18613 47073 18647 47107
rect 18797 47073 18831 47107
rect 22569 47073 22603 47107
rect 18521 47005 18555 47039
rect 22385 47005 22419 47039
rect 22477 47005 22511 47039
rect 25329 47005 25363 47039
rect 10517 46937 10551 46971
rect 12265 46937 12299 46971
rect 14197 46937 14231 46971
rect 24869 46937 24903 46971
rect 11989 46869 12023 46903
rect 17693 46869 17727 46903
rect 22017 46869 22051 46903
rect 7205 46665 7239 46699
rect 10885 46665 10919 46699
rect 18613 46665 18647 46699
rect 20821 46665 20855 46699
rect 22661 46665 22695 46699
rect 22753 46665 22787 46699
rect 12633 46597 12667 46631
rect 21097 46597 21131 46631
rect 23489 46597 23523 46631
rect 7389 46529 7423 46563
rect 11069 46529 11103 46563
rect 24777 46529 24811 46563
rect 12357 46461 12391 46495
rect 14565 46461 14599 46495
rect 14841 46461 14875 46495
rect 16865 46461 16899 46495
rect 17141 46461 17175 46495
rect 19073 46461 19107 46495
rect 19349 46461 19383 46495
rect 22845 46461 22879 46495
rect 23305 46461 23339 46495
rect 24501 46461 24535 46495
rect 14105 46325 14139 46359
rect 16313 46325 16347 46359
rect 22293 46325 22327 46359
rect 8125 46121 8159 46155
rect 9137 46121 9171 46155
rect 10701 46121 10735 46155
rect 18705 46121 18739 46155
rect 19441 46121 19475 46155
rect 25421 46121 25455 46155
rect 10057 46053 10091 46087
rect 1869 45985 1903 46019
rect 11345 45985 11379 46019
rect 11897 45985 11931 46019
rect 12173 45985 12207 46019
rect 14105 45985 14139 46019
rect 20177 45985 20211 46019
rect 20361 45985 20395 46019
rect 21373 45985 21407 46019
rect 21557 45985 21591 46019
rect 1593 45917 1627 45951
rect 9321 45917 9355 45951
rect 10241 45917 10275 45951
rect 11069 45917 11103 45951
rect 20085 45917 20119 45951
rect 21281 45917 21315 45951
rect 21925 45917 21959 45951
rect 23213 45917 23247 45951
rect 23489 45917 23523 45951
rect 8033 45849 8067 45883
rect 8493 45849 8527 45883
rect 11161 45781 11195 45815
rect 13645 45781 13679 45815
rect 16405 45781 16439 45815
rect 19717 45781 19751 45815
rect 20913 45781 20947 45815
rect 24501 45781 24535 45815
rect 1409 45577 1443 45611
rect 20177 45577 20211 45611
rect 23765 45577 23799 45611
rect 8861 45509 8895 45543
rect 9229 45441 9263 45475
rect 9505 45373 9539 45407
rect 11529 45373 11563 45407
rect 14381 45373 14415 45407
rect 14657 45373 14691 45407
rect 18429 45373 18463 45407
rect 18705 45373 18739 45407
rect 22017 45373 22051 45407
rect 22293 45373 22327 45407
rect 24501 45373 24535 45407
rect 24777 45373 24811 45407
rect 10977 45305 11011 45339
rect 16405 45305 16439 45339
rect 11253 45237 11287 45271
rect 12173 45237 12207 45271
rect 16129 45237 16163 45271
rect 20545 45237 20579 45271
rect 24133 45237 24167 45271
rect 9321 45033 9355 45067
rect 11621 45033 11655 45067
rect 12449 45033 12483 45067
rect 13001 45033 13035 45067
rect 17141 45033 17175 45067
rect 7941 44965 7975 44999
rect 13553 44897 13587 44931
rect 21649 44897 21683 44931
rect 13369 44829 13403 44863
rect 15117 44829 15151 44863
rect 19533 44829 19567 44863
rect 22293 44829 22327 44863
rect 7757 44761 7791 44795
rect 9229 44761 9263 44795
rect 11161 44761 11195 44795
rect 11529 44761 11563 44795
rect 12357 44761 12391 44795
rect 15393 44761 15427 44795
rect 19809 44761 19843 44795
rect 22569 44761 22603 44795
rect 6469 44693 6503 44727
rect 7205 44693 7239 44727
rect 8309 44693 8343 44727
rect 9781 44693 9815 44727
rect 13461 44693 13495 44727
rect 16865 44693 16899 44727
rect 21281 44693 21315 44727
rect 24041 44693 24075 44727
rect 24409 44693 24443 44727
rect 25513 44693 25547 44727
rect 5825 44489 5859 44523
rect 6745 44489 6779 44523
rect 7481 44489 7515 44523
rect 8033 44489 8067 44523
rect 11069 44489 11103 44523
rect 11897 44489 11931 44523
rect 12265 44489 12299 44523
rect 18889 44489 18923 44523
rect 21281 44489 21315 44523
rect 21649 44489 21683 44523
rect 24041 44489 24075 44523
rect 9137 44421 9171 44455
rect 15393 44421 15427 44455
rect 6009 44353 6043 44387
rect 6653 44353 6687 44387
rect 7389 44353 7423 44387
rect 8217 44353 8251 44387
rect 8953 44353 8987 44387
rect 9413 44353 9447 44387
rect 10977 44353 11011 44387
rect 13185 44353 13219 44387
rect 24501 44353 24535 44387
rect 12357 44285 12391 44319
rect 12449 44285 12483 44319
rect 14933 44285 14967 44319
rect 16865 44285 16899 44319
rect 17141 44285 17175 44319
rect 19533 44285 19567 44319
rect 19809 44285 19843 44319
rect 22293 44285 22327 44319
rect 22569 44285 22603 44319
rect 24777 44285 24811 44319
rect 11621 44217 11655 44251
rect 13448 44149 13482 44183
rect 15209 44149 15243 44183
rect 18613 44149 18647 44183
rect 8401 43945 8435 43979
rect 11621 43945 11655 43979
rect 6929 43877 6963 43911
rect 9137 43809 9171 43843
rect 22477 43809 22511 43843
rect 22661 43809 22695 43843
rect 8585 43741 8619 43775
rect 6745 43673 6779 43707
rect 9413 43673 9447 43707
rect 11529 43673 11563 43707
rect 25421 43673 25455 43707
rect 1409 43605 1443 43639
rect 7205 43605 7239 43639
rect 10885 43605 10919 43639
rect 12081 43605 12115 43639
rect 17969 43605 18003 43639
rect 22017 43605 22051 43639
rect 22385 43605 22419 43639
rect 23029 43605 23063 43639
rect 24225 43605 24259 43639
rect 25329 43605 25363 43639
rect 7757 43401 7791 43435
rect 9505 43401 9539 43435
rect 10609 43401 10643 43435
rect 15025 43401 15059 43435
rect 17417 43401 17451 43435
rect 17509 43401 17543 43435
rect 20085 43401 20119 43435
rect 20453 43401 20487 43435
rect 21465 43401 21499 43435
rect 22477 43401 22511 43435
rect 8677 43333 8711 43367
rect 11069 43333 11103 43367
rect 12633 43333 12667 43367
rect 1593 43265 1627 43299
rect 7941 43265 7975 43299
rect 8493 43265 8527 43299
rect 9597 43265 9631 43299
rect 10517 43265 10551 43299
rect 12357 43265 12391 43299
rect 15117 43265 15151 43299
rect 22385 43265 22419 43299
rect 9689 43197 9723 43231
rect 15209 43197 15243 43231
rect 17601 43197 17635 43231
rect 18337 43197 18371 43231
rect 18613 43197 18647 43231
rect 22661 43197 22695 43231
rect 23581 43197 23615 43231
rect 23857 43197 23891 43231
rect 9137 43129 9171 43163
rect 2237 43061 2271 43095
rect 14105 43061 14139 43095
rect 14657 43061 14691 43095
rect 15761 43061 15795 43095
rect 16681 43061 16715 43095
rect 17049 43061 17083 43095
rect 21649 43061 21683 43095
rect 22017 43061 22051 43095
rect 25329 43061 25363 43095
rect 8585 42857 8619 42891
rect 8953 42857 8987 42891
rect 9229 42857 9263 42891
rect 12909 42857 12943 42891
rect 14289 42857 14323 42891
rect 19796 42857 19830 42891
rect 4997 42721 5031 42755
rect 9321 42721 9355 42755
rect 10793 42721 10827 42755
rect 14841 42721 14875 42755
rect 17785 42721 17819 42755
rect 18153 42721 18187 42755
rect 18429 42721 18463 42755
rect 19533 42721 19567 42755
rect 22293 42721 22327 42755
rect 22477 42721 22511 42755
rect 25329 42721 25363 42755
rect 1685 42653 1719 42687
rect 17601 42653 17635 42687
rect 23213 42653 23247 42687
rect 23489 42653 23523 42687
rect 1869 42585 1903 42619
rect 4813 42585 4847 42619
rect 5273 42585 5307 42619
rect 11069 42585 11103 42619
rect 15117 42585 15151 42619
rect 22201 42585 22235 42619
rect 8309 42517 8343 42551
rect 9505 42517 9539 42551
rect 10333 42517 10367 42551
rect 12541 42517 12575 42551
rect 16589 42517 16623 42551
rect 17141 42517 17175 42551
rect 17509 42517 17543 42551
rect 21281 42517 21315 42551
rect 21833 42517 21867 42551
rect 24501 42517 24535 42551
rect 4353 42313 4387 42347
rect 5089 42313 5123 42347
rect 6745 42313 6779 42347
rect 9689 42313 9723 42347
rect 11805 42313 11839 42347
rect 13001 42313 13035 42347
rect 15393 42313 15427 42347
rect 15853 42313 15887 42347
rect 16865 42313 16899 42347
rect 17233 42313 17267 42347
rect 18153 42313 18187 42347
rect 20269 42313 20303 42347
rect 20729 42313 20763 42347
rect 21373 42313 21407 42347
rect 25237 42313 25271 42347
rect 12265 42245 12299 42279
rect 15761 42245 15795 42279
rect 3893 42177 3927 42211
rect 4261 42177 4295 42211
rect 4997 42177 5031 42211
rect 6653 42177 6687 42211
rect 7481 42177 7515 42211
rect 10057 42177 10091 42211
rect 12173 42177 12207 42211
rect 13369 42177 13403 42211
rect 14197 42177 14231 42211
rect 18889 42177 18923 42211
rect 20637 42177 20671 42211
rect 22017 42177 22051 42211
rect 7757 42109 7791 42143
rect 10149 42109 10183 42143
rect 10241 42109 10275 42143
rect 12449 42109 12483 42143
rect 13461 42109 13495 42143
rect 13645 42109 13679 42143
rect 15945 42109 15979 42143
rect 17325 42109 17359 42143
rect 17509 42109 17543 42143
rect 17877 42109 17911 42143
rect 19625 42109 19659 42143
rect 20821 42109 20855 42143
rect 22845 42109 22879 42143
rect 23489 42109 23523 42143
rect 23765 42109 23799 42143
rect 18613 42041 18647 42075
rect 21557 42041 21591 42075
rect 5549 41973 5583 42007
rect 7113 41973 7147 42007
rect 9229 41973 9263 42007
rect 10701 41973 10735 42007
rect 16405 41973 16439 42007
rect 5181 41769 5215 41803
rect 7665 41769 7699 41803
rect 8125 41769 8159 41803
rect 10701 41769 10735 41803
rect 21189 41769 21223 41803
rect 8033 41701 8067 41735
rect 17325 41701 17359 41735
rect 22845 41701 22879 41735
rect 5917 41633 5951 41667
rect 10057 41633 10091 41667
rect 11253 41633 11287 41667
rect 12725 41633 12759 41667
rect 16773 41633 16807 41667
rect 18613 41633 18647 41667
rect 18797 41633 18831 41667
rect 19441 41633 19475 41667
rect 22293 41633 22327 41667
rect 23305 41633 23339 41667
rect 23397 41633 23431 41667
rect 9321 41565 9355 41599
rect 11989 41565 12023 41599
rect 16681 41565 16715 41599
rect 24501 41565 24535 41599
rect 25329 41565 25363 41599
rect 5089 41497 5123 41531
rect 6193 41497 6227 41531
rect 13185 41497 13219 41531
rect 19717 41497 19751 41531
rect 22109 41497 22143 41531
rect 23213 41497 23247 41531
rect 24225 41497 24259 41531
rect 1409 41429 1443 41463
rect 5641 41429 5675 41463
rect 11069 41429 11103 41463
rect 11161 41429 11195 41463
rect 16221 41429 16255 41463
rect 16589 41429 16623 41463
rect 18153 41429 18187 41463
rect 18521 41429 18555 41463
rect 21649 41429 21683 41463
rect 22017 41429 22051 41463
rect 24593 41429 24627 41463
rect 24869 41429 24903 41463
rect 25145 41429 25179 41463
rect 3341 41225 3375 41259
rect 8033 41225 8067 41259
rect 10977 41225 11011 41259
rect 11713 41225 11747 41259
rect 12173 41225 12207 41259
rect 15761 41225 15795 41259
rect 19901 41225 19935 41259
rect 22017 41225 22051 41259
rect 24685 41225 24719 41259
rect 18889 41157 18923 41191
rect 1593 41089 1627 41123
rect 3249 41089 3283 41123
rect 3709 41089 3743 41123
rect 8953 41089 8987 41123
rect 12081 41089 12115 41123
rect 13645 41089 13679 41123
rect 16865 41089 16899 41123
rect 19809 41089 19843 41123
rect 21097 41089 21131 41123
rect 25329 41089 25363 41123
rect 9229 41021 9263 41055
rect 12265 41021 12299 41055
rect 13921 41021 13955 41055
rect 17141 41021 17175 41055
rect 19993 41021 20027 41055
rect 21189 41021 21223 41055
rect 21281 41021 21315 41055
rect 22937 41021 22971 41055
rect 23213 41021 23247 41055
rect 15393 40953 15427 40987
rect 25145 40953 25179 40987
rect 2237 40885 2271 40919
rect 10701 40885 10735 40919
rect 18613 40885 18647 40919
rect 19165 40885 19199 40919
rect 19441 40885 19475 40919
rect 20729 40885 20763 40919
rect 7941 40681 7975 40715
rect 8493 40681 8527 40715
rect 10609 40681 10643 40715
rect 20913 40681 20947 40715
rect 22201 40681 22235 40715
rect 6469 40545 6503 40579
rect 9781 40545 9815 40579
rect 10241 40545 10275 40579
rect 11529 40545 11563 40579
rect 13277 40545 13311 40579
rect 14749 40545 14783 40579
rect 15853 40545 15887 40579
rect 17141 40545 17175 40579
rect 17233 40545 17267 40579
rect 21557 40545 21591 40579
rect 21925 40545 21959 40579
rect 22937 40545 22971 40579
rect 23121 40545 23155 40579
rect 1777 40477 1811 40511
rect 6193 40477 6227 40511
rect 8769 40477 8803 40511
rect 9689 40477 9723 40511
rect 13001 40477 13035 40511
rect 13093 40477 13127 40511
rect 13737 40477 13771 40511
rect 21281 40477 21315 40511
rect 22845 40477 22879 40511
rect 24685 40477 24719 40511
rect 25329 40477 25363 40511
rect 11069 40409 11103 40443
rect 11345 40409 11379 40443
rect 11805 40409 11839 40443
rect 14841 40409 14875 40443
rect 15669 40409 15703 40443
rect 17049 40409 17083 40443
rect 24041 40409 24075 40443
rect 24869 40409 24903 40443
rect 1593 40341 1627 40375
rect 8309 40341 8343 40375
rect 9229 40341 9263 40375
rect 9597 40341 9631 40375
rect 11713 40341 11747 40375
rect 12173 40341 12207 40375
rect 12633 40341 12667 40375
rect 15209 40341 15243 40375
rect 15577 40341 15611 40375
rect 16313 40341 16347 40375
rect 16681 40341 16715 40375
rect 20361 40341 20395 40375
rect 21373 40341 21407 40375
rect 22477 40341 22511 40375
rect 24225 40341 24259 40375
rect 24501 40341 24535 40375
rect 25145 40341 25179 40375
rect 7297 40137 7331 40171
rect 11529 40137 11563 40171
rect 12265 40137 12299 40171
rect 15025 40137 15059 40171
rect 15577 40137 15611 40171
rect 25237 40137 25271 40171
rect 7665 40069 7699 40103
rect 10517 40069 10551 40103
rect 15945 40069 15979 40103
rect 18613 40069 18647 40103
rect 20177 40069 20211 40103
rect 8493 40001 8527 40035
rect 12909 40001 12943 40035
rect 20269 40001 20303 40035
rect 21097 40001 21131 40035
rect 22293 40001 22327 40035
rect 22569 40001 22603 40035
rect 23489 40001 23523 40035
rect 7757 39933 7791 39967
rect 7849 39933 7883 39967
rect 8769 39933 8803 39967
rect 10977 39933 11011 39967
rect 13185 39933 13219 39967
rect 16037 39933 16071 39967
rect 16129 39933 16163 39967
rect 18705 39933 18739 39967
rect 18797 39933 18831 39967
rect 20453 39933 20487 39967
rect 23765 39933 23799 39967
rect 18245 39865 18279 39899
rect 19809 39865 19843 39899
rect 14657 39797 14691 39831
rect 16681 39797 16715 39831
rect 20913 39797 20947 39831
rect 6653 39593 6687 39627
rect 9781 39593 9815 39627
rect 11240 39593 11274 39627
rect 13093 39593 13127 39627
rect 15577 39593 15611 39627
rect 18797 39593 18831 39627
rect 19073 39593 19107 39627
rect 20453 39593 20487 39627
rect 21281 39593 21315 39627
rect 12725 39525 12759 39559
rect 13277 39525 13311 39559
rect 14381 39525 14415 39559
rect 4905 39457 4939 39491
rect 7113 39457 7147 39491
rect 10241 39457 10275 39491
rect 10333 39457 10367 39491
rect 10977 39457 11011 39491
rect 15025 39457 15059 39491
rect 16221 39457 16255 39491
rect 19901 39457 19935 39491
rect 20085 39457 20119 39491
rect 21925 39457 21959 39491
rect 22293 39457 22327 39491
rect 23305 39457 23339 39491
rect 25053 39457 25087 39491
rect 25237 39457 25271 39491
rect 23121 39389 23155 39423
rect 5181 39321 5215 39355
rect 6929 39321 6963 39355
rect 10149 39321 10183 39355
rect 14841 39321 14875 39355
rect 19809 39321 19843 39355
rect 21741 39321 21775 39355
rect 23029 39321 23063 39355
rect 23857 39321 23891 39355
rect 24961 39321 24995 39355
rect 9137 39253 9171 39287
rect 13829 39253 13863 39287
rect 14749 39253 14783 39287
rect 15945 39253 15979 39287
rect 16037 39253 16071 39287
rect 18613 39253 18647 39287
rect 19441 39253 19475 39287
rect 21649 39253 21683 39287
rect 22661 39253 22695 39287
rect 24593 39253 24627 39287
rect 7297 39049 7331 39083
rect 8217 39049 8251 39083
rect 9505 39049 9539 39083
rect 10793 39049 10827 39083
rect 14289 39049 14323 39083
rect 15301 39049 15335 39083
rect 19165 39049 19199 39083
rect 20729 39049 20763 39083
rect 24501 39049 24535 39083
rect 8677 38981 8711 39015
rect 10885 38981 10919 39015
rect 18337 38981 18371 39015
rect 19625 38981 19659 39015
rect 24133 38981 24167 39015
rect 8309 38913 8343 38947
rect 9597 38913 9631 38947
rect 12081 38913 12115 38947
rect 19533 38913 19567 38947
rect 24685 38913 24719 38947
rect 25329 38913 25363 38947
rect 9689 38845 9723 38879
rect 11069 38845 11103 38879
rect 12357 38845 12391 38879
rect 15393 38845 15427 38879
rect 15577 38845 15611 38879
rect 16865 38845 16899 38879
rect 18429 38845 18463 38879
rect 18613 38845 18647 38879
rect 19717 38845 19751 38879
rect 20821 38845 20855 38879
rect 21005 38845 21039 38879
rect 22116 38845 22150 38879
rect 22385 38845 22419 38879
rect 8585 38777 8619 38811
rect 10425 38777 10459 38811
rect 14933 38777 14967 38811
rect 1409 38709 1443 38743
rect 9137 38709 9171 38743
rect 11529 38709 11563 38743
rect 13829 38709 13863 38743
rect 16037 38709 16071 38743
rect 17969 38709 18003 38743
rect 20361 38709 20395 38743
rect 23857 38709 23891 38743
rect 25145 38709 25179 38743
rect 7849 38505 7883 38539
rect 10425 38505 10459 38539
rect 14289 38505 14323 38539
rect 19441 38505 19475 38539
rect 11897 38437 11931 38471
rect 18153 38437 18187 38471
rect 5733 38369 5767 38403
rect 7205 38369 7239 38403
rect 8493 38369 8527 38403
rect 9689 38369 9723 38403
rect 9781 38369 9815 38403
rect 10977 38369 11011 38403
rect 12357 38369 12391 38403
rect 12449 38369 12483 38403
rect 13277 38369 13311 38403
rect 13921 38369 13955 38403
rect 14841 38369 14875 38403
rect 18705 38369 18739 38403
rect 19993 38369 20027 38403
rect 21097 38369 21131 38403
rect 21281 38369 21315 38403
rect 22477 38369 22511 38403
rect 22661 38369 22695 38403
rect 23765 38369 23799 38403
rect 25053 38369 25087 38403
rect 25145 38369 25179 38403
rect 1593 38301 1627 38335
rect 5457 38301 5491 38335
rect 8217 38301 8251 38335
rect 14749 38301 14783 38335
rect 15945 38301 15979 38335
rect 18521 38301 18555 38335
rect 18613 38301 18647 38335
rect 19901 38301 19935 38335
rect 21649 38301 21683 38335
rect 16221 38233 16255 38267
rect 19809 38233 19843 38267
rect 21005 38233 21039 38267
rect 22385 38233 22419 38267
rect 2237 38165 2271 38199
rect 7481 38165 7515 38199
rect 8309 38165 8343 38199
rect 9229 38165 9263 38199
rect 9597 38165 9631 38199
rect 10793 38165 10827 38199
rect 10885 38165 10919 38199
rect 12265 38165 12299 38199
rect 12909 38165 12943 38199
rect 14657 38165 14691 38199
rect 17693 38165 17727 38199
rect 20637 38165 20671 38199
rect 22017 38165 22051 38199
rect 23213 38165 23247 38199
rect 23581 38165 23615 38199
rect 23673 38165 23707 38199
rect 24593 38165 24627 38199
rect 24961 38165 24995 38199
rect 5273 37961 5307 37995
rect 5733 37961 5767 37995
rect 10057 37961 10091 37995
rect 11713 37961 11747 37995
rect 14105 37961 14139 37995
rect 16405 37961 16439 37995
rect 17233 37961 17267 37995
rect 18061 37961 18095 37995
rect 18337 37961 18371 37995
rect 18981 37961 19015 37995
rect 19441 37961 19475 37995
rect 20729 37961 20763 37995
rect 21557 37961 21591 37995
rect 22017 37961 22051 37995
rect 6837 37893 6871 37927
rect 8585 37893 8619 37927
rect 11253 37893 11287 37927
rect 12817 37893 12851 37927
rect 22477 37893 22511 37927
rect 1777 37825 1811 37859
rect 5641 37825 5675 37859
rect 9137 37825 9171 37859
rect 9413 37825 9447 37859
rect 10425 37825 10459 37859
rect 10517 37825 10551 37859
rect 12725 37825 12759 37859
rect 14381 37825 14415 37859
rect 15393 37825 15427 37859
rect 15485 37825 15519 37859
rect 18429 37825 18463 37859
rect 19349 37825 19383 37859
rect 20637 37825 20671 37859
rect 21281 37825 21315 37859
rect 22385 37825 22419 37859
rect 23213 37825 23247 37859
rect 5825 37757 5859 37791
rect 6561 37757 6595 37791
rect 10701 37757 10735 37791
rect 13001 37757 13035 37791
rect 13553 37757 13587 37791
rect 15669 37757 15703 37791
rect 17325 37757 17359 37791
rect 17509 37757 17543 37791
rect 19625 37757 19659 37791
rect 20913 37757 20947 37791
rect 22569 37757 22603 37791
rect 23581 37757 23615 37791
rect 23857 37757 23891 37791
rect 25329 37757 25363 37791
rect 17877 37689 17911 37723
rect 1593 37621 1627 37655
rect 8861 37621 8895 37655
rect 12357 37621 12391 37655
rect 15025 37621 15059 37655
rect 16129 37621 16163 37655
rect 16865 37621 16899 37655
rect 18705 37621 18739 37655
rect 20269 37621 20303 37655
rect 23029 37621 23063 37655
rect 8585 37417 8619 37451
rect 10425 37417 10459 37451
rect 10885 37417 10919 37451
rect 14657 37417 14691 37451
rect 23949 37417 23983 37451
rect 24685 37417 24719 37451
rect 14197 37349 14231 37383
rect 20637 37349 20671 37383
rect 7113 37281 7147 37315
rect 11805 37281 11839 37315
rect 12449 37281 12483 37315
rect 13369 37281 13403 37315
rect 13461 37281 13495 37315
rect 15485 37281 15519 37315
rect 16589 37281 16623 37315
rect 16681 37281 16715 37315
rect 17877 37281 17911 37315
rect 19073 37281 19107 37315
rect 24593 37281 24627 37315
rect 6837 37213 6871 37247
rect 9873 37213 9907 37247
rect 11621 37213 11655 37247
rect 13277 37213 13311 37247
rect 16497 37213 16531 37247
rect 17785 37213 17819 37247
rect 21097 37213 21131 37247
rect 21465 37213 21499 37247
rect 25329 37213 25363 37247
rect 9137 37145 9171 37179
rect 11713 37145 11747 37179
rect 15393 37145 15427 37179
rect 17693 37145 17727 37179
rect 19441 37145 19475 37179
rect 20177 37145 20211 37179
rect 22293 37145 22327 37179
rect 24225 37145 24259 37179
rect 10609 37077 10643 37111
rect 11253 37077 11287 37111
rect 12633 37077 12667 37111
rect 12909 37077 12943 37111
rect 14473 37077 14507 37111
rect 14933 37077 14967 37111
rect 15301 37077 15335 37111
rect 16129 37077 16163 37111
rect 17325 37077 17359 37111
rect 18521 37077 18555 37111
rect 23857 37077 23891 37111
rect 25145 37077 25179 37111
rect 7481 36873 7515 36907
rect 7941 36873 7975 36907
rect 9045 36873 9079 36907
rect 12081 36873 12115 36907
rect 12541 36873 12575 36907
rect 13829 36873 13863 36907
rect 15025 36873 15059 36907
rect 15577 36873 15611 36907
rect 17049 36873 17083 36907
rect 17417 36873 17451 36907
rect 20361 36873 20395 36907
rect 6009 36805 6043 36839
rect 10241 36805 10275 36839
rect 11529 36805 11563 36839
rect 3985 36737 4019 36771
rect 7849 36737 7883 36771
rect 9413 36737 9447 36771
rect 13737 36737 13771 36771
rect 14933 36737 14967 36771
rect 16681 36737 16715 36771
rect 17509 36737 17543 36771
rect 20453 36737 20487 36771
rect 21005 36737 21039 36771
rect 25329 36737 25363 36771
rect 4261 36669 4295 36703
rect 5733 36669 5767 36703
rect 8033 36669 8067 36703
rect 9505 36669 9539 36703
rect 9597 36669 9631 36703
rect 10977 36669 11011 36703
rect 11897 36669 11931 36703
rect 12633 36669 12667 36703
rect 12817 36669 12851 36703
rect 14013 36669 14047 36703
rect 15209 36669 15243 36703
rect 15853 36669 15887 36703
rect 17693 36669 17727 36703
rect 20545 36669 20579 36703
rect 22845 36669 22879 36703
rect 23121 36669 23155 36703
rect 24593 36669 24627 36703
rect 19349 36601 19383 36635
rect 25145 36601 25179 36635
rect 1501 36533 1535 36567
rect 8677 36533 8711 36567
rect 12173 36533 12207 36567
rect 13369 36533 13403 36567
rect 14565 36533 14599 36567
rect 19993 36533 20027 36567
rect 7665 36329 7699 36363
rect 9137 36329 9171 36363
rect 12449 36329 12483 36363
rect 12725 36329 12759 36363
rect 14289 36329 14323 36363
rect 16129 36329 16163 36363
rect 19441 36329 19475 36363
rect 12173 36261 12207 36295
rect 13829 36261 13863 36295
rect 19073 36261 19107 36295
rect 23305 36261 23339 36295
rect 8217 36193 8251 36227
rect 9689 36193 9723 36227
rect 13185 36193 13219 36227
rect 13369 36193 13403 36227
rect 14749 36193 14783 36227
rect 14933 36193 14967 36227
rect 16773 36193 16807 36227
rect 19993 36193 20027 36227
rect 21281 36193 21315 36227
rect 21373 36193 21407 36227
rect 23765 36193 23799 36227
rect 23949 36193 23983 36227
rect 1593 36125 1627 36159
rect 9597 36125 9631 36159
rect 16589 36125 16623 36159
rect 21189 36125 21223 36159
rect 24869 36125 24903 36159
rect 25329 36125 25363 36159
rect 8125 36057 8159 36091
rect 15761 36057 15795 36091
rect 16497 36057 16531 36091
rect 17325 36057 17359 36091
rect 19901 36057 19935 36091
rect 2237 35989 2271 36023
rect 8033 35989 8067 36023
rect 9505 35989 9539 36023
rect 13093 35989 13127 36023
rect 14657 35989 14691 36023
rect 19809 35989 19843 36023
rect 20821 35989 20855 36023
rect 23673 35989 23707 36023
rect 25145 35989 25179 36023
rect 6009 35785 6043 35819
rect 13921 35785 13955 35819
rect 14473 35785 14507 35819
rect 20177 35785 20211 35819
rect 24869 35785 24903 35819
rect 17877 35717 17911 35751
rect 20269 35717 20303 35751
rect 1777 35649 1811 35683
rect 4261 35649 4295 35683
rect 6377 35649 6411 35683
rect 23121 35649 23155 35683
rect 4537 35581 4571 35615
rect 8125 35581 8159 35615
rect 8401 35581 8435 35615
rect 11713 35581 11747 35615
rect 11989 35581 12023 35615
rect 17601 35581 17635 35615
rect 19349 35581 19383 35615
rect 20361 35581 20395 35615
rect 22477 35581 22511 35615
rect 23397 35581 23431 35615
rect 1593 35445 1627 35479
rect 9873 35445 9907 35479
rect 10241 35445 10275 35479
rect 13461 35445 13495 35479
rect 13829 35445 13863 35479
rect 19809 35445 19843 35479
rect 20821 35445 20855 35479
rect 25237 35445 25271 35479
rect 25421 35445 25455 35479
rect 7849 35241 7883 35275
rect 9321 35241 9355 35275
rect 13001 35241 13035 35275
rect 17141 35241 17175 35275
rect 17509 35241 17543 35275
rect 21649 35241 21683 35275
rect 21741 35173 21775 35207
rect 6101 35105 6135 35139
rect 6377 35105 6411 35139
rect 9873 35105 9907 35139
rect 13553 35105 13587 35139
rect 15393 35105 15427 35139
rect 19441 35105 19475 35139
rect 13461 35037 13495 35071
rect 22293 35037 22327 35071
rect 25329 35037 25363 35071
rect 9689 34969 9723 35003
rect 9781 34969 9815 35003
rect 15669 34969 15703 35003
rect 19717 34969 19751 35003
rect 22569 34969 22603 35003
rect 8125 34901 8159 34935
rect 13369 34901 13403 34935
rect 21189 34901 21223 34935
rect 24041 34901 24075 34935
rect 24409 34901 24443 34935
rect 25145 34901 25179 34935
rect 8309 34697 8343 34731
rect 10609 34697 10643 34731
rect 15945 34697 15979 34731
rect 20269 34697 20303 34731
rect 20729 34697 20763 34731
rect 21097 34697 21131 34731
rect 22385 34697 22419 34731
rect 23213 34697 23247 34731
rect 24409 34697 24443 34731
rect 6837 34629 6871 34663
rect 11989 34629 12023 34663
rect 16037 34629 16071 34663
rect 23581 34629 23615 34663
rect 6561 34561 6595 34595
rect 8861 34561 8895 34595
rect 21189 34561 21223 34595
rect 24593 34561 24627 34595
rect 25329 34561 25363 34595
rect 11713 34493 11747 34527
rect 13461 34493 13495 34527
rect 16129 34493 16163 34527
rect 21281 34493 21315 34527
rect 22477 34493 22511 34527
rect 22661 34493 22695 34527
rect 23673 34493 23707 34527
rect 23857 34493 23891 34527
rect 25145 34425 25179 34459
rect 9124 34357 9158 34391
rect 10977 34357 11011 34391
rect 13829 34357 13863 34391
rect 15577 34357 15611 34391
rect 22017 34357 22051 34391
rect 7573 34153 7607 34187
rect 7757 34153 7791 34187
rect 9137 34153 9171 34187
rect 12173 34153 12207 34187
rect 17693 34153 17727 34187
rect 18061 34153 18095 34187
rect 20545 34153 20579 34187
rect 23305 34153 23339 34187
rect 25329 34153 25363 34187
rect 8493 34085 8527 34119
rect 19441 34085 19475 34119
rect 22293 34085 22327 34119
rect 5549 34017 5583 34051
rect 7297 34017 7331 34051
rect 9689 34017 9723 34051
rect 10701 34017 10735 34051
rect 13461 34017 13495 34051
rect 13553 34017 13587 34051
rect 15945 34017 15979 34051
rect 19073 34017 19107 34051
rect 19993 34017 20027 34051
rect 21649 34017 21683 34051
rect 22753 34017 22787 34051
rect 22937 34017 22971 34051
rect 10425 33949 10459 33983
rect 12541 33949 12575 33983
rect 19809 33949 19843 33983
rect 21557 33949 21591 33983
rect 24777 33949 24811 33983
rect 5825 33881 5859 33915
rect 9505 33881 9539 33915
rect 16221 33881 16255 33915
rect 19901 33881 19935 33915
rect 25421 33881 25455 33915
rect 1409 33813 1443 33847
rect 9597 33813 9631 33847
rect 13001 33813 13035 33847
rect 13369 33813 13403 33847
rect 14105 33813 14139 33847
rect 20637 33813 20671 33847
rect 21097 33813 21131 33847
rect 21465 33813 21499 33847
rect 22661 33813 22695 33847
rect 24593 33813 24627 33847
rect 7113 33609 7147 33643
rect 10425 33609 10459 33643
rect 10885 33609 10919 33643
rect 12909 33609 12943 33643
rect 13369 33609 13403 33643
rect 16221 33609 16255 33643
rect 19809 33609 19843 33643
rect 22661 33609 22695 33643
rect 25237 33609 25271 33643
rect 12817 33541 12851 33575
rect 1593 33473 1627 33507
rect 10793 33473 10827 33507
rect 13277 33473 13311 33507
rect 14105 33473 14139 33507
rect 18061 33473 18095 33507
rect 20637 33473 20671 33507
rect 20729 33473 20763 33507
rect 23489 33473 23523 33507
rect 5365 33405 5399 33439
rect 9781 33405 9815 33439
rect 10977 33405 11011 33439
rect 13461 33405 13495 33439
rect 14381 33405 14415 33439
rect 18337 33405 18371 33439
rect 20821 33405 20855 33439
rect 22017 33405 22051 33439
rect 23765 33405 23799 33439
rect 20269 33337 20303 33371
rect 2237 33269 2271 33303
rect 12541 33269 12575 33303
rect 15853 33269 15887 33303
rect 21373 33269 21407 33303
rect 7481 33065 7515 33099
rect 9413 33065 9447 33099
rect 10609 33065 10643 33099
rect 11161 33065 11195 33099
rect 12265 33065 12299 33099
rect 19441 33065 19475 33099
rect 19809 33065 19843 33099
rect 25145 33065 25179 33099
rect 7021 32997 7055 33031
rect 21005 32997 21039 33031
rect 22937 32997 22971 33031
rect 5273 32929 5307 32963
rect 8125 32929 8159 32963
rect 10057 32929 10091 32963
rect 10885 32929 10919 32963
rect 11621 32929 11655 32963
rect 11805 32929 11839 32963
rect 14749 32929 14783 32963
rect 14841 32929 14875 32963
rect 16681 32929 16715 32963
rect 20269 32929 20303 32963
rect 20453 32929 20487 32963
rect 21557 32929 21591 32963
rect 1777 32861 1811 32895
rect 9781 32861 9815 32895
rect 11529 32861 11563 32895
rect 15761 32861 15795 32895
rect 16589 32861 16623 32895
rect 17325 32861 17359 32895
rect 20177 32861 20211 32895
rect 22385 32857 22419 32891
rect 24869 32861 24903 32895
rect 25329 32861 25363 32895
rect 5549 32793 5583 32827
rect 7941 32793 7975 32827
rect 17233 32793 17267 32827
rect 1593 32725 1627 32759
rect 7849 32725 7883 32759
rect 9873 32725 9907 32759
rect 14289 32725 14323 32759
rect 14657 32725 14691 32759
rect 16129 32725 16163 32759
rect 16497 32725 16531 32759
rect 17969 32725 18003 32759
rect 21373 32725 21407 32759
rect 21465 32725 21499 32759
rect 22201 32725 22235 32759
rect 22753 32725 22787 32759
rect 4629 32521 4663 32555
rect 4997 32521 5031 32555
rect 5365 32521 5399 32555
rect 6929 32521 6963 32555
rect 11989 32521 12023 32555
rect 18429 32521 18463 32555
rect 18521 32521 18555 32555
rect 19073 32521 19107 32555
rect 21189 32521 21223 32555
rect 21925 32521 21959 32555
rect 5457 32453 5491 32487
rect 17233 32453 17267 32487
rect 7573 32385 7607 32419
rect 12357 32385 12391 32419
rect 13185 32385 13219 32419
rect 14565 32385 14599 32419
rect 20269 32385 20303 32419
rect 21097 32385 21131 32419
rect 22385 32385 22419 32419
rect 23029 32385 23063 32419
rect 24869 32385 24903 32419
rect 25329 32385 25363 32419
rect 5549 32317 5583 32351
rect 7849 32317 7883 32351
rect 9873 32317 9907 32351
rect 11713 32317 11747 32351
rect 12449 32317 12483 32351
rect 12541 32317 12575 32351
rect 14841 32317 14875 32351
rect 16313 32317 16347 32351
rect 17325 32317 17359 32351
rect 17509 32317 17543 32351
rect 18613 32317 18647 32351
rect 19257 32317 19291 32351
rect 21373 32317 21407 32351
rect 23305 32317 23339 32351
rect 25145 32249 25179 32283
rect 9321 32181 9355 32215
rect 10425 32181 10459 32215
rect 16865 32181 16899 32215
rect 18061 32181 18095 32215
rect 20085 32181 20119 32215
rect 20729 32181 20763 32215
rect 22201 32181 22235 32215
rect 22845 32181 22879 32215
rect 7941 31977 7975 32011
rect 8401 31977 8435 32011
rect 8585 31977 8619 32011
rect 11161 31977 11195 32011
rect 16405 31977 16439 32011
rect 18061 31977 18095 32011
rect 13645 31909 13679 31943
rect 13921 31909 13955 31943
rect 14289 31909 14323 31943
rect 19441 31909 19475 31943
rect 20637 31909 20671 31943
rect 21925 31909 21959 31943
rect 25145 31909 25179 31943
rect 6193 31841 6227 31875
rect 6469 31841 6503 31875
rect 9689 31841 9723 31875
rect 14749 31841 14783 31875
rect 14841 31841 14875 31875
rect 16957 31841 16991 31875
rect 19993 31841 20027 31875
rect 21189 31841 21223 31875
rect 22385 31841 22419 31875
rect 22569 31841 22603 31875
rect 9402 31773 9436 31807
rect 19901 31773 19935 31807
rect 21097 31773 21131 31807
rect 24041 31773 24075 31807
rect 24869 31773 24903 31807
rect 25329 31773 25363 31807
rect 16865 31705 16899 31739
rect 18429 31705 18463 31739
rect 19809 31705 19843 31739
rect 21005 31705 21039 31739
rect 22293 31705 22327 31739
rect 9137 31637 9171 31671
rect 11529 31637 11563 31671
rect 14657 31637 14691 31671
rect 16773 31637 16807 31671
rect 18245 31637 18279 31671
rect 7481 31433 7515 31467
rect 8677 31433 8711 31467
rect 9045 31433 9079 31467
rect 14657 31433 14691 31467
rect 18337 31433 18371 31467
rect 19533 31433 19567 31467
rect 21557 31433 21591 31467
rect 25145 31433 25179 31467
rect 19901 31365 19935 31399
rect 20545 31365 20579 31399
rect 22477 31365 22511 31399
rect 1777 31297 1811 31331
rect 7849 31297 7883 31331
rect 15025 31297 15059 31331
rect 17509 31297 17543 31331
rect 17601 31297 17635 31331
rect 18705 31297 18739 31331
rect 20729 31297 20763 31331
rect 24593 31297 24627 31331
rect 25329 31297 25363 31331
rect 2053 31229 2087 31263
rect 7941 31229 7975 31263
rect 8125 31229 8159 31263
rect 9137 31229 9171 31263
rect 9229 31229 9263 31263
rect 9689 31229 9723 31263
rect 12909 31229 12943 31263
rect 13185 31229 13219 31263
rect 17693 31229 17727 31263
rect 18797 31229 18831 31263
rect 18889 31229 18923 31263
rect 19993 31229 20027 31263
rect 20177 31229 20211 31263
rect 22201 31229 22235 31263
rect 7205 31161 7239 31195
rect 16773 31093 16807 31127
rect 17141 31093 17175 31127
rect 23949 31093 23983 31127
rect 24409 31093 24443 31127
rect 12817 30889 12851 30923
rect 24869 30889 24903 30923
rect 11713 30821 11747 30855
rect 15945 30821 15979 30855
rect 18245 30821 18279 30855
rect 20453 30821 20487 30855
rect 25145 30821 25179 30855
rect 4077 30753 4111 30787
rect 4629 30753 4663 30787
rect 7941 30753 7975 30787
rect 9597 30753 9631 30787
rect 9873 30753 9907 30787
rect 12541 30753 12575 30787
rect 13369 30753 13403 30787
rect 16221 30753 16255 30787
rect 16497 30753 16531 30787
rect 19901 30753 19935 30787
rect 19993 30753 20027 30787
rect 22569 30753 22603 30787
rect 12265 30685 12299 30719
rect 13185 30685 13219 30719
rect 19809 30685 19843 30719
rect 22477 30685 22511 30719
rect 23029 30685 23063 30719
rect 23857 30685 23891 30719
rect 25329 30685 25363 30719
rect 4169 30617 4203 30651
rect 13277 30617 13311 30651
rect 13921 30617 13955 30651
rect 22385 30617 22419 30651
rect 8585 30549 8619 30583
rect 11345 30549 11379 30583
rect 17969 30549 18003 30583
rect 19441 30549 19475 30583
rect 22017 30549 22051 30583
rect 23673 30549 23707 30583
rect 10057 30345 10091 30379
rect 10885 30345 10919 30379
rect 8953 30277 8987 30311
rect 23673 30277 23707 30311
rect 25421 30277 25455 30311
rect 10793 30209 10827 30243
rect 11713 30209 11747 30243
rect 14473 30209 14507 30243
rect 17969 30209 18003 30243
rect 18613 30209 18647 30243
rect 18797 30209 18831 30243
rect 19625 30209 19659 30243
rect 23397 30209 23431 30243
rect 11069 30141 11103 30175
rect 16221 30141 16255 30175
rect 16957 30141 16991 30175
rect 18061 30141 18095 30175
rect 18245 30141 18279 30175
rect 25145 30141 25179 30175
rect 10425 30005 10459 30039
rect 12265 30005 12299 30039
rect 12541 30005 12575 30039
rect 14736 30005 14770 30039
rect 17601 30005 17635 30039
rect 19441 30005 19475 30039
rect 7297 29801 7331 29835
rect 7849 29801 7883 29835
rect 9505 29801 9539 29835
rect 16037 29801 16071 29835
rect 21557 29801 21591 29835
rect 12633 29733 12667 29767
rect 22937 29733 22971 29767
rect 4353 29665 4387 29699
rect 8401 29665 8435 29699
rect 9229 29665 9263 29699
rect 10057 29665 10091 29699
rect 11989 29665 12023 29699
rect 13185 29665 13219 29699
rect 17509 29665 17543 29699
rect 18797 29665 18831 29699
rect 20085 29665 20119 29699
rect 20269 29665 20303 29699
rect 22201 29665 22235 29699
rect 23397 29665 23431 29699
rect 23581 29665 23615 29699
rect 13001 29597 13035 29631
rect 17417 29597 17451 29631
rect 19993 29597 20027 29631
rect 21925 29597 21959 29631
rect 25329 29597 25363 29631
rect 4445 29529 4479 29563
rect 5365 29529 5399 29563
rect 7481 29529 7515 29563
rect 8309 29529 8343 29563
rect 9873 29529 9907 29563
rect 11805 29529 11839 29563
rect 13093 29529 13127 29563
rect 14749 29529 14783 29563
rect 17325 29529 17359 29563
rect 18613 29529 18647 29563
rect 8217 29461 8251 29495
rect 9045 29461 9079 29495
rect 9965 29461 9999 29495
rect 11437 29461 11471 29495
rect 11897 29461 11931 29495
rect 13737 29461 13771 29495
rect 16957 29461 16991 29495
rect 18153 29461 18187 29495
rect 18521 29461 18555 29495
rect 19625 29461 19659 29495
rect 20913 29461 20947 29495
rect 22017 29461 22051 29495
rect 23305 29461 23339 29495
rect 25145 29461 25179 29495
rect 12909 29257 12943 29291
rect 14197 29257 14231 29291
rect 16037 29257 16071 29291
rect 17233 29257 17267 29291
rect 17325 29257 17359 29291
rect 17969 29257 18003 29291
rect 22385 29257 22419 29291
rect 23949 29257 23983 29291
rect 25329 29257 25363 29291
rect 25513 29257 25547 29291
rect 9781 29189 9815 29223
rect 16221 29189 16255 29223
rect 21097 29189 21131 29223
rect 21557 29189 21591 29223
rect 22477 29189 22511 29223
rect 24685 29189 24719 29223
rect 13001 29121 13035 29155
rect 14105 29121 14139 29155
rect 15301 29121 15335 29155
rect 20453 29121 20487 29155
rect 23673 29121 23707 29155
rect 24133 29121 24167 29155
rect 7757 29053 7791 29087
rect 9505 29053 9539 29087
rect 13093 29053 13127 29087
rect 14381 29053 14415 29087
rect 15393 29053 15427 29087
rect 15485 29053 15519 29087
rect 17417 29053 17451 29087
rect 19717 29053 19751 29087
rect 20545 29053 20579 29087
rect 20637 29053 20671 29087
rect 22661 29053 22695 29087
rect 12541 28985 12575 29019
rect 13737 28985 13771 29019
rect 14933 28985 14967 29019
rect 16405 28985 16439 29019
rect 18153 28985 18187 29019
rect 20085 28985 20119 29019
rect 22017 28985 22051 29019
rect 24869 28985 24903 29019
rect 8020 28917 8054 28951
rect 16865 28917 16899 28951
rect 8677 28713 8711 28747
rect 12817 28713 12851 28747
rect 21189 28713 21223 28747
rect 8309 28645 8343 28679
rect 23857 28645 23891 28679
rect 2053 28577 2087 28611
rect 4353 28577 4387 28611
rect 5181 28577 5215 28611
rect 6561 28577 6595 28611
rect 6837 28577 6871 28611
rect 10885 28577 10919 28611
rect 13369 28577 13403 28611
rect 14841 28577 14875 28611
rect 16221 28577 16255 28611
rect 17693 28577 17727 28611
rect 17785 28577 17819 28611
rect 19441 28577 19475 28611
rect 1777 28509 1811 28543
rect 10609 28509 10643 28543
rect 14657 28509 14691 28543
rect 16037 28509 16071 28543
rect 17601 28509 17635 28543
rect 24041 28509 24075 28543
rect 24777 28509 24811 28543
rect 4445 28441 4479 28475
rect 16129 28441 16163 28475
rect 19717 28441 19751 28475
rect 21465 28441 21499 28475
rect 12357 28373 12391 28407
rect 13185 28373 13219 28407
rect 13277 28373 13311 28407
rect 13921 28373 13955 28407
rect 14289 28373 14323 28407
rect 14749 28373 14783 28407
rect 15301 28373 15335 28407
rect 15669 28373 15703 28407
rect 16773 28373 16807 28407
rect 17233 28373 17267 28407
rect 24593 28373 24627 28407
rect 2053 28169 2087 28203
rect 3755 28169 3789 28203
rect 12633 28169 12667 28203
rect 13369 28169 13403 28203
rect 15945 28169 15979 28203
rect 16865 28169 16899 28203
rect 18337 28169 18371 28203
rect 23765 28169 23799 28203
rect 16681 28101 16715 28135
rect 24685 28101 24719 28135
rect 2237 28033 2271 28067
rect 3652 28033 3686 28067
rect 13185 28033 13219 28067
rect 18245 28033 18279 28067
rect 19441 28033 19475 28067
rect 22017 28033 22051 28067
rect 8309 27965 8343 27999
rect 8585 27965 8619 27999
rect 16037 27965 16071 27999
rect 16221 27965 16255 27999
rect 18521 27965 18555 27999
rect 19533 27965 19567 27999
rect 19717 27965 19751 27999
rect 22293 27965 22327 27999
rect 10057 27897 10091 27931
rect 17049 27897 17083 27931
rect 24869 27897 24903 27931
rect 10425 27829 10459 27863
rect 15117 27829 15151 27863
rect 15577 27829 15611 27863
rect 17509 27829 17543 27863
rect 17877 27829 17911 27863
rect 19073 27829 19107 27863
rect 20085 27829 20119 27863
rect 24133 27829 24167 27863
rect 6456 27625 6490 27659
rect 13185 27625 13219 27659
rect 18705 27625 18739 27659
rect 24225 27625 24259 27659
rect 7941 27557 7975 27591
rect 8309 27557 8343 27591
rect 8401 27557 8435 27591
rect 18153 27557 18187 27591
rect 6193 27489 6227 27523
rect 15669 27489 15703 27523
rect 16405 27489 16439 27523
rect 20545 27489 20579 27523
rect 20637 27489 20671 27523
rect 21925 27489 21959 27523
rect 11161 27421 11195 27455
rect 15485 27421 15519 27455
rect 18337 27421 18371 27455
rect 24685 27421 24719 27455
rect 11437 27353 11471 27387
rect 15577 27353 15611 27387
rect 16129 27353 16163 27387
rect 19717 27353 19751 27387
rect 20453 27353 20487 27387
rect 22201 27353 22235 27387
rect 24869 27353 24903 27387
rect 12909 27285 12943 27319
rect 15117 27285 15151 27319
rect 18889 27285 18923 27319
rect 20085 27285 20119 27319
rect 23673 27285 23707 27319
rect 25237 27285 25271 27319
rect 3203 27081 3237 27115
rect 11805 27081 11839 27115
rect 15209 27081 15243 27115
rect 17601 27081 17635 27115
rect 19993 27081 20027 27115
rect 3801 27013 3835 27047
rect 3893 27013 3927 27047
rect 10517 27013 10551 27047
rect 12817 27013 12851 27047
rect 18061 27013 18095 27047
rect 23121 27013 23155 27047
rect 25145 27013 25179 27047
rect 3132 26945 3166 26979
rect 6561 26945 6595 26979
rect 9137 26945 9171 26979
rect 12541 26945 12575 26979
rect 15117 26945 15151 26979
rect 17969 26945 18003 26979
rect 19901 26945 19935 26979
rect 20729 26945 20763 26979
rect 22385 26945 22419 26979
rect 4445 26877 4479 26911
rect 6837 26877 6871 26911
rect 9229 26877 9263 26911
rect 9413 26877 9447 26911
rect 15301 26877 15335 26911
rect 18245 26877 18279 26911
rect 20177 26877 20211 26911
rect 22845 26877 22879 26911
rect 24593 26877 24627 26911
rect 8309 26809 8343 26843
rect 10701 26809 10735 26843
rect 25329 26809 25363 26843
rect 8769 26741 8803 26775
rect 14289 26741 14323 26775
rect 14749 26741 14783 26775
rect 17325 26741 17359 26775
rect 19533 26741 19567 26775
rect 22201 26741 22235 26775
rect 4077 26537 4111 26571
rect 8217 26537 8251 26571
rect 14381 26537 14415 26571
rect 17141 26537 17175 26571
rect 23857 26537 23891 26571
rect 25145 26537 25179 26571
rect 12173 26469 12207 26503
rect 19441 26469 19475 26503
rect 22385 26469 22419 26503
rect 22845 26469 22879 26503
rect 6469 26401 6503 26435
rect 6745 26401 6779 26435
rect 9137 26401 9171 26435
rect 10241 26401 10275 26435
rect 12725 26401 12759 26435
rect 15669 26401 15703 26435
rect 19901 26401 19935 26435
rect 20085 26401 20119 26435
rect 20637 26401 20671 26435
rect 23489 26401 23523 26435
rect 1777 26333 1811 26367
rect 9965 26333 9999 26367
rect 12541 26333 12575 26367
rect 12633 26333 12667 26367
rect 15393 26333 15427 26367
rect 19809 26333 19843 26367
rect 23213 26333 23247 26367
rect 24685 26333 24719 26367
rect 2789 26265 2823 26299
rect 8677 26265 8711 26299
rect 17509 26265 17543 26299
rect 20913 26265 20947 26299
rect 23305 26265 23339 26299
rect 24869 26265 24903 26299
rect 11713 26197 11747 26231
rect 17601 26197 17635 26231
rect 2145 25993 2179 26027
rect 9229 25993 9263 26027
rect 10793 25993 10827 26027
rect 10885 25993 10919 26027
rect 15853 25993 15887 26027
rect 19349 25993 19383 26027
rect 20269 25993 20303 26027
rect 20361 25993 20395 26027
rect 22477 25993 22511 26027
rect 8493 25925 8527 25959
rect 14749 25925 14783 25959
rect 20913 25925 20947 25959
rect 23305 25925 23339 25959
rect 2329 25857 2363 25891
rect 3065 25857 3099 25891
rect 4169 25857 4203 25891
rect 9597 25857 9631 25891
rect 12725 25857 12759 25891
rect 15761 25857 15795 25891
rect 17601 25857 17635 25891
rect 22385 25857 22419 25891
rect 23949 25857 23983 25891
rect 3249 25789 3283 25823
rect 8033 25789 8067 25823
rect 9689 25789 9723 25823
rect 9781 25789 9815 25823
rect 10977 25789 11011 25823
rect 11989 25789 12023 25823
rect 13001 25789 13035 25823
rect 14473 25789 14507 25823
rect 16037 25789 16071 25823
rect 17877 25789 17911 25823
rect 20545 25789 20579 25823
rect 21281 25789 21315 25823
rect 22569 25789 22603 25823
rect 25145 25789 25179 25823
rect 3433 25721 3467 25755
rect 4629 25721 4663 25755
rect 19901 25721 19935 25755
rect 23489 25721 23523 25755
rect 4261 25653 4295 25687
rect 8861 25653 8895 25687
rect 10425 25653 10459 25687
rect 15393 25653 15427 25687
rect 22017 25653 22051 25687
rect 11437 25449 11471 25483
rect 14749 25449 14783 25483
rect 17969 25449 18003 25483
rect 23121 25449 23155 25483
rect 23397 25449 23431 25483
rect 25145 25449 25179 25483
rect 25513 25449 25547 25483
rect 22109 25381 22143 25415
rect 6837 25313 6871 25347
rect 9413 25313 9447 25347
rect 10609 25313 10643 25347
rect 11989 25313 12023 25347
rect 13185 25313 13219 25347
rect 15301 25313 15335 25347
rect 15945 25313 15979 25347
rect 16221 25313 16255 25347
rect 19901 25313 19935 25347
rect 20085 25313 20119 25347
rect 22661 25313 22695 25347
rect 4052 25245 4086 25279
rect 10425 25245 10459 25279
rect 10517 25245 10551 25279
rect 11805 25245 11839 25279
rect 13093 25245 13127 25279
rect 19809 25245 19843 25279
rect 22477 25245 22511 25279
rect 23857 25245 23891 25279
rect 24685 25245 24719 25279
rect 7113 25177 7147 25211
rect 8953 25177 8987 25211
rect 22569 25177 22603 25211
rect 24869 25177 24903 25211
rect 4123 25109 4157 25143
rect 8585 25109 8619 25143
rect 10057 25109 10091 25143
rect 11161 25109 11195 25143
rect 11897 25109 11931 25143
rect 12633 25109 12667 25143
rect 13001 25109 13035 25143
rect 15117 25109 15151 25143
rect 15209 25109 15243 25143
rect 17693 25109 17727 25143
rect 18245 25109 18279 25143
rect 19441 25109 19475 25143
rect 23949 25109 23983 25143
rect 5457 24905 5491 24939
rect 8033 24905 8067 24939
rect 15209 24905 15243 24939
rect 16865 24905 16899 24939
rect 9229 24837 9263 24871
rect 12081 24837 12115 24871
rect 17233 24837 17267 24871
rect 18429 24837 18463 24871
rect 23213 24837 23247 24871
rect 7389 24769 7423 24803
rect 10057 24769 10091 24803
rect 12173 24769 12207 24803
rect 13185 24769 13219 24803
rect 13829 24769 13863 24803
rect 15301 24769 15335 24803
rect 17325 24769 17359 24803
rect 20637 24769 20671 24803
rect 25329 24769 25363 24803
rect 3709 24701 3743 24735
rect 3985 24701 4019 24735
rect 8125 24701 8159 24735
rect 8217 24701 8251 24735
rect 9321 24701 9355 24735
rect 9413 24701 9447 24735
rect 12265 24701 12299 24735
rect 13921 24701 13955 24735
rect 14105 24701 14139 24735
rect 15393 24701 15427 24735
rect 17509 24701 17543 24735
rect 18521 24701 18555 24735
rect 18613 24701 18647 24735
rect 20729 24701 20763 24735
rect 20821 24701 20855 24735
rect 22937 24701 22971 24735
rect 24685 24701 24719 24735
rect 7665 24633 7699 24667
rect 11713 24633 11747 24667
rect 13461 24633 13495 24667
rect 5825 24565 5859 24599
rect 8861 24565 8895 24599
rect 12725 24565 12759 24599
rect 13001 24565 13035 24599
rect 14565 24565 14599 24599
rect 14841 24565 14875 24599
rect 16497 24565 16531 24599
rect 18061 24565 18095 24599
rect 19901 24565 19935 24599
rect 20269 24565 20303 24599
rect 25145 24565 25179 24599
rect 3249 24361 3283 24395
rect 3433 24361 3467 24395
rect 5733 24361 5767 24395
rect 6193 24361 6227 24395
rect 8769 24361 8803 24395
rect 13737 24361 13771 24395
rect 18245 24293 18279 24327
rect 4261 24225 4295 24259
rect 10057 24225 10091 24259
rect 10517 24225 10551 24259
rect 11345 24225 11379 24259
rect 12541 24225 12575 24259
rect 13185 24225 13219 24259
rect 14289 24225 14323 24259
rect 16865 24225 16899 24259
rect 17049 24225 17083 24259
rect 19717 24225 19751 24259
rect 23857 24225 23891 24259
rect 25145 24225 25179 24259
rect 2237 24157 2271 24191
rect 2973 24157 3007 24191
rect 3985 24157 4019 24191
rect 6377 24157 6411 24191
rect 11161 24157 11195 24191
rect 11253 24157 11287 24191
rect 16773 24157 16807 24191
rect 17785 24157 17819 24191
rect 22017 24157 22051 24191
rect 22845 24157 22879 24191
rect 24961 24157 24995 24191
rect 25053 24157 25087 24191
rect 2697 24089 2731 24123
rect 9873 24089 9907 24123
rect 12449 24089 12483 24123
rect 19993 24089 20027 24123
rect 22201 24089 22235 24123
rect 2053 24021 2087 24055
rect 6745 24021 6779 24055
rect 9413 24021 9447 24055
rect 9781 24021 9815 24055
rect 10793 24021 10827 24055
rect 11989 24021 12023 24055
rect 12357 24021 12391 24055
rect 16405 24021 16439 24055
rect 17601 24021 17635 24055
rect 18153 24021 18187 24055
rect 21465 24021 21499 24055
rect 24593 24021 24627 24055
rect 6009 23817 6043 23851
rect 9413 23817 9447 23851
rect 9873 23817 9907 23851
rect 21649 23817 21683 23851
rect 25145 23817 25179 23851
rect 6469 23749 6503 23783
rect 10333 23749 10367 23783
rect 11805 23749 11839 23783
rect 1777 23681 1811 23715
rect 25329 23681 25363 23715
rect 2053 23613 2087 23647
rect 4261 23613 4295 23647
rect 4537 23613 4571 23647
rect 7665 23613 7699 23647
rect 7941 23613 7975 23647
rect 10885 23613 10919 23647
rect 12449 23613 12483 23647
rect 17049 23613 17083 23647
rect 18797 23613 18831 23647
rect 19073 23613 19107 23647
rect 20821 23613 20855 23647
rect 22937 23613 22971 23647
rect 23213 23613 23247 23647
rect 24685 23613 24719 23647
rect 11529 23477 11563 23511
rect 12173 23477 12207 23511
rect 12541 23477 12575 23511
rect 13921 23477 13955 23511
rect 21097 23477 21131 23511
rect 2053 23273 2087 23307
rect 3157 23273 3191 23307
rect 7573 23273 7607 23307
rect 16037 23273 16071 23307
rect 18521 23273 18555 23307
rect 21189 23273 21223 23307
rect 7849 23205 7883 23239
rect 11345 23205 11379 23239
rect 13001 23205 13035 23239
rect 2973 23137 3007 23171
rect 5825 23137 5859 23171
rect 11897 23137 11931 23171
rect 13553 23137 13587 23171
rect 14289 23137 14323 23171
rect 16497 23137 16531 23171
rect 19441 23137 19475 23171
rect 22017 23137 22051 23171
rect 23857 23137 23891 23171
rect 25053 23137 25087 23171
rect 25145 23137 25179 23171
rect 2237 23069 2271 23103
rect 2789 23069 2823 23103
rect 4112 23069 4146 23103
rect 4215 23069 4249 23103
rect 9965 23069 9999 23103
rect 11713 23069 11747 23103
rect 11805 23069 11839 23103
rect 13369 23069 13403 23103
rect 22845 23069 22879 23103
rect 24961 23069 24995 23103
rect 6101 23001 6135 23035
rect 10701 23001 10735 23035
rect 12541 23001 12575 23035
rect 13461 23001 13495 23035
rect 14565 23001 14599 23035
rect 16773 23001 16807 23035
rect 19717 23001 19751 23035
rect 12633 22933 12667 22967
rect 18245 22933 18279 22967
rect 21465 22933 21499 22967
rect 24593 22933 24627 22967
rect 2053 22729 2087 22763
rect 5641 22729 5675 22763
rect 6837 22729 6871 22763
rect 7205 22729 7239 22763
rect 10149 22729 10183 22763
rect 10885 22729 10919 22763
rect 12357 22729 12391 22763
rect 13093 22729 13127 22763
rect 15209 22729 15243 22763
rect 16221 22729 16255 22763
rect 17509 22729 17543 22763
rect 23765 22729 23799 22763
rect 24225 22729 24259 22763
rect 24317 22729 24351 22763
rect 24777 22729 24811 22763
rect 25421 22729 25455 22763
rect 12449 22661 12483 22695
rect 13277 22661 13311 22695
rect 16313 22661 16347 22695
rect 17877 22661 17911 22695
rect 18613 22661 18647 22695
rect 19717 22661 19751 22695
rect 20545 22661 20579 22695
rect 2237 22593 2271 22627
rect 5733 22593 5767 22627
rect 8033 22593 8067 22627
rect 9229 22593 9263 22627
rect 10793 22593 10827 22627
rect 15117 22593 15151 22627
rect 19625 22593 19659 22627
rect 21373 22593 21407 22627
rect 22017 22593 22051 22627
rect 5917 22525 5951 22559
rect 7297 22525 7331 22559
rect 7481 22525 7515 22559
rect 8861 22525 8895 22559
rect 10977 22525 11011 22559
rect 12633 22525 12667 22559
rect 13921 22525 13955 22559
rect 15393 22525 15427 22559
rect 19809 22525 19843 22559
rect 22293 22525 22327 22559
rect 10425 22457 10459 22491
rect 11989 22457 12023 22491
rect 5273 22389 5307 22423
rect 11621 22389 11655 22423
rect 14749 22389 14783 22423
rect 19257 22389 19291 22423
rect 16313 22185 16347 22219
rect 19698 22185 19732 22219
rect 21189 22185 21223 22219
rect 16865 22117 16899 22151
rect 18061 22117 18095 22151
rect 11989 22049 12023 22083
rect 14289 22049 14323 22083
rect 16037 22049 16071 22083
rect 17509 22049 17543 22083
rect 18521 22049 18555 22083
rect 18705 22049 18739 22083
rect 22017 22049 22051 22083
rect 22293 22049 22327 22083
rect 24041 22049 24075 22083
rect 11161 21981 11195 22015
rect 13277 21981 13311 22015
rect 17233 21981 17267 22015
rect 19441 21981 19475 22015
rect 24869 21981 24903 22015
rect 11805 21913 11839 21947
rect 12541 21913 12575 21947
rect 14565 21913 14599 21947
rect 18429 21913 18463 21947
rect 21465 21913 21499 21947
rect 24685 21913 24719 21947
rect 4445 21845 4479 21879
rect 10885 21845 10919 21879
rect 11437 21845 11471 21879
rect 11897 21845 11931 21879
rect 13093 21845 13127 21879
rect 16589 21845 16623 21879
rect 17325 21845 17359 21879
rect 7113 21641 7147 21675
rect 7481 21641 7515 21675
rect 8309 21641 8343 21675
rect 8677 21641 8711 21675
rect 9873 21641 9907 21675
rect 11713 21641 11747 21675
rect 12081 21641 12115 21675
rect 13553 21641 13587 21675
rect 13921 21641 13955 21675
rect 14013 21641 14047 21675
rect 22569 21641 22603 21675
rect 23673 21573 23707 21607
rect 1777 21505 1811 21539
rect 3433 21505 3467 21539
rect 4537 21505 4571 21539
rect 7573 21505 7607 21539
rect 12173 21505 12207 21539
rect 15209 21505 15243 21539
rect 16221 21505 16255 21539
rect 17049 21505 17083 21539
rect 18705 21505 18739 21539
rect 22477 21505 22511 21539
rect 23397 21505 23431 21539
rect 2053 21437 2087 21471
rect 3617 21437 3651 21471
rect 4997 21437 5031 21471
rect 7665 21437 7699 21471
rect 8769 21437 8803 21471
rect 8861 21437 8895 21471
rect 9965 21437 9999 21471
rect 10057 21437 10091 21471
rect 12265 21437 12299 21471
rect 14197 21437 14231 21471
rect 15301 21437 15335 21471
rect 15393 21437 15427 21471
rect 17693 21437 17727 21471
rect 22753 21437 22787 21471
rect 25145 21437 25179 21471
rect 3801 21369 3835 21403
rect 9505 21369 9539 21403
rect 16037 21369 16071 21403
rect 4813 21301 4847 21335
rect 14841 21301 14875 21335
rect 16865 21301 16899 21335
rect 18521 21301 18555 21335
rect 20453 21301 20487 21335
rect 22109 21301 22143 21335
rect 3157 21097 3191 21131
rect 7849 21097 7883 21131
rect 11897 21097 11931 21131
rect 13737 21097 13771 21131
rect 22017 21097 22051 21131
rect 4077 21029 4111 21063
rect 16313 21029 16347 21063
rect 17233 21029 17267 21063
rect 2789 20961 2823 20995
rect 8493 20961 8527 20995
rect 11529 20961 11563 20995
rect 13829 20961 13863 20995
rect 14933 20961 14967 20995
rect 17877 20961 17911 20995
rect 19901 20961 19935 20995
rect 23857 20961 23891 20995
rect 2237 20893 2271 20927
rect 2973 20893 3007 20927
rect 4261 20893 4295 20927
rect 9781 20893 9815 20927
rect 14841 20893 14875 20927
rect 15761 20893 15795 20927
rect 16129 20893 16163 20927
rect 17601 20893 17635 20927
rect 18889 20893 18923 20927
rect 22661 20893 22695 20927
rect 8309 20825 8343 20859
rect 10057 20825 10091 20859
rect 14749 20825 14783 20859
rect 20177 20825 20211 20859
rect 2053 20757 2087 20791
rect 7481 20757 7515 20791
rect 8217 20757 8251 20791
rect 14381 20757 14415 20791
rect 15577 20757 15611 20791
rect 16865 20757 16899 20791
rect 17693 20757 17727 20791
rect 18705 20757 18739 20791
rect 21649 20757 21683 20791
rect 22385 20757 22419 20791
rect 9965 20553 9999 20587
rect 12449 20553 12483 20587
rect 13277 20553 13311 20587
rect 17325 20553 17359 20587
rect 19349 20553 19383 20587
rect 19441 20553 19475 20587
rect 4261 20485 4295 20519
rect 6009 20485 6043 20519
rect 10425 20485 10459 20519
rect 17693 20485 17727 20519
rect 23305 20485 23339 20519
rect 3985 20417 4019 20451
rect 6561 20417 6595 20451
rect 9137 20417 9171 20451
rect 10333 20417 10367 20451
rect 15669 20417 15703 20451
rect 18521 20417 18555 20451
rect 22293 20417 22327 20451
rect 24133 20417 24167 20451
rect 6837 20349 6871 20383
rect 9229 20349 9263 20383
rect 9413 20349 9447 20383
rect 10517 20349 10551 20383
rect 12541 20349 12575 20383
rect 12725 20349 12759 20383
rect 19625 20349 19659 20383
rect 24685 20349 24719 20383
rect 8769 20281 8803 20315
rect 17877 20281 17911 20315
rect 5733 20213 5767 20247
rect 8309 20213 8343 20247
rect 12081 20213 12115 20247
rect 13737 20213 13771 20247
rect 14657 20213 14691 20247
rect 15485 20213 15519 20247
rect 18337 20213 18371 20247
rect 18981 20213 19015 20247
rect 5089 20009 5123 20043
rect 11713 20009 11747 20043
rect 14289 20009 14323 20043
rect 20361 20009 20395 20043
rect 15393 19941 15427 19975
rect 5733 19873 5767 19907
rect 6009 19873 6043 19907
rect 9137 19873 9171 19907
rect 11161 19873 11195 19907
rect 12265 19873 12299 19907
rect 14841 19873 14875 19907
rect 23857 19873 23891 19907
rect 5273 19805 5307 19839
rect 7757 19805 7791 19839
rect 8401 19805 8435 19839
rect 12081 19805 12115 19839
rect 13921 19805 13955 19839
rect 17233 19805 17267 19839
rect 17785 19805 17819 19839
rect 18705 19805 18739 19839
rect 22017 19805 22051 19839
rect 22845 19805 22879 19839
rect 9413 19737 9447 19771
rect 12173 19737 12207 19771
rect 14657 19737 14691 19771
rect 17325 19737 17359 19771
rect 17969 19737 18003 19771
rect 22201 19737 22235 19771
rect 7481 19669 7515 19703
rect 8677 19669 8711 19703
rect 14749 19669 14783 19703
rect 18521 19669 18555 19703
rect 19349 19669 19383 19703
rect 2053 19465 2087 19499
rect 4721 19465 4755 19499
rect 9229 19465 9263 19499
rect 11713 19465 11747 19499
rect 12081 19465 12115 19499
rect 16865 19465 16899 19499
rect 17509 19465 17543 19499
rect 19441 19465 19475 19499
rect 19809 19465 19843 19499
rect 19901 19465 19935 19499
rect 20729 19465 20763 19499
rect 21189 19465 21223 19499
rect 23765 19465 23799 19499
rect 18797 19397 18831 19431
rect 2237 19329 2271 19363
rect 3065 19329 3099 19363
rect 3893 19329 3927 19363
rect 4905 19329 4939 19363
rect 6561 19329 6595 19363
rect 9137 19329 9171 19363
rect 12173 19329 12207 19363
rect 13921 19329 13955 19363
rect 17049 19329 17083 19363
rect 17877 19329 17911 19363
rect 21097 19329 21131 19363
rect 6837 19261 6871 19295
rect 9321 19261 9355 19295
rect 11161 19261 11195 19295
rect 12265 19261 12299 19295
rect 13277 19261 13311 19295
rect 14013 19261 14047 19295
rect 14197 19261 14231 19295
rect 17969 19261 18003 19295
rect 18153 19261 18187 19295
rect 20085 19261 20119 19295
rect 21373 19261 21407 19295
rect 22017 19261 22051 19295
rect 22293 19261 22327 19295
rect 18981 19193 19015 19227
rect 8309 19125 8343 19159
rect 8769 19125 8803 19159
rect 10885 19125 10919 19159
rect 11253 19125 11287 19159
rect 13553 19125 13587 19159
rect 14657 19125 14691 19159
rect 14841 19125 14875 19159
rect 24041 19125 24075 19159
rect 8953 18921 8987 18955
rect 14289 18921 14323 18955
rect 17969 18921 18003 18955
rect 18981 18921 19015 18955
rect 24041 18921 24075 18955
rect 2053 18785 2087 18819
rect 5089 18785 5123 18819
rect 13553 18785 13587 18819
rect 14841 18785 14875 18819
rect 18337 18785 18371 18819
rect 1777 18717 1811 18751
rect 4077 18717 4111 18751
rect 9781 18717 9815 18751
rect 11897 18717 11931 18751
rect 13461 18717 13495 18751
rect 14657 18717 14691 18751
rect 16221 18717 16255 18751
rect 19625 18717 19659 18751
rect 20361 18717 20395 18751
rect 21557 18717 21591 18751
rect 22293 18717 22327 18751
rect 9229 18649 9263 18683
rect 10057 18649 10091 18683
rect 14749 18649 14783 18683
rect 16497 18649 16531 18683
rect 18521 18649 18555 18683
rect 21097 18649 21131 18683
rect 22569 18649 22603 18683
rect 8493 18581 8527 18615
rect 8677 18581 8711 18615
rect 9413 18581 9447 18615
rect 11529 18581 11563 18615
rect 12081 18581 12115 18615
rect 13001 18581 13035 18615
rect 13369 18581 13403 18615
rect 19717 18581 19751 18615
rect 21741 18581 21775 18615
rect 24409 18581 24443 18615
rect 7757 18377 7791 18411
rect 9689 18377 9723 18411
rect 11713 18377 11747 18411
rect 14289 18377 14323 18411
rect 14657 18377 14691 18411
rect 15393 18377 15427 18411
rect 21833 18377 21867 18411
rect 8493 18309 8527 18343
rect 12081 18309 12115 18343
rect 13829 18309 13863 18343
rect 19165 18309 19199 18343
rect 3341 18241 3375 18275
rect 7665 18241 7699 18275
rect 10793 18241 10827 18275
rect 14749 18241 14783 18275
rect 17509 18241 17543 18275
rect 21281 18241 21315 18275
rect 22385 18241 22419 18275
rect 3801 18173 3835 18207
rect 7849 18173 7883 18207
rect 9229 18173 9263 18207
rect 10885 18173 10919 18207
rect 10977 18173 11011 18207
rect 12173 18173 12207 18207
rect 12265 18173 12299 18207
rect 14933 18173 14967 18207
rect 18337 18173 18371 18207
rect 18889 18173 18923 18207
rect 23397 18173 23431 18207
rect 10425 18105 10459 18139
rect 13921 18105 13955 18139
rect 21465 18105 21499 18139
rect 6929 18037 6963 18071
rect 7297 18037 7331 18071
rect 10149 18037 10183 18071
rect 13553 18037 13587 18071
rect 17141 18037 17175 18071
rect 20637 18037 20671 18071
rect 23949 18037 23983 18071
rect 6285 17833 6319 17867
rect 9137 17833 9171 17867
rect 12541 17833 12575 17867
rect 21649 17833 21683 17867
rect 23857 17833 23891 17867
rect 17233 17765 17267 17799
rect 6837 17697 6871 17731
rect 8125 17697 8159 17731
rect 9689 17697 9723 17731
rect 12725 17697 12759 17731
rect 13553 17697 13587 17731
rect 14841 17697 14875 17731
rect 16681 17697 16715 17731
rect 16865 17697 16899 17731
rect 19901 17697 19935 17731
rect 22109 17697 22143 17731
rect 22385 17697 22419 17731
rect 7941 17629 7975 17663
rect 11897 17629 11931 17663
rect 13461 17629 13495 17663
rect 14657 17629 14691 17663
rect 15577 17629 15611 17663
rect 24869 17629 24903 17663
rect 6653 17561 6687 17595
rect 10517 17561 10551 17595
rect 11345 17561 11379 17595
rect 13369 17561 13403 17595
rect 20177 17561 20211 17595
rect 24133 17561 24167 17595
rect 6745 17493 6779 17527
rect 7481 17493 7515 17527
rect 7849 17493 7883 17527
rect 8769 17493 8803 17527
rect 9505 17493 9539 17527
rect 9597 17493 9631 17527
rect 13001 17493 13035 17527
rect 14289 17493 14323 17527
rect 14749 17493 14783 17527
rect 15669 17493 15703 17527
rect 16221 17493 16255 17527
rect 16589 17493 16623 17527
rect 24685 17493 24719 17527
rect 10057 17289 10091 17323
rect 11529 17289 11563 17323
rect 3985 17221 4019 17255
rect 10425 17221 10459 17255
rect 15117 17221 15151 17255
rect 19809 17221 19843 17255
rect 23305 17221 23339 17255
rect 3157 17153 3191 17187
rect 9045 17153 9079 17187
rect 17049 17153 17083 17187
rect 17693 17153 17727 17187
rect 21281 17153 21315 17187
rect 22109 17153 22143 17187
rect 23949 17153 23983 17187
rect 6561 17085 6595 17119
rect 6837 17085 6871 17119
rect 8585 17085 8619 17119
rect 10517 17085 10551 17119
rect 10701 17085 10735 17119
rect 12633 17085 12667 17119
rect 12909 17085 12943 17119
rect 14933 17085 14967 17119
rect 17969 17085 18003 17119
rect 19441 17085 19475 17119
rect 20453 17085 20487 17119
rect 24409 17085 24443 17119
rect 14381 17017 14415 17051
rect 16037 17017 16071 17051
rect 21465 17017 21499 17051
rect 9137 16949 9171 16983
rect 9505 16949 9539 16983
rect 14749 16949 14783 16983
rect 16865 16949 16899 16983
rect 5628 16745 5662 16779
rect 7113 16745 7147 16779
rect 7481 16745 7515 16779
rect 9137 16745 9171 16779
rect 10517 16745 10551 16779
rect 19349 16745 19383 16779
rect 8677 16677 8711 16711
rect 10241 16677 10275 16711
rect 5365 16609 5399 16643
rect 7665 16609 7699 16643
rect 9689 16609 9723 16643
rect 11069 16609 11103 16643
rect 12265 16609 12299 16643
rect 12357 16609 12391 16643
rect 14933 16609 14967 16643
rect 15761 16609 15795 16643
rect 15945 16609 15979 16643
rect 20637 16609 20671 16643
rect 21741 16609 21775 16643
rect 22017 16609 22051 16643
rect 23765 16609 23799 16643
rect 1593 16541 1627 16575
rect 9505 16541 9539 16575
rect 10885 16541 10919 16575
rect 12173 16541 12207 16575
rect 20453 16541 20487 16575
rect 20545 16541 20579 16575
rect 2513 16473 2547 16507
rect 8493 16405 8527 16439
rect 9597 16405 9631 16439
rect 10977 16405 11011 16439
rect 11805 16405 11839 16439
rect 15301 16405 15335 16439
rect 15669 16405 15703 16439
rect 16405 16405 16439 16439
rect 20085 16405 20119 16439
rect 23489 16405 23523 16439
rect 8953 16201 8987 16235
rect 10149 16201 10183 16235
rect 10609 16201 10643 16235
rect 11713 16201 11747 16235
rect 12081 16201 12115 16235
rect 13737 16201 13771 16235
rect 14749 16201 14783 16235
rect 18613 16201 18647 16235
rect 18889 16201 18923 16235
rect 19257 16201 19291 16235
rect 2513 16133 2547 16167
rect 9321 16133 9355 16167
rect 13093 16133 13127 16167
rect 14197 16133 14231 16167
rect 15945 16133 15979 16167
rect 16405 16133 16439 16167
rect 17141 16133 17175 16167
rect 22477 16133 22511 16167
rect 6653 16065 6687 16099
rect 10517 16065 10551 16099
rect 12173 16065 12207 16099
rect 16865 16065 16899 16099
rect 19625 16065 19659 16099
rect 20453 16065 20487 16099
rect 21281 16065 21315 16099
rect 22385 16065 22419 16099
rect 23489 16065 23523 16099
rect 24133 16065 24167 16099
rect 6929 15997 6963 16031
rect 8401 15997 8435 16031
rect 9413 15997 9447 16031
rect 9505 15997 9539 16031
rect 10701 15997 10735 16031
rect 12265 15997 12299 16031
rect 19717 15997 19751 16031
rect 19901 15997 19935 16031
rect 22569 15997 22603 16031
rect 24409 15997 24443 16031
rect 21465 15929 21499 15963
rect 2605 15861 2639 15895
rect 14289 15861 14323 15895
rect 16037 15861 16071 15895
rect 22017 15861 22051 15895
rect 23305 15861 23339 15895
rect 8769 15657 8803 15691
rect 9965 15657 9999 15691
rect 14289 15657 14323 15691
rect 21097 15657 21131 15691
rect 17325 15589 17359 15623
rect 11069 15521 11103 15555
rect 14841 15521 14875 15555
rect 17877 15521 17911 15555
rect 20085 15521 20119 15555
rect 13461 15453 13495 15487
rect 14657 15453 14691 15487
rect 19901 15453 19935 15487
rect 20821 15453 20855 15487
rect 21833 15453 21867 15487
rect 22845 15453 22879 15487
rect 11345 15385 11379 15419
rect 13645 15385 13679 15419
rect 17785 15385 17819 15419
rect 18337 15385 18371 15419
rect 23857 15385 23891 15419
rect 8493 15317 8527 15351
rect 10241 15317 10275 15351
rect 10793 15317 10827 15351
rect 12817 15317 12851 15351
rect 14749 15317 14783 15351
rect 17049 15317 17083 15351
rect 17693 15317 17727 15351
rect 18705 15317 18739 15351
rect 19441 15317 19475 15351
rect 19809 15317 19843 15351
rect 20637 15317 20671 15351
rect 21925 15317 21959 15351
rect 13001 15113 13035 15147
rect 14197 15113 14231 15147
rect 18797 15113 18831 15147
rect 18889 15113 18923 15147
rect 22293 15113 22327 15147
rect 9413 15045 9447 15079
rect 11621 15045 11655 15079
rect 13369 15045 13403 15079
rect 15669 15045 15703 15079
rect 16129 15045 16163 15079
rect 20085 15045 20119 15079
rect 14565 14977 14599 15011
rect 14657 14977 14691 15011
rect 15301 14977 15335 15011
rect 17233 14977 17267 15011
rect 17693 14977 17727 15011
rect 19809 14977 19843 15011
rect 23397 14977 23431 15011
rect 24133 14977 24167 15011
rect 9137 14909 9171 14943
rect 11161 14909 11195 14943
rect 13461 14909 13495 14943
rect 13553 14909 13587 14943
rect 14841 14909 14875 14943
rect 18981 14909 19015 14943
rect 24777 14909 24811 14943
rect 12725 14841 12759 14875
rect 17417 14841 17451 14875
rect 15761 14773 15795 14807
rect 18429 14773 18463 14807
rect 19625 14773 19659 14807
rect 23213 14773 23247 14807
rect 13001 14569 13035 14603
rect 14381 14569 14415 14603
rect 14473 14569 14507 14603
rect 17141 14569 17175 14603
rect 18705 14569 18739 14603
rect 12081 14501 12115 14535
rect 14105 14501 14139 14535
rect 9965 14433 9999 14467
rect 12725 14433 12759 14467
rect 13553 14433 13587 14467
rect 15393 14433 15427 14467
rect 21189 14433 21223 14467
rect 13369 14365 13403 14399
rect 18245 14365 18279 14399
rect 18613 14365 18647 14399
rect 20913 14365 20947 14399
rect 22937 14365 22971 14399
rect 10241 14297 10275 14331
rect 12541 14297 12575 14331
rect 13461 14297 13495 14331
rect 15669 14297 15703 14331
rect 11713 14229 11747 14263
rect 17417 14229 17451 14263
rect 19441 14229 19475 14263
rect 19993 14229 20027 14263
rect 22661 14229 22695 14263
rect 11897 14025 11931 14059
rect 12725 14025 12759 14059
rect 18889 14025 18923 14059
rect 19809 14025 19843 14059
rect 23029 14025 23063 14059
rect 10057 13957 10091 13991
rect 13553 13957 13587 13991
rect 14013 13957 14047 13991
rect 17417 13957 17451 13991
rect 19717 13957 19751 13991
rect 21189 13957 21223 13991
rect 21833 13957 21867 13991
rect 1777 13889 1811 13923
rect 8033 13889 8067 13923
rect 12633 13889 12667 13923
rect 17141 13889 17175 13923
rect 20453 13889 20487 13923
rect 23213 13889 23247 13923
rect 23949 13889 23983 13923
rect 2053 13821 2087 13855
rect 9781 13821 9815 13855
rect 12817 13821 12851 13855
rect 13737 13821 13771 13855
rect 20637 13821 20671 13855
rect 21373 13821 21407 13855
rect 24685 13821 24719 13855
rect 8296 13685 8330 13719
rect 12265 13685 12299 13719
rect 19165 13685 19199 13719
rect 11621 13481 11655 13515
rect 11989 13481 12023 13515
rect 12357 13481 12391 13515
rect 13369 13481 13403 13515
rect 16313 13481 16347 13515
rect 20729 13481 20763 13515
rect 9045 13413 9079 13447
rect 17785 13413 17819 13447
rect 9137 13345 9171 13379
rect 9873 13345 9907 13379
rect 10149 13345 10183 13379
rect 12909 13345 12943 13379
rect 14565 13345 14599 13379
rect 18245 13345 18279 13379
rect 18429 13345 18463 13379
rect 19993 13345 20027 13379
rect 6837 13277 6871 13311
rect 12725 13277 12759 13311
rect 18797 13277 18831 13311
rect 19809 13277 19843 13311
rect 22661 13277 22695 13311
rect 7113 13209 7147 13243
rect 12817 13209 12851 13243
rect 14841 13209 14875 13243
rect 19901 13209 19935 13243
rect 23857 13209 23891 13243
rect 8585 13141 8619 13175
rect 16865 13141 16899 13175
rect 17509 13141 17543 13175
rect 18153 13141 18187 13175
rect 19441 13141 19475 13175
rect 21557 13141 21591 13175
rect 22017 13141 22051 13175
rect 8677 12937 8711 12971
rect 11161 12937 11195 12971
rect 16129 12937 16163 12971
rect 17233 12937 17267 12971
rect 17325 12937 17359 12971
rect 18981 12937 19015 12971
rect 11529 12869 11563 12903
rect 13277 12869 13311 12903
rect 13737 12869 13771 12903
rect 14473 12869 14507 12903
rect 14933 12869 14967 12903
rect 15393 12869 15427 12903
rect 15853 12869 15887 12903
rect 16405 12869 16439 12903
rect 18521 12869 18555 12903
rect 8585 12801 8619 12835
rect 9413 12801 9447 12835
rect 22293 12801 22327 12835
rect 23305 12801 23339 12835
rect 23949 12801 23983 12835
rect 8769 12733 8803 12767
rect 9689 12733 9723 12767
rect 17417 12733 17451 12767
rect 19717 12733 19751 12767
rect 19993 12733 20027 12767
rect 21465 12733 21499 12767
rect 24777 12733 24811 12767
rect 13921 12665 13955 12699
rect 14657 12665 14691 12699
rect 16865 12665 16899 12699
rect 8217 12597 8251 12631
rect 15485 12597 15519 12631
rect 18613 12597 18647 12631
rect 13829 12393 13863 12427
rect 14105 12393 14139 12427
rect 14473 12393 14507 12427
rect 15669 12393 15703 12427
rect 18889 12393 18923 12427
rect 22661 12325 22695 12359
rect 11529 12257 11563 12291
rect 11805 12257 11839 12291
rect 15025 12257 15059 12291
rect 16129 12257 16163 12291
rect 16221 12257 16255 12291
rect 17141 12257 17175 12291
rect 17417 12257 17451 12291
rect 21557 12257 21591 12291
rect 21741 12257 21775 12291
rect 14841 12189 14875 12223
rect 20637 12189 20671 12223
rect 21465 12189 21499 12223
rect 22845 12189 22879 12223
rect 23489 12189 23523 12223
rect 16037 12121 16071 12155
rect 13277 12053 13311 12087
rect 13737 12053 13771 12087
rect 14933 12053 14967 12087
rect 19349 12053 19383 12087
rect 20453 12053 20487 12087
rect 21097 12053 21131 12087
rect 23305 12053 23339 12087
rect 15485 11849 15519 11883
rect 16037 11849 16071 11883
rect 19993 11849 20027 11883
rect 20361 11849 20395 11883
rect 13093 11781 13127 11815
rect 16957 11781 16991 11815
rect 17417 11781 17451 11815
rect 18521 11781 18555 11815
rect 20913 11781 20947 11815
rect 21373 11781 21407 11815
rect 12817 11713 12851 11747
rect 15393 11713 15427 11747
rect 18245 11713 18279 11747
rect 23305 11713 23339 11747
rect 15577 11645 15611 11679
rect 24041 11645 24075 11679
rect 14565 11577 14599 11611
rect 15025 11577 15059 11611
rect 21097 11577 21131 11611
rect 17049 11509 17083 11543
rect 15485 11305 15519 11339
rect 14749 11169 14783 11203
rect 16037 11169 16071 11203
rect 15853 11101 15887 11135
rect 15945 11033 15979 11067
rect 20821 11033 20855 11067
rect 21005 11033 21039 11067
rect 19625 10965 19659 10999
rect 15301 10761 15335 10795
rect 19533 10761 19567 10795
rect 20361 10761 20395 10795
rect 12081 10693 12115 10727
rect 12541 10693 12575 10727
rect 14841 10625 14875 10659
rect 18429 10625 18463 10659
rect 19625 10625 19659 10659
rect 20545 10625 20579 10659
rect 23397 10625 23431 10659
rect 23949 10625 23983 10659
rect 19809 10557 19843 10591
rect 24777 10557 24811 10591
rect 12265 10489 12299 10523
rect 14657 10489 14691 10523
rect 15209 10421 15243 10455
rect 18245 10421 18279 10455
rect 19165 10421 19199 10455
rect 23213 10421 23247 10455
rect 14657 10013 14691 10047
rect 16773 10013 16807 10047
rect 21465 10013 21499 10047
rect 22201 10013 22235 10047
rect 22661 10013 22695 10047
rect 23857 10013 23891 10047
rect 14841 9945 14875 9979
rect 24685 9945 24719 9979
rect 16865 9877 16899 9911
rect 21281 9877 21315 9911
rect 22017 9877 22051 9911
rect 24777 9877 24811 9911
rect 16957 9605 16991 9639
rect 5825 9537 5859 9571
rect 6929 9537 6963 9571
rect 19257 9537 19291 9571
rect 22937 9537 22971 9571
rect 23949 9537 23983 9571
rect 7021 9469 7055 9503
rect 7113 9469 7147 9503
rect 24409 9469 24443 9503
rect 6561 9401 6595 9435
rect 17141 9401 17175 9435
rect 19073 9333 19107 9367
rect 22753 9333 22787 9367
rect 24685 9061 24719 9095
rect 21741 8925 21775 8959
rect 23949 8925 23983 8959
rect 24869 8925 24903 8959
rect 21557 8789 21591 8823
rect 23765 8789 23799 8823
rect 19165 8517 19199 8551
rect 19625 8517 19659 8551
rect 20729 8517 20763 8551
rect 22293 8449 22327 8483
rect 23949 8449 23983 8483
rect 23305 8381 23339 8415
rect 24685 8381 24719 8415
rect 19349 8313 19383 8347
rect 20913 8313 20947 8347
rect 6469 8041 6503 8075
rect 6653 8041 6687 8075
rect 24593 8041 24627 8075
rect 4077 7905 4111 7939
rect 20453 7837 20487 7871
rect 21281 7837 21315 7871
rect 22845 7837 22879 7871
rect 24777 7837 24811 7871
rect 4353 7769 4387 7803
rect 6101 7769 6135 7803
rect 23857 7769 23891 7803
rect 20269 7701 20303 7735
rect 21097 7701 21131 7735
rect 18797 7429 18831 7463
rect 25145 7429 25179 7463
rect 20269 7361 20303 7395
rect 22109 7361 22143 7395
rect 23949 7361 23983 7395
rect 21281 7293 21315 7327
rect 22569 7293 22603 7327
rect 18981 7225 19015 7259
rect 19717 6749 19751 6783
rect 19993 6749 20027 6783
rect 20821 6749 20855 6783
rect 22845 6749 22879 6783
rect 24869 6749 24903 6783
rect 21833 6681 21867 6715
rect 23857 6681 23891 6715
rect 19533 6613 19567 6647
rect 24685 6613 24719 6647
rect 1869 6409 1903 6443
rect 3709 6409 3743 6443
rect 17969 6409 18003 6443
rect 1685 6273 1719 6307
rect 2605 6273 2639 6307
rect 3065 6273 3099 6307
rect 18245 6273 18279 6307
rect 20269 6273 20303 6307
rect 22017 6273 22051 6307
rect 23949 6273 23983 6307
rect 19441 6205 19475 6239
rect 21281 6205 21315 6239
rect 22477 6205 22511 6239
rect 24777 6205 24811 6239
rect 2421 6069 2455 6103
rect 3157 5865 3191 5899
rect 24777 5865 24811 5899
rect 2053 5797 2087 5831
rect 21005 5729 21039 5763
rect 22845 5729 22879 5763
rect 2513 5661 2547 5695
rect 17693 5661 17727 5695
rect 20545 5661 20579 5695
rect 22385 5661 22419 5695
rect 1869 5593 1903 5627
rect 3801 5593 3835 5627
rect 18705 5593 18739 5627
rect 24685 5593 24719 5627
rect 3617 5525 3651 5559
rect 3985 5525 4019 5559
rect 3065 5321 3099 5355
rect 3801 5321 3835 5355
rect 4353 5321 4387 5355
rect 5181 5321 5215 5355
rect 2421 5253 2455 5287
rect 20361 5253 20395 5287
rect 1777 5185 1811 5219
rect 2881 5185 2915 5219
rect 3617 5185 3651 5219
rect 4537 5185 4571 5219
rect 4997 5185 5031 5219
rect 17785 5185 17819 5219
rect 19533 5185 19567 5219
rect 22201 5185 22235 5219
rect 24041 5185 24075 5219
rect 18797 5117 18831 5151
rect 22477 5117 22511 5151
rect 24593 5117 24627 5151
rect 1501 4981 1535 5015
rect 6101 4981 6135 5015
rect 7389 4981 7423 5015
rect 4169 4777 4203 4811
rect 5917 4777 5951 4811
rect 6745 4777 6779 4811
rect 7757 4777 7791 4811
rect 8493 4777 8527 4811
rect 9781 4777 9815 4811
rect 23857 4777 23891 4811
rect 5181 4709 5215 4743
rect 11713 4709 11747 4743
rect 24869 4709 24903 4743
rect 3341 4641 3375 4675
rect 4537 4641 4571 4675
rect 19901 4641 19935 4675
rect 21741 4641 21775 4675
rect 1593 4573 1627 4607
rect 2697 4573 2731 4607
rect 3985 4573 4019 4607
rect 4997 4573 5031 4607
rect 5733 4573 5767 4607
rect 6561 4573 6595 4607
rect 8309 4573 8343 4607
rect 9597 4573 9631 4607
rect 11897 4573 11931 4607
rect 12173 4573 12207 4607
rect 17693 4573 17727 4607
rect 19441 4573 19475 4607
rect 21281 4573 21315 4607
rect 24041 4573 24075 4607
rect 7665 4505 7699 4539
rect 8953 4505 8987 4539
rect 10149 4505 10183 4539
rect 18705 4505 18739 4539
rect 24685 4505 24719 4539
rect 2237 4437 2271 4471
rect 7113 4437 7147 4471
rect 9137 4437 9171 4471
rect 10333 4437 10367 4471
rect 1777 4097 1811 4131
rect 2421 4097 2455 4131
rect 2973 4097 3007 4131
rect 3709 4097 3743 4131
rect 4629 4097 4663 4131
rect 5365 4097 5399 4131
rect 6009 4097 6043 4131
rect 6561 4097 6595 4131
rect 7205 4097 7239 4131
rect 7941 4097 7975 4131
rect 8677 4097 8711 4131
rect 9413 4097 9447 4131
rect 10333 4097 10367 4131
rect 11713 4097 11747 4131
rect 13645 4097 13679 4131
rect 16129 4097 16163 4131
rect 16865 4097 16899 4131
rect 18705 4097 18739 4131
rect 22201 4097 22235 4131
rect 24133 4097 24167 4131
rect 4353 4029 4387 4063
rect 10057 4029 10091 4063
rect 14013 4029 14047 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 22477 4029 22511 4063
rect 24777 4029 24811 4063
rect 8125 3961 8159 3995
rect 8861 3961 8895 3995
rect 11069 3961 11103 3995
rect 1501 3893 1535 3927
rect 3157 3893 3191 3927
rect 4905 3893 4939 3927
rect 5089 3893 5123 3927
rect 7573 3893 7607 3927
rect 10517 3893 10551 3927
rect 10885 3893 10919 3927
rect 11253 3893 11287 3927
rect 12357 3893 12391 3927
rect 16221 3893 16255 3927
rect 2329 3689 2363 3723
rect 3433 3689 3467 3723
rect 5273 3689 5307 3723
rect 6377 3689 6411 3723
rect 8585 3689 8619 3723
rect 9321 3689 9355 3723
rect 18613 3689 18647 3723
rect 3985 3621 4019 3655
rect 10977 3553 11011 3587
rect 11253 3553 11287 3587
rect 12817 3553 12851 3587
rect 15485 3553 15519 3587
rect 17325 3553 17359 3587
rect 19901 3553 19935 3587
rect 21741 3553 21775 3587
rect 1685 3485 1719 3519
rect 2789 3485 2823 3519
rect 4169 3485 4203 3519
rect 4629 3485 4663 3519
rect 5733 3485 5767 3519
rect 6837 3485 6871 3519
rect 7941 3485 7975 3519
rect 9137 3485 9171 3519
rect 9873 3485 9907 3519
rect 12541 3485 12575 3519
rect 15117 3485 15151 3519
rect 16865 3485 16899 3519
rect 19441 3485 19475 3519
rect 21465 3485 21499 3519
rect 23397 3485 23431 3519
rect 24041 3485 24075 3519
rect 24593 3485 24627 3519
rect 10517 3417 10551 3451
rect 7481 3349 7515 3383
rect 25237 3349 25271 3383
rect 2789 3145 2823 3179
rect 6009 3145 6043 3179
rect 8585 3145 8619 3179
rect 11897 3145 11931 3179
rect 23121 3145 23155 3179
rect 25145 3145 25179 3179
rect 2145 3009 2179 3043
rect 4629 3009 4663 3043
rect 5365 3009 5399 3043
rect 6561 3009 6595 3043
rect 6837 3009 6871 3043
rect 7941 3009 7975 3043
rect 9045 3009 9079 3043
rect 9321 3009 9355 3043
rect 10333 3009 10367 3043
rect 10609 3009 10643 3043
rect 11713 3009 11747 3043
rect 12633 3009 12667 3043
rect 14289 3009 14323 3043
rect 17049 3009 17083 3043
rect 18797 3009 18831 3043
rect 22477 3009 22511 3043
rect 25329 3009 25363 3043
rect 1869 2941 1903 2975
rect 3249 2941 3283 2975
rect 3525 2941 3559 2975
rect 13369 2941 13403 2975
rect 14749 2941 14783 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 1501 2873 1535 2907
rect 4813 2873 4847 2907
rect 1685 2805 1719 2839
rect 7481 2805 7515 2839
rect 23489 2805 23523 2839
rect 2329 2601 2363 2635
rect 3433 2601 3467 2635
rect 9873 2601 9907 2635
rect 11713 2601 11747 2635
rect 18613 2601 18647 2635
rect 25237 2601 25271 2635
rect 7205 2533 7239 2567
rect 14289 2533 14323 2567
rect 4997 2465 5031 2499
rect 6009 2465 6043 2499
rect 10333 2465 10367 2499
rect 14105 2465 14139 2499
rect 15209 2465 15243 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 22477 2465 22511 2499
rect 24041 2465 24075 2499
rect 1685 2397 1719 2431
rect 2789 2397 2823 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 6561 2397 6595 2431
rect 7665 2397 7699 2431
rect 7941 2397 7975 2431
rect 9229 2397 9263 2431
rect 10609 2397 10643 2431
rect 11897 2397 11931 2431
rect 12449 2397 12483 2431
rect 14657 2397 14691 2431
rect 16865 2397 16899 2431
rect 19533 2397 19567 2431
rect 22017 2397 22051 2431
rect 24593 2397 24627 2431
rect 13553 2329 13587 2363
rect 4169 2261 4203 2295
rect 6101 2261 6135 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 3970 54272 3976 54324
rect 4028 54272 4034 54324
rect 9950 54272 9956 54324
rect 10008 54272 10014 54324
rect 13998 54272 14004 54324
rect 14056 54312 14062 54324
rect 14093 54315 14151 54321
rect 14093 54312 14105 54315
rect 14056 54284 14105 54312
rect 14056 54272 14062 54284
rect 14093 54281 14105 54284
rect 14139 54281 14151 54315
rect 14093 54275 14151 54281
rect 14553 54315 14611 54321
rect 14553 54281 14565 54315
rect 14599 54312 14611 54315
rect 14734 54312 14740 54324
rect 14599 54284 14740 54312
rect 14599 54281 14611 54284
rect 14553 54275 14611 54281
rect 14734 54272 14740 54284
rect 14792 54272 14798 54324
rect 5813 54247 5871 54253
rect 5813 54213 5825 54247
rect 5859 54244 5871 54247
rect 7834 54244 7840 54256
rect 5859 54216 7840 54244
rect 5859 54213 5871 54216
rect 5813 54207 5871 54213
rect 7834 54204 7840 54216
rect 7892 54204 7898 54256
rect 8389 54247 8447 54253
rect 8389 54213 8401 54247
rect 8435 54244 8447 54247
rect 9968 54244 9996 54272
rect 8435 54216 9996 54244
rect 10965 54247 11023 54253
rect 8435 54213 8447 54216
rect 8389 54207 8447 54213
rect 10965 54213 10977 54247
rect 11011 54244 11023 54247
rect 11422 54244 11428 54256
rect 11011 54216 11428 54244
rect 11011 54213 11023 54216
rect 10965 54207 11023 54213
rect 11422 54204 11428 54216
rect 11480 54204 11486 54256
rect 12894 54244 12900 54256
rect 11900 54216 12900 54244
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 2314 54176 2320 54188
rect 2271 54148 2320 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 2314 54136 2320 54148
rect 2372 54136 2378 54188
rect 4614 54136 4620 54188
rect 4672 54136 4678 54188
rect 7377 54179 7435 54185
rect 7377 54145 7389 54179
rect 7423 54145 7435 54179
rect 7377 54139 7435 54145
rect 3237 54111 3295 54117
rect 3237 54077 3249 54111
rect 3283 54108 3295 54111
rect 5902 54108 5908 54120
rect 3283 54080 5908 54108
rect 3283 54077 3295 54080
rect 3237 54071 3295 54077
rect 5902 54068 5908 54080
rect 5960 54068 5966 54120
rect 7392 54108 7420 54139
rect 9950 54136 9956 54188
rect 10008 54136 10014 54188
rect 11606 54136 11612 54188
rect 11664 54176 11670 54188
rect 11900 54185 11928 54216
rect 12894 54204 12900 54216
rect 12952 54204 12958 54256
rect 13630 54204 13636 54256
rect 13688 54244 13694 54256
rect 14277 54247 14335 54253
rect 14277 54244 14289 54247
rect 13688 54216 14289 54244
rect 13688 54204 13694 54216
rect 14277 54213 14289 54216
rect 14323 54213 14335 54247
rect 14277 54207 14335 54213
rect 11885 54179 11943 54185
rect 11885 54176 11897 54179
rect 11664 54148 11897 54176
rect 11664 54136 11670 54148
rect 11885 54145 11897 54148
rect 11931 54145 11943 54179
rect 11885 54139 11943 54145
rect 12342 54136 12348 54188
rect 12400 54136 12406 54188
rect 14752 54176 14780 54272
rect 15562 54204 15568 54256
rect 15620 54244 15626 54256
rect 24121 54247 24179 54253
rect 24121 54244 24133 54247
rect 15620 54216 16574 54244
rect 15620 54204 15626 54216
rect 14829 54179 14887 54185
rect 14829 54176 14841 54179
rect 14752 54148 14841 54176
rect 14829 54145 14841 54148
rect 14875 54145 14887 54179
rect 14829 54139 14887 54145
rect 15473 54179 15531 54185
rect 15473 54145 15485 54179
rect 15519 54176 15531 54179
rect 15933 54179 15991 54185
rect 15933 54176 15945 54179
rect 15519 54148 15945 54176
rect 15519 54145 15531 54148
rect 15473 54139 15531 54145
rect 15933 54145 15945 54148
rect 15979 54145 15991 54179
rect 16546 54176 16574 54216
rect 22020 54216 24133 54244
rect 16853 54179 16911 54185
rect 16853 54176 16865 54179
rect 16546 54148 16865 54176
rect 15933 54139 15991 54145
rect 16853 54145 16865 54148
rect 16899 54176 16911 54179
rect 17402 54176 17408 54188
rect 16899 54148 17408 54176
rect 16899 54145 16911 54148
rect 16853 54139 16911 54145
rect 17402 54136 17408 54148
rect 17460 54136 17466 54188
rect 17954 54136 17960 54188
rect 18012 54176 18018 54188
rect 18877 54179 18935 54185
rect 18877 54176 18889 54179
rect 18012 54148 18889 54176
rect 18012 54136 18018 54148
rect 18877 54145 18889 54148
rect 18923 54145 18935 54179
rect 18877 54139 18935 54145
rect 19426 54136 19432 54188
rect 19484 54136 19490 54188
rect 20533 54179 20591 54185
rect 20533 54145 20545 54179
rect 20579 54145 20591 54179
rect 20533 54139 20591 54145
rect 11238 54108 11244 54120
rect 7392 54080 11244 54108
rect 11238 54068 11244 54080
rect 11296 54068 11302 54120
rect 12526 54068 12532 54120
rect 12584 54108 12590 54120
rect 12805 54111 12863 54117
rect 12805 54108 12817 54111
rect 12584 54080 12817 54108
rect 12584 54068 12590 54080
rect 12805 54077 12817 54080
rect 12851 54077 12863 54111
rect 12805 54071 12863 54077
rect 18690 54068 18696 54120
rect 18748 54108 18754 54120
rect 19150 54108 19156 54120
rect 18748 54080 19156 54108
rect 18748 54068 18754 54080
rect 19150 54068 19156 54080
rect 19208 54108 19214 54120
rect 20548 54108 20576 54139
rect 20714 54136 20720 54188
rect 20772 54176 20778 54188
rect 22020 54185 22048 54216
rect 24121 54213 24133 54216
rect 24167 54213 24179 54247
rect 24121 54207 24179 54213
rect 22005 54179 22063 54185
rect 22005 54176 22017 54179
rect 20772 54148 22017 54176
rect 20772 54136 20778 54148
rect 22005 54145 22017 54148
rect 22051 54145 22063 54179
rect 22005 54139 22063 54145
rect 23109 54179 23167 54185
rect 23109 54145 23121 54179
rect 23155 54145 23167 54179
rect 23109 54139 23167 54145
rect 19208 54080 20576 54108
rect 19208 54068 19214 54080
rect 21358 54068 21364 54120
rect 21416 54108 21422 54120
rect 23124 54108 23152 54139
rect 24026 54136 24032 54188
rect 24084 54176 24090 54188
rect 24581 54179 24639 54185
rect 24581 54176 24593 54179
rect 24084 54148 24593 54176
rect 24084 54136 24090 54148
rect 24581 54145 24593 54148
rect 24627 54176 24639 54179
rect 24670 54176 24676 54188
rect 24627 54148 24676 54176
rect 24627 54145 24639 54148
rect 24581 54139 24639 54145
rect 24670 54136 24676 54148
rect 24728 54136 24734 54188
rect 25133 54111 25191 54117
rect 25133 54108 25145 54111
rect 21416 54080 25145 54108
rect 21416 54068 21422 54080
rect 25133 54077 25145 54080
rect 25179 54077 25191 54111
rect 25133 54071 25191 54077
rect 20530 54000 20536 54052
rect 20588 54040 20594 54052
rect 21453 54043 21511 54049
rect 21453 54040 21465 54043
rect 20588 54012 21465 54040
rect 20588 54000 20594 54012
rect 21453 54009 21465 54012
rect 21499 54009 21511 54043
rect 21453 54003 21511 54009
rect 25038 54000 25044 54052
rect 25096 54040 25102 54052
rect 25409 54043 25467 54049
rect 25409 54040 25421 54043
rect 25096 54012 25421 54040
rect 25096 54000 25102 54012
rect 25409 54009 25421 54012
rect 25455 54009 25467 54043
rect 25409 54003 25467 54009
rect 3786 53932 3792 53984
rect 3844 53932 3850 53984
rect 11701 53975 11759 53981
rect 11701 53941 11713 53975
rect 11747 53972 11759 53975
rect 12710 53972 12716 53984
rect 11747 53944 12716 53972
rect 11747 53941 11759 53944
rect 11701 53935 11759 53941
rect 12710 53932 12716 53944
rect 12768 53932 12774 53984
rect 15286 53932 15292 53984
rect 15344 53972 15350 53984
rect 16117 53975 16175 53981
rect 16117 53972 16129 53975
rect 15344 53944 16129 53972
rect 15344 53932 15350 53944
rect 16117 53941 16129 53944
rect 16163 53941 16175 53975
rect 16117 53935 16175 53941
rect 17494 53932 17500 53984
rect 17552 53932 17558 53984
rect 18598 53932 18604 53984
rect 18656 53932 18662 53984
rect 19334 53932 19340 53984
rect 19392 53972 19398 53984
rect 20073 53975 20131 53981
rect 20073 53972 20085 53975
rect 19392 53944 20085 53972
rect 19392 53932 19398 53944
rect 20073 53941 20085 53944
rect 20119 53941 20131 53975
rect 20073 53935 20131 53941
rect 21174 53932 21180 53984
rect 21232 53932 21238 53984
rect 22094 53932 22100 53984
rect 22152 53972 22158 53984
rect 22649 53975 22707 53981
rect 22649 53972 22661 53975
rect 22152 53944 22661 53972
rect 22152 53932 22158 53944
rect 22649 53941 22661 53944
rect 22695 53941 22707 53975
rect 22649 53935 22707 53941
rect 23750 53932 23756 53984
rect 23808 53932 23814 53984
rect 23842 53932 23848 53984
rect 23900 53972 23906 53984
rect 24765 53975 24823 53981
rect 24765 53972 24777 53975
rect 23900 53944 24777 53972
rect 23900 53932 23906 53944
rect 24765 53941 24777 53944
rect 24811 53941 24823 53975
rect 24765 53935 24823 53941
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 16574 53728 16580 53780
rect 16632 53768 16638 53780
rect 17954 53768 17960 53780
rect 16632 53740 17960 53768
rect 16632 53728 16638 53740
rect 17954 53728 17960 53740
rect 18012 53728 18018 53780
rect 18414 53728 18420 53780
rect 18472 53768 18478 53780
rect 18969 53771 19027 53777
rect 18969 53768 18981 53771
rect 18472 53740 18981 53768
rect 18472 53728 18478 53740
rect 18969 53737 18981 53740
rect 19015 53737 19027 53771
rect 18969 53731 19027 53737
rect 2222 53660 2228 53712
rect 2280 53700 2286 53712
rect 3418 53700 3424 53712
rect 2280 53672 3424 53700
rect 2280 53660 2286 53672
rect 3418 53660 3424 53672
rect 3476 53660 3482 53712
rect 5534 53660 5540 53712
rect 5592 53660 5598 53712
rect 17678 53660 17684 53712
rect 17736 53700 17742 53712
rect 18785 53703 18843 53709
rect 18785 53700 18797 53703
rect 17736 53672 18797 53700
rect 17736 53660 17742 53672
rect 18785 53669 18797 53672
rect 18831 53669 18843 53703
rect 18785 53663 18843 53669
rect 3237 53635 3295 53641
rect 3237 53601 3249 53635
rect 3283 53632 3295 53635
rect 5552 53632 5580 53660
rect 3283 53604 5580 53632
rect 6549 53635 6607 53641
rect 3283 53601 3295 53604
rect 3237 53595 3295 53601
rect 6549 53601 6561 53635
rect 6595 53632 6607 53635
rect 7374 53632 7380 53644
rect 6595 53604 7380 53632
rect 6595 53601 6607 53604
rect 6549 53595 6607 53601
rect 7374 53592 7380 53604
rect 7432 53592 7438 53644
rect 8389 53635 8447 53641
rect 8389 53601 8401 53635
rect 8435 53632 8447 53635
rect 8846 53632 8852 53644
rect 8435 53604 8852 53632
rect 8435 53601 8447 53604
rect 8389 53595 8447 53601
rect 8846 53592 8852 53604
rect 8904 53592 8910 53644
rect 11054 53592 11060 53644
rect 11112 53592 11118 53644
rect 12158 53592 12164 53644
rect 12216 53632 12222 53644
rect 12713 53635 12771 53641
rect 12713 53632 12725 53635
rect 12216 53604 12725 53632
rect 12216 53592 12222 53604
rect 12713 53601 12725 53604
rect 12759 53601 12771 53635
rect 12713 53595 12771 53601
rect 18690 53592 18696 53644
rect 18748 53592 18754 53644
rect 2222 53524 2228 53576
rect 2280 53524 2286 53576
rect 3970 53524 3976 53576
rect 4028 53524 4034 53576
rect 5537 53567 5595 53573
rect 5537 53533 5549 53567
rect 5583 53564 5595 53567
rect 6822 53564 6828 53576
rect 5583 53536 6828 53564
rect 5583 53533 5595 53536
rect 5537 53527 5595 53533
rect 6822 53524 6828 53536
rect 6880 53524 6886 53576
rect 7285 53567 7343 53573
rect 7285 53533 7297 53567
rect 7331 53564 7343 53567
rect 8662 53564 8668 53576
rect 7331 53536 8668 53564
rect 7331 53533 7343 53536
rect 7285 53527 7343 53533
rect 8662 53524 8668 53536
rect 8720 53524 8726 53576
rect 10597 53567 10655 53573
rect 10597 53533 10609 53567
rect 10643 53564 10655 53567
rect 12066 53564 12072 53576
rect 10643 53536 12072 53564
rect 10643 53533 10655 53536
rect 10597 53527 10655 53533
rect 12066 53524 12072 53536
rect 12124 53524 12130 53576
rect 12437 53567 12495 53573
rect 12437 53533 12449 53567
rect 12483 53564 12495 53567
rect 12618 53564 12624 53576
rect 12483 53536 12624 53564
rect 12483 53533 12495 53536
rect 12437 53527 12495 53533
rect 12618 53524 12624 53536
rect 12676 53524 12682 53576
rect 13998 53524 14004 53576
rect 14056 53564 14062 53576
rect 14277 53567 14335 53573
rect 14277 53564 14289 53567
rect 14056 53536 14289 53564
rect 14056 53524 14062 53536
rect 14277 53533 14289 53536
rect 14323 53533 14335 53567
rect 14277 53527 14335 53533
rect 15102 53524 15108 53576
rect 15160 53564 15166 53576
rect 15381 53567 15439 53573
rect 15381 53564 15393 53567
rect 15160 53536 15393 53564
rect 15160 53524 15166 53536
rect 15381 53533 15393 53536
rect 15427 53533 15439 53567
rect 15381 53527 15439 53533
rect 16206 53524 16212 53576
rect 16264 53564 16270 53576
rect 16577 53567 16635 53573
rect 16577 53564 16589 53567
rect 16264 53536 16589 53564
rect 16264 53524 16270 53536
rect 16577 53533 16589 53536
rect 16623 53533 16635 53567
rect 16577 53527 16635 53533
rect 16942 53524 16948 53576
rect 17000 53564 17006 53576
rect 17678 53564 17684 53576
rect 17000 53536 17684 53564
rect 17000 53524 17006 53536
rect 17678 53524 17684 53536
rect 17736 53524 17742 53576
rect 4617 53431 4675 53437
rect 4617 53397 4629 53431
rect 4663 53428 4675 53431
rect 6546 53428 6552 53440
rect 4663 53400 6552 53428
rect 4663 53397 4675 53400
rect 4617 53391 4675 53397
rect 6546 53388 6552 53400
rect 6604 53388 6610 53440
rect 14274 53388 14280 53440
rect 14332 53428 14338 53440
rect 14921 53431 14979 53437
rect 14921 53428 14933 53431
rect 14332 53400 14933 53428
rect 14332 53388 14338 53400
rect 14921 53397 14933 53400
rect 14967 53397 14979 53431
rect 14921 53391 14979 53397
rect 15562 53388 15568 53440
rect 15620 53428 15626 53440
rect 16025 53431 16083 53437
rect 16025 53428 16037 53431
rect 15620 53400 16037 53428
rect 15620 53388 15626 53400
rect 16025 53397 16037 53400
rect 16071 53397 16083 53431
rect 16025 53391 16083 53397
rect 16850 53388 16856 53440
rect 16908 53428 16914 53440
rect 17221 53431 17279 53437
rect 17221 53428 17233 53431
rect 16908 53400 17233 53428
rect 16908 53388 16914 53400
rect 17221 53397 17233 53400
rect 17267 53397 17279 53431
rect 17221 53391 17279 53397
rect 17586 53388 17592 53440
rect 17644 53428 17650 53440
rect 18325 53431 18383 53437
rect 18325 53428 18337 53431
rect 17644 53400 18337 53428
rect 17644 53388 17650 53400
rect 18325 53397 18337 53400
rect 18371 53397 18383 53431
rect 18800 53428 18828 53663
rect 18984 53564 19012 53731
rect 22646 53660 22652 53712
rect 22704 53700 22710 53712
rect 23845 53703 23903 53709
rect 23845 53700 23857 53703
rect 22704 53672 23857 53700
rect 22704 53660 22710 53672
rect 23845 53669 23857 53672
rect 23891 53669 23903 53703
rect 23845 53663 23903 53669
rect 22462 53592 22468 53644
rect 22520 53632 22526 53644
rect 25133 53635 25191 53641
rect 25133 53632 25145 53635
rect 22520 53604 25145 53632
rect 22520 53592 22526 53604
rect 19429 53567 19487 53573
rect 19429 53564 19441 53567
rect 18984 53536 19441 53564
rect 19429 53533 19441 53536
rect 19475 53533 19487 53567
rect 19429 53527 19487 53533
rect 19518 53524 19524 53576
rect 19576 53564 19582 53576
rect 20530 53564 20536 53576
rect 19576 53536 20536 53564
rect 19576 53524 19582 53536
rect 20530 53524 20536 53536
rect 20588 53524 20594 53576
rect 20990 53524 20996 53576
rect 21048 53564 21054 53576
rect 21450 53564 21456 53576
rect 21048 53536 21456 53564
rect 21048 53524 21054 53536
rect 21450 53524 21456 53536
rect 21508 53564 21514 53576
rect 22756 53573 22784 53604
rect 25133 53601 25145 53604
rect 25179 53601 25191 53635
rect 25133 53595 25191 53601
rect 21637 53567 21695 53573
rect 21637 53564 21649 53567
rect 21508 53536 21649 53564
rect 21508 53524 21514 53536
rect 21637 53533 21649 53536
rect 21683 53533 21695 53567
rect 21637 53527 21695 53533
rect 22741 53567 22799 53573
rect 22741 53533 22753 53567
rect 22787 53533 22799 53567
rect 22741 53527 22799 53533
rect 24029 53567 24087 53573
rect 24029 53533 24041 53567
rect 24075 53533 24087 53567
rect 24029 53527 24087 53533
rect 22186 53456 22192 53508
rect 22244 53496 22250 53508
rect 24044 53496 24072 53527
rect 24578 53524 24584 53576
rect 24636 53564 24642 53576
rect 24673 53567 24731 53573
rect 24673 53564 24685 53567
rect 24636 53536 24685 53564
rect 24636 53524 24642 53536
rect 24673 53533 24685 53536
rect 24719 53533 24731 53567
rect 24673 53527 24731 53533
rect 24857 53567 24915 53573
rect 24857 53533 24869 53567
rect 24903 53564 24915 53567
rect 25958 53564 25964 53576
rect 24903 53536 25964 53564
rect 24903 53533 24915 53536
rect 24857 53527 24915 53533
rect 25958 53524 25964 53536
rect 26016 53524 26022 53576
rect 25317 53499 25375 53505
rect 25317 53496 25329 53499
rect 22244 53468 25329 53496
rect 22244 53456 22250 53468
rect 25317 53465 25329 53468
rect 25363 53465 25375 53499
rect 25317 53459 25375 53465
rect 19426 53428 19432 53440
rect 18800 53400 19432 53428
rect 18325 53391 18383 53397
rect 19426 53388 19432 53400
rect 19484 53388 19490 53440
rect 20073 53431 20131 53437
rect 20073 53397 20085 53431
rect 20119 53428 20131 53431
rect 20162 53428 20168 53440
rect 20119 53400 20168 53428
rect 20119 53397 20131 53400
rect 20073 53391 20131 53397
rect 20162 53388 20168 53400
rect 20220 53388 20226 53440
rect 20898 53388 20904 53440
rect 20956 53428 20962 53440
rect 21177 53431 21235 53437
rect 21177 53428 21189 53431
rect 20956 53400 21189 53428
rect 20956 53388 20962 53400
rect 21177 53397 21189 53400
rect 21223 53397 21235 53431
rect 21177 53391 21235 53397
rect 22002 53388 22008 53440
rect 22060 53428 22066 53440
rect 22281 53431 22339 53437
rect 22281 53428 22293 53431
rect 22060 53400 22293 53428
rect 22060 53388 22066 53400
rect 22281 53397 22293 53400
rect 22327 53397 22339 53431
rect 22281 53391 22339 53397
rect 23385 53431 23443 53437
rect 23385 53397 23397 53431
rect 23431 53428 23443 53431
rect 23474 53428 23480 53440
rect 23431 53400 23480 53428
rect 23431 53397 23443 53400
rect 23385 53391 23443 53397
rect 23474 53388 23480 53400
rect 23532 53388 23538 53440
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 11606 53184 11612 53236
rect 11664 53184 11670 53236
rect 17402 53184 17408 53236
rect 17460 53184 17466 53236
rect 17678 53184 17684 53236
rect 17736 53184 17742 53236
rect 3973 53159 4031 53165
rect 3973 53125 3985 53159
rect 4019 53156 4031 53159
rect 4430 53156 4436 53168
rect 4019 53128 4436 53156
rect 4019 53125 4031 53128
rect 3973 53119 4031 53125
rect 4430 53116 4436 53128
rect 4488 53116 4494 53168
rect 5813 53159 5871 53165
rect 5813 53125 5825 53159
rect 5859 53156 5871 53159
rect 6270 53156 6276 53168
rect 5859 53128 6276 53156
rect 5859 53125 5871 53128
rect 5813 53119 5871 53125
rect 6270 53116 6276 53128
rect 6328 53116 6334 53168
rect 9125 53159 9183 53165
rect 9125 53125 9137 53159
rect 9171 53156 9183 53159
rect 9214 53156 9220 53168
rect 9171 53128 9220 53156
rect 9171 53125 9183 53128
rect 9125 53119 9183 53125
rect 9214 53116 9220 53128
rect 9272 53116 9278 53168
rect 13354 53116 13360 53168
rect 13412 53156 13418 53168
rect 16025 53159 16083 53165
rect 13412 53128 14872 53156
rect 13412 53116 13418 53128
rect 14844 53100 14872 53128
rect 16025 53125 16037 53159
rect 16071 53156 16083 53159
rect 17494 53156 17500 53168
rect 16071 53128 17500 53156
rect 16071 53125 16083 53128
rect 16025 53119 16083 53125
rect 17494 53116 17500 53128
rect 17552 53116 17558 53168
rect 18598 53156 18604 53168
rect 17696 53128 18604 53156
rect 1673 53091 1731 53097
rect 1673 53057 1685 53091
rect 1719 53057 1731 53091
rect 1673 53051 1731 53057
rect 2961 53091 3019 53097
rect 2961 53057 2973 53091
rect 3007 53088 3019 53091
rect 4522 53088 4528 53100
rect 3007 53060 4528 53088
rect 3007 53057 3019 53060
rect 2961 53051 3019 53057
rect 1688 52952 1716 53051
rect 4522 53048 4528 53060
rect 4580 53048 4586 53100
rect 4706 53048 4712 53100
rect 4764 53048 4770 53100
rect 6546 53048 6552 53100
rect 6604 53048 6610 53100
rect 7558 53048 7564 53100
rect 7616 53088 7622 53100
rect 7929 53091 7987 53097
rect 7929 53088 7941 53091
rect 7616 53060 7941 53088
rect 7616 53048 7622 53060
rect 7929 53057 7941 53060
rect 7975 53057 7987 53091
rect 7929 53051 7987 53057
rect 9306 53048 9312 53100
rect 9364 53088 9370 53100
rect 9769 53091 9827 53097
rect 9769 53088 9781 53091
rect 9364 53060 9781 53088
rect 9364 53048 9370 53060
rect 9769 53057 9781 53060
rect 9815 53057 9827 53091
rect 9769 53051 9827 53057
rect 11882 53048 11888 53100
rect 11940 53048 11946 53100
rect 13630 53048 13636 53100
rect 13688 53088 13694 53100
rect 13725 53091 13783 53097
rect 13725 53088 13737 53091
rect 13688 53060 13737 53088
rect 13688 53048 13694 53060
rect 13725 53057 13737 53060
rect 13771 53057 13783 53091
rect 13725 53051 13783 53057
rect 14826 53048 14832 53100
rect 14884 53048 14890 53100
rect 16853 53091 16911 53097
rect 16853 53057 16865 53091
rect 16899 53088 16911 53091
rect 17696 53088 17724 53128
rect 18598 53116 18604 53128
rect 18656 53116 18662 53168
rect 19334 53116 19340 53168
rect 19392 53116 19398 53168
rect 23750 53156 23756 53168
rect 22756 53128 23756 53156
rect 16899 53060 17724 53088
rect 17865 53091 17923 53097
rect 16899 53057 16911 53060
rect 16853 53051 16911 53057
rect 17865 53057 17877 53091
rect 17911 53088 17923 53091
rect 18141 53091 18199 53097
rect 18141 53088 18153 53091
rect 17911 53060 18153 53088
rect 17911 53057 17923 53060
rect 17865 53051 17923 53057
rect 18141 53057 18153 53060
rect 18187 53088 18199 53091
rect 18322 53088 18328 53100
rect 18187 53060 18328 53088
rect 18187 53057 18199 53060
rect 18141 53051 18199 53057
rect 18322 53048 18328 53060
rect 18380 53048 18386 53100
rect 19886 53048 19892 53100
rect 19944 53088 19950 53100
rect 20073 53091 20131 53097
rect 20073 53088 20085 53091
rect 19944 53060 20085 53088
rect 19944 53048 19950 53060
rect 20073 53057 20085 53060
rect 20119 53057 20131 53091
rect 20073 53051 20131 53057
rect 20717 53091 20775 53097
rect 20717 53057 20729 53091
rect 20763 53088 20775 53091
rect 21269 53091 21327 53097
rect 21269 53088 21281 53091
rect 20763 53060 21281 53088
rect 20763 53057 20775 53060
rect 20717 53051 20775 53057
rect 21269 53057 21281 53060
rect 21315 53057 21327 53091
rect 21269 53051 21327 53057
rect 22002 53048 22008 53100
rect 22060 53048 22066 53100
rect 22756 53097 22784 53128
rect 23750 53116 23756 53128
rect 23808 53116 23814 53168
rect 22741 53091 22799 53097
rect 22741 53057 22753 53091
rect 22787 53057 22799 53091
rect 22741 53051 22799 53057
rect 23474 53048 23480 53100
rect 23532 53048 23538 53100
rect 24305 53091 24363 53097
rect 24305 53057 24317 53091
rect 24351 53088 24363 53091
rect 24762 53088 24768 53100
rect 24351 53060 24768 53088
rect 24351 53057 24363 53060
rect 24305 53051 24363 53057
rect 24762 53048 24768 53060
rect 24820 53048 24826 53100
rect 25038 53048 25044 53100
rect 25096 53048 25102 53100
rect 10318 52980 10324 53032
rect 10376 52980 10382 53032
rect 11790 52980 11796 53032
rect 11848 53020 11854 53032
rect 12345 53023 12403 53029
rect 12345 53020 12357 53023
rect 11848 52992 12357 53020
rect 11848 52980 11854 52992
rect 12345 52989 12357 52992
rect 12391 52989 12403 53023
rect 12345 52983 12403 52989
rect 7193 52955 7251 52961
rect 7193 52952 7205 52955
rect 1688 52924 7205 52952
rect 7193 52921 7205 52924
rect 7239 52921 7251 52955
rect 7193 52915 7251 52921
rect 16209 52955 16267 52961
rect 16209 52921 16221 52955
rect 16255 52952 16267 52955
rect 16390 52952 16396 52964
rect 16255 52924 16396 52952
rect 16255 52921 16267 52924
rect 16209 52915 16267 52921
rect 16390 52912 16396 52924
rect 16448 52912 16454 52964
rect 21453 52955 21511 52961
rect 21453 52921 21465 52955
rect 21499 52952 21511 52955
rect 21634 52952 21640 52964
rect 21499 52924 21640 52952
rect 21499 52921 21511 52924
rect 21453 52915 21511 52921
rect 21634 52912 21640 52924
rect 21692 52912 21698 52964
rect 22189 52955 22247 52961
rect 22189 52921 22201 52955
rect 22235 52952 22247 52955
rect 22738 52952 22744 52964
rect 22235 52924 22744 52952
rect 22235 52921 22247 52924
rect 22189 52915 22247 52921
rect 22738 52912 22744 52924
rect 22796 52912 22802 52964
rect 1762 52844 1768 52896
rect 1820 52884 1826 52896
rect 2317 52887 2375 52893
rect 2317 52884 2329 52887
rect 1820 52856 2329 52884
rect 1820 52844 1826 52856
rect 2317 52853 2329 52856
rect 2363 52853 2375 52887
rect 2317 52847 2375 52853
rect 14366 52844 14372 52896
rect 14424 52844 14430 52896
rect 14550 52844 14556 52896
rect 14608 52884 14614 52896
rect 15473 52887 15531 52893
rect 15473 52884 15485 52887
rect 14608 52856 15485 52884
rect 14608 52844 14614 52856
rect 15473 52853 15485 52856
rect 15519 52853 15531 52887
rect 15473 52847 15531 52853
rect 17034 52844 17040 52896
rect 17092 52844 17098 52896
rect 18782 52844 18788 52896
rect 18840 52844 18846 52896
rect 19426 52844 19432 52896
rect 19484 52844 19490 52896
rect 22554 52844 22560 52896
rect 22612 52884 22618 52896
rect 22925 52887 22983 52893
rect 22925 52884 22937 52887
rect 22612 52856 22937 52884
rect 22612 52844 22618 52856
rect 22925 52853 22937 52856
rect 22971 52853 22983 52887
rect 22925 52847 22983 52853
rect 23658 52844 23664 52896
rect 23716 52844 23722 52896
rect 23934 52844 23940 52896
rect 23992 52884 23998 52896
rect 24489 52887 24547 52893
rect 24489 52884 24501 52887
rect 23992 52856 24501 52884
rect 23992 52844 23998 52856
rect 24489 52853 24501 52856
rect 24535 52853 24547 52887
rect 24489 52847 24547 52853
rect 24946 52844 24952 52896
rect 25004 52884 25010 52896
rect 25225 52887 25283 52893
rect 25225 52884 25237 52887
rect 25004 52856 25237 52884
rect 25004 52844 25010 52856
rect 25225 52853 25237 52856
rect 25271 52853 25283 52887
rect 25225 52847 25283 52853
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 1854 52640 1860 52692
rect 1912 52680 1918 52692
rect 3510 52680 3516 52692
rect 1912 52652 3516 52680
rect 1912 52640 1918 52652
rect 3510 52640 3516 52652
rect 3568 52640 3574 52692
rect 12618 52640 12624 52692
rect 12676 52640 12682 52692
rect 14826 52640 14832 52692
rect 14884 52640 14890 52692
rect 15102 52640 15108 52692
rect 15160 52680 15166 52692
rect 15197 52683 15255 52689
rect 15197 52680 15209 52683
rect 15160 52652 15209 52680
rect 15160 52640 15166 52652
rect 15197 52649 15209 52652
rect 15243 52649 15255 52683
rect 15197 52643 15255 52649
rect 16206 52640 16212 52692
rect 16264 52680 16270 52692
rect 16393 52683 16451 52689
rect 16393 52680 16405 52683
rect 16264 52652 16405 52680
rect 16264 52640 16270 52652
rect 16393 52649 16405 52652
rect 16439 52649 16451 52683
rect 16393 52643 16451 52649
rect 17037 52683 17095 52689
rect 17037 52649 17049 52683
rect 17083 52680 17095 52683
rect 17126 52680 17132 52692
rect 17083 52652 17132 52680
rect 17083 52649 17095 52652
rect 17037 52643 17095 52649
rect 17126 52640 17132 52652
rect 17184 52640 17190 52692
rect 21358 52640 21364 52692
rect 21416 52680 21422 52692
rect 22373 52683 22431 52689
rect 22373 52680 22385 52683
rect 21416 52652 22385 52680
rect 21416 52640 21422 52652
rect 22373 52649 22385 52652
rect 22419 52649 22431 52683
rect 22373 52643 22431 52649
rect 24026 52640 24032 52692
rect 24084 52640 24090 52692
rect 24213 52683 24271 52689
rect 24213 52649 24225 52683
rect 24259 52680 24271 52683
rect 24578 52680 24584 52692
rect 24259 52652 24584 52680
rect 24259 52649 24271 52652
rect 24213 52643 24271 52649
rect 24578 52640 24584 52652
rect 24636 52640 24642 52692
rect 24762 52640 24768 52692
rect 24820 52640 24826 52692
rect 1302 52572 1308 52624
rect 1360 52612 1366 52624
rect 3786 52612 3792 52624
rect 1360 52584 3792 52612
rect 1360 52572 1366 52584
rect 3786 52572 3792 52584
rect 3844 52612 3850 52624
rect 3844 52584 4016 52612
rect 3844 52572 3850 52584
rect 3237 52547 3295 52553
rect 3237 52513 3249 52547
rect 3283 52544 3295 52547
rect 3694 52544 3700 52556
rect 3283 52516 3700 52544
rect 3283 52513 3295 52516
rect 3237 52507 3295 52513
rect 3694 52504 3700 52516
rect 3752 52504 3758 52556
rect 3988 52553 4016 52584
rect 15654 52572 15660 52624
rect 15712 52612 15718 52624
rect 17773 52615 17831 52621
rect 17773 52612 17785 52615
rect 15712 52584 17785 52612
rect 15712 52572 15718 52584
rect 17773 52581 17785 52584
rect 17819 52581 17831 52615
rect 17773 52575 17831 52581
rect 21542 52572 21548 52624
rect 21600 52612 21606 52624
rect 21821 52615 21879 52621
rect 21821 52612 21833 52615
rect 21600 52584 21833 52612
rect 21600 52572 21606 52584
rect 21821 52581 21833 52584
rect 21867 52581 21879 52615
rect 21821 52575 21879 52581
rect 22462 52572 22468 52624
rect 22520 52612 22526 52624
rect 23293 52615 23351 52621
rect 23293 52612 23305 52615
rect 22520 52584 23305 52612
rect 22520 52572 22526 52584
rect 23293 52581 23305 52584
rect 23339 52581 23351 52615
rect 23293 52575 23351 52581
rect 25130 52572 25136 52624
rect 25188 52612 25194 52624
rect 25225 52615 25283 52621
rect 25225 52612 25237 52615
rect 25188 52584 25237 52612
rect 25188 52572 25194 52584
rect 25225 52581 25237 52584
rect 25271 52581 25283 52615
rect 25225 52575 25283 52581
rect 3973 52547 4031 52553
rect 3973 52513 3985 52547
rect 4019 52513 4031 52547
rect 3973 52507 4031 52513
rect 4249 52547 4307 52553
rect 4249 52513 4261 52547
rect 4295 52544 4307 52547
rect 4295 52516 7696 52544
rect 4295 52513 4307 52516
rect 4249 52507 4307 52513
rect 2225 52479 2283 52485
rect 2225 52445 2237 52479
rect 2271 52476 2283 52479
rect 5166 52476 5172 52488
rect 2271 52448 5172 52476
rect 2271 52445 2283 52448
rect 2225 52439 2283 52445
rect 5166 52436 5172 52448
rect 5224 52436 5230 52488
rect 5445 52479 5503 52485
rect 5445 52445 5457 52479
rect 5491 52476 5503 52479
rect 5902 52476 5908 52488
rect 5491 52448 5908 52476
rect 5491 52445 5503 52448
rect 5445 52439 5503 52445
rect 5902 52436 5908 52448
rect 5960 52436 5966 52488
rect 6549 52479 6607 52485
rect 6549 52445 6561 52479
rect 6595 52476 6607 52479
rect 6638 52476 6644 52488
rect 6595 52448 6644 52476
rect 6595 52445 6607 52448
rect 6549 52439 6607 52445
rect 6638 52436 6644 52448
rect 6696 52436 6702 52488
rect 7282 52436 7288 52488
rect 7340 52436 7346 52488
rect 7668 52476 7696 52516
rect 7742 52504 7748 52556
rect 7800 52504 7806 52556
rect 10686 52504 10692 52556
rect 10744 52544 10750 52556
rect 11241 52547 11299 52553
rect 11241 52544 11253 52547
rect 10744 52516 11253 52544
rect 10744 52504 10750 52516
rect 11241 52513 11253 52516
rect 11287 52513 11299 52547
rect 21174 52544 21180 52556
rect 11241 52507 11299 52513
rect 19444 52516 21180 52544
rect 8570 52476 8576 52488
rect 7668 52448 8576 52476
rect 8570 52436 8576 52448
rect 8628 52436 8634 52488
rect 9582 52436 9588 52488
rect 9640 52476 9646 52488
rect 10781 52479 10839 52485
rect 10781 52476 10793 52479
rect 9640 52448 10793 52476
rect 9640 52436 9646 52448
rect 10781 52445 10793 52448
rect 10827 52445 10839 52479
rect 10781 52439 10839 52445
rect 12802 52436 12808 52488
rect 12860 52436 12866 52488
rect 13538 52436 13544 52488
rect 13596 52476 13602 52488
rect 13633 52479 13691 52485
rect 13633 52476 13645 52479
rect 13596 52448 13645 52476
rect 13596 52436 13602 52448
rect 13633 52445 13645 52448
rect 13679 52445 13691 52479
rect 13633 52439 13691 52445
rect 14274 52436 14280 52488
rect 14332 52436 14338 52488
rect 15562 52436 15568 52488
rect 15620 52436 15626 52488
rect 16850 52436 16856 52488
rect 16908 52436 16914 52488
rect 17586 52436 17592 52488
rect 17644 52436 17650 52488
rect 18417 52479 18475 52485
rect 18417 52445 18429 52479
rect 18463 52476 18475 52479
rect 18782 52476 18788 52488
rect 18463 52448 18788 52476
rect 18463 52445 18475 52448
rect 18417 52439 18475 52445
rect 18782 52436 18788 52448
rect 18840 52436 18846 52488
rect 19444 52485 19472 52516
rect 21174 52504 21180 52516
rect 21232 52504 21238 52556
rect 21726 52504 21732 52556
rect 21784 52544 21790 52556
rect 22833 52547 22891 52553
rect 22833 52544 22845 52547
rect 21784 52516 22845 52544
rect 21784 52504 21790 52516
rect 19429 52479 19487 52485
rect 19429 52445 19441 52479
rect 19475 52445 19487 52479
rect 19429 52439 19487 52445
rect 20162 52436 20168 52488
rect 20220 52436 20226 52488
rect 20898 52436 20904 52488
rect 20956 52436 20962 52488
rect 21637 52479 21695 52485
rect 21637 52445 21649 52479
rect 21683 52476 21695 52479
rect 22094 52476 22100 52488
rect 21683 52448 22100 52476
rect 21683 52445 21695 52448
rect 21637 52439 21695 52445
rect 22094 52436 22100 52448
rect 22152 52436 22158 52488
rect 22572 52485 22600 52516
rect 22833 52513 22845 52516
rect 22879 52513 22891 52547
rect 22833 52507 22891 52513
rect 22557 52479 22615 52485
rect 22557 52445 22569 52479
rect 22603 52445 22615 52479
rect 22557 52439 22615 52445
rect 22738 52436 22744 52488
rect 22796 52476 22802 52488
rect 22922 52476 22928 52488
rect 22796 52448 22928 52476
rect 22796 52436 22802 52448
rect 22922 52436 22928 52448
rect 22980 52436 22986 52488
rect 23290 52436 23296 52488
rect 23348 52476 23354 52488
rect 23477 52479 23535 52485
rect 23477 52476 23489 52479
rect 23348 52448 23489 52476
rect 23348 52436 23354 52448
rect 23477 52445 23489 52448
rect 23523 52476 23535 52479
rect 23753 52479 23811 52485
rect 23753 52476 23765 52479
rect 23523 52448 23765 52476
rect 23523 52445 23535 52448
rect 23477 52439 23535 52445
rect 23753 52445 23765 52448
rect 23799 52445 23811 52479
rect 23753 52439 23811 52445
rect 24581 52479 24639 52485
rect 24581 52445 24593 52479
rect 24627 52476 24639 52479
rect 24762 52476 24768 52488
rect 24627 52448 24768 52476
rect 24627 52445 24639 52448
rect 24581 52439 24639 52445
rect 24762 52436 24768 52448
rect 24820 52476 24826 52488
rect 25041 52479 25099 52485
rect 25041 52476 25053 52479
rect 24820 52448 25053 52476
rect 24820 52436 24826 52448
rect 25041 52445 25053 52448
rect 25087 52445 25099 52479
rect 25041 52439 25099 52445
rect 13449 52411 13507 52417
rect 13449 52377 13461 52411
rect 13495 52408 13507 52411
rect 14550 52408 14556 52420
rect 13495 52380 14556 52408
rect 13495 52377 13507 52380
rect 13449 52371 13507 52377
rect 14550 52368 14556 52380
rect 14608 52368 14614 52420
rect 14458 52300 14464 52352
rect 14516 52300 14522 52352
rect 15746 52300 15752 52352
rect 15804 52300 15810 52352
rect 18506 52300 18512 52352
rect 18564 52300 18570 52352
rect 19610 52300 19616 52352
rect 19668 52300 19674 52352
rect 20346 52300 20352 52352
rect 20404 52300 20410 52352
rect 21082 52300 21088 52352
rect 21140 52300 21146 52352
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 4522 52096 4528 52148
rect 4580 52136 4586 52148
rect 7009 52139 7067 52145
rect 7009 52136 7021 52139
rect 4580 52108 7021 52136
rect 4580 52096 4586 52108
rect 7009 52105 7021 52108
rect 7055 52105 7067 52139
rect 7009 52099 7067 52105
rect 11701 52139 11759 52145
rect 11701 52105 11713 52139
rect 11747 52136 11759 52139
rect 11882 52136 11888 52148
rect 11747 52108 11888 52136
rect 11747 52105 11759 52108
rect 11701 52099 11759 52105
rect 11882 52096 11888 52108
rect 11940 52096 11946 52148
rect 12342 52096 12348 52148
rect 12400 52096 12406 52148
rect 19886 52096 19892 52148
rect 19944 52096 19950 52148
rect 21450 52096 21456 52148
rect 21508 52096 21514 52148
rect 6917 52071 6975 52077
rect 6917 52037 6929 52071
rect 6963 52068 6975 52071
rect 9122 52068 9128 52080
rect 6963 52040 9128 52068
rect 6963 52037 6975 52040
rect 6917 52031 6975 52037
rect 9122 52028 9128 52040
rect 9180 52028 9186 52080
rect 13817 52071 13875 52077
rect 13817 52037 13829 52071
rect 13863 52068 13875 52071
rect 14366 52068 14372 52080
rect 13863 52040 14372 52068
rect 13863 52037 13875 52040
rect 13817 52031 13875 52037
rect 14366 52028 14372 52040
rect 14424 52028 14430 52080
rect 1670 51960 1676 52012
rect 1728 51960 1734 52012
rect 2961 52003 3019 52009
rect 2961 51969 2973 52003
rect 3007 52000 3019 52003
rect 4801 52003 4859 52009
rect 3007 51972 3832 52000
rect 3007 51969 3019 51972
rect 2961 51963 3019 51969
rect 3326 51892 3332 51944
rect 3384 51892 3390 51944
rect 3804 51864 3832 51972
rect 4801 51969 4813 52003
rect 4847 52000 4859 52003
rect 7190 52000 7196 52012
rect 4847 51972 7196 52000
rect 4847 51969 4859 51972
rect 4801 51963 4859 51969
rect 7190 51960 7196 51972
rect 7248 51960 7254 52012
rect 8021 52003 8079 52009
rect 8021 51969 8033 52003
rect 8067 51969 8079 52003
rect 8021 51963 8079 51969
rect 4890 51892 4896 51944
rect 4948 51932 4954 51944
rect 5077 51935 5135 51941
rect 5077 51932 5089 51935
rect 4948 51904 5089 51932
rect 4948 51892 4954 51904
rect 5077 51901 5089 51904
rect 5123 51901 5135 51935
rect 5077 51895 5135 51901
rect 8036 51864 8064 51963
rect 9674 51960 9680 52012
rect 9732 51960 9738 52012
rect 10870 51960 10876 52012
rect 10928 52000 10934 52012
rect 11885 52003 11943 52009
rect 11885 52000 11897 52003
rect 10928 51972 11897 52000
rect 10928 51960 10934 51972
rect 11885 51969 11897 51972
rect 11931 51969 11943 52003
rect 11885 51963 11943 51969
rect 11974 51960 11980 52012
rect 12032 52000 12038 52012
rect 12529 52003 12587 52009
rect 12529 52000 12541 52003
rect 12032 51972 12541 52000
rect 12032 51960 12038 51972
rect 12529 51969 12541 51972
rect 12575 51969 12587 52003
rect 12529 51963 12587 51969
rect 14642 51960 14648 52012
rect 14700 52000 14706 52012
rect 14921 52003 14979 52009
rect 14921 52000 14933 52003
rect 14700 51972 14933 52000
rect 14700 51960 14706 51972
rect 14921 51969 14933 51972
rect 14967 51969 14979 52003
rect 14921 51963 14979 51969
rect 15838 51960 15844 52012
rect 15896 52000 15902 52012
rect 16117 52003 16175 52009
rect 16117 52000 16129 52003
rect 15896 51972 16129 52000
rect 15896 51960 15902 51972
rect 16117 51969 16129 51972
rect 16163 52000 16175 52003
rect 16393 52003 16451 52009
rect 16393 52000 16405 52003
rect 16163 51972 16405 52000
rect 16163 51969 16175 51972
rect 16117 51963 16175 51969
rect 16393 51969 16405 51972
rect 16439 51969 16451 52003
rect 16393 51963 16451 51969
rect 17310 51960 17316 52012
rect 17368 52000 17374 52012
rect 17589 52003 17647 52009
rect 17589 52000 17601 52003
rect 17368 51972 17601 52000
rect 17368 51960 17374 51972
rect 17589 51969 17601 51972
rect 17635 52000 17647 52003
rect 17865 52003 17923 52009
rect 17865 52000 17877 52003
rect 17635 51972 17877 52000
rect 17635 51969 17647 51972
rect 17589 51963 17647 51969
rect 17865 51969 17877 51972
rect 17911 51969 17923 52003
rect 17865 51963 17923 51969
rect 18874 51960 18880 52012
rect 18932 52000 18938 52012
rect 19061 52003 19119 52009
rect 19061 52000 19073 52003
rect 18932 51972 19073 52000
rect 18932 51960 18938 51972
rect 19061 51969 19073 51972
rect 19107 52000 19119 52003
rect 19337 52003 19395 52009
rect 19337 52000 19349 52003
rect 19107 51972 19349 52000
rect 19107 51969 19119 51972
rect 19061 51963 19119 51969
rect 19337 51969 19349 51972
rect 19383 51969 19395 52003
rect 19337 51963 19395 51969
rect 20254 51960 20260 52012
rect 20312 52000 20318 52012
rect 20533 52003 20591 52009
rect 20533 52000 20545 52003
rect 20312 51972 20545 52000
rect 20312 51960 20318 51972
rect 20533 51969 20545 51972
rect 20579 52000 20591 52003
rect 20809 52003 20867 52009
rect 20809 52000 20821 52003
rect 20579 51972 20821 52000
rect 20579 51969 20591 51972
rect 20533 51963 20591 51969
rect 20809 51969 20821 51972
rect 20855 51969 20867 52003
rect 20809 51963 20867 51969
rect 22830 51960 22836 52012
rect 22888 52000 22894 52012
rect 23293 52003 23351 52009
rect 23293 52000 23305 52003
rect 22888 51972 23305 52000
rect 22888 51960 22894 51972
rect 23293 51969 23305 51972
rect 23339 52000 23351 52003
rect 23569 52003 23627 52009
rect 23569 52000 23581 52003
rect 23339 51972 23581 52000
rect 23339 51969 23351 51972
rect 23293 51963 23351 51969
rect 23569 51969 23581 51972
rect 23615 51969 23627 52003
rect 23569 51963 23627 51969
rect 23658 51960 23664 52012
rect 23716 52000 23722 52012
rect 24121 52003 24179 52009
rect 24121 52000 24133 52003
rect 23716 51972 24133 52000
rect 23716 51960 23722 51972
rect 24121 51969 24133 51972
rect 24167 52000 24179 52003
rect 24397 52003 24455 52009
rect 24397 52000 24409 52003
rect 24167 51972 24409 52000
rect 24167 51969 24179 51972
rect 24121 51963 24179 51969
rect 24397 51969 24409 51972
rect 24443 51969 24455 52003
rect 24397 51963 24455 51969
rect 24670 51960 24676 52012
rect 24728 52000 24734 52012
rect 25041 52003 25099 52009
rect 25041 52000 25053 52003
rect 24728 51972 25053 52000
rect 24728 51960 24734 51972
rect 25041 51969 25053 51972
rect 25087 51969 25099 52003
rect 25041 51963 25099 51969
rect 8478 51892 8484 51944
rect 8536 51892 8542 51944
rect 9766 51892 9772 51944
rect 9824 51932 9830 51944
rect 10137 51935 10195 51941
rect 10137 51932 10149 51935
rect 9824 51904 10149 51932
rect 9824 51892 9830 51904
rect 10137 51901 10149 51904
rect 10183 51901 10195 51935
rect 10137 51895 10195 51901
rect 10410 51864 10416 51876
rect 3804 51836 4936 51864
rect 8036 51836 10416 51864
rect 4908 51808 4936 51836
rect 10410 51824 10416 51836
rect 10468 51824 10474 51876
rect 14001 51867 14059 51873
rect 14001 51833 14013 51867
rect 14047 51864 14059 51867
rect 14090 51864 14096 51876
rect 14047 51836 14096 51864
rect 14047 51833 14059 51836
rect 14001 51827 14059 51833
rect 14090 51824 14096 51836
rect 14148 51824 14154 51876
rect 14461 51867 14519 51873
rect 14461 51833 14473 51867
rect 14507 51864 14519 51867
rect 15010 51864 15016 51876
rect 14507 51836 15016 51864
rect 14507 51833 14519 51836
rect 14461 51827 14519 51833
rect 15010 51824 15016 51836
rect 15068 51824 15074 51876
rect 15933 51867 15991 51873
rect 15933 51833 15945 51867
rect 15979 51864 15991 51867
rect 17218 51864 17224 51876
rect 15979 51836 17224 51864
rect 15979 51833 15991 51836
rect 15933 51827 15991 51833
rect 17218 51824 17224 51836
rect 17276 51824 17282 51876
rect 17405 51867 17463 51873
rect 17405 51833 17417 51867
rect 17451 51864 17463 51867
rect 18414 51864 18420 51876
rect 17451 51836 18420 51864
rect 17451 51833 17463 51836
rect 17405 51827 17463 51833
rect 18414 51824 18420 51836
rect 18472 51824 18478 51876
rect 22738 51824 22744 51876
rect 22796 51864 22802 51876
rect 23937 51867 23995 51873
rect 23937 51864 23949 51867
rect 22796 51836 23949 51864
rect 22796 51824 22802 51836
rect 23937 51833 23949 51836
rect 23983 51833 23995 51867
rect 23937 51827 23995 51833
rect 2317 51799 2375 51805
rect 2317 51765 2329 51799
rect 2363 51796 2375 51799
rect 3970 51796 3976 51808
rect 2363 51768 3976 51796
rect 2363 51765 2375 51768
rect 2317 51759 2375 51765
rect 3970 51756 3976 51768
rect 4028 51756 4034 51808
rect 4890 51756 4896 51808
rect 4948 51756 4954 51808
rect 18598 51756 18604 51808
rect 18656 51796 18662 51808
rect 18877 51799 18935 51805
rect 18877 51796 18889 51799
rect 18656 51768 18889 51796
rect 18656 51756 18662 51768
rect 18877 51765 18889 51768
rect 18923 51765 18935 51799
rect 18877 51759 18935 51765
rect 20162 51756 20168 51808
rect 20220 51796 20226 51808
rect 20349 51799 20407 51805
rect 20349 51796 20361 51799
rect 20220 51768 20361 51796
rect 20220 51756 20226 51768
rect 20349 51765 20361 51768
rect 20395 51765 20407 51799
rect 20349 51759 20407 51765
rect 22370 51756 22376 51808
rect 22428 51796 22434 51808
rect 23109 51799 23167 51805
rect 23109 51796 23121 51799
rect 22428 51768 23121 51796
rect 22428 51756 22434 51768
rect 23109 51765 23121 51768
rect 23155 51765 23167 51799
rect 23109 51759 23167 51765
rect 25225 51799 25283 51805
rect 25225 51765 25237 51799
rect 25271 51796 25283 51799
rect 25774 51796 25780 51808
rect 25271 51768 25780 51796
rect 25271 51765 25283 51768
rect 25225 51759 25283 51765
rect 25774 51756 25780 51768
rect 25832 51756 25838 51808
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 9950 51552 9956 51604
rect 10008 51592 10014 51604
rect 10229 51595 10287 51601
rect 10229 51592 10241 51595
rect 10008 51564 10241 51592
rect 10008 51552 10014 51564
rect 10229 51561 10241 51564
rect 10275 51561 10287 51595
rect 10229 51555 10287 51561
rect 2866 51416 2872 51468
rect 2924 51416 2930 51468
rect 6914 51456 6920 51468
rect 3896 51428 6920 51456
rect 2225 51391 2283 51397
rect 2225 51357 2237 51391
rect 2271 51388 2283 51391
rect 3896 51388 3924 51428
rect 6914 51416 6920 51428
rect 6972 51416 6978 51468
rect 7006 51416 7012 51468
rect 7064 51456 7070 51468
rect 7561 51459 7619 51465
rect 7561 51456 7573 51459
rect 7064 51428 7573 51456
rect 7064 51416 7070 51428
rect 7561 51425 7573 51428
rect 7607 51425 7619 51459
rect 7561 51419 7619 51425
rect 2271 51360 3924 51388
rect 2271 51357 2283 51360
rect 2225 51351 2283 51357
rect 3970 51348 3976 51400
rect 4028 51348 4034 51400
rect 5445 51391 5503 51397
rect 5445 51357 5457 51391
rect 5491 51357 5503 51391
rect 5445 51351 5503 51357
rect 5460 51320 5488 51351
rect 5534 51348 5540 51400
rect 5592 51388 5598 51400
rect 6181 51391 6239 51397
rect 6181 51388 6193 51391
rect 5592 51360 6193 51388
rect 5592 51348 5598 51360
rect 6181 51357 6193 51360
rect 6227 51357 6239 51391
rect 6181 51351 6239 51357
rect 7098 51348 7104 51400
rect 7156 51348 7162 51400
rect 9214 51348 9220 51400
rect 9272 51388 9278 51400
rect 10413 51391 10471 51397
rect 10413 51388 10425 51391
rect 9272 51360 10425 51388
rect 9272 51348 9278 51360
rect 10413 51357 10425 51360
rect 10459 51357 10471 51391
rect 10413 51351 10471 51357
rect 24765 51391 24823 51397
rect 24765 51357 24777 51391
rect 24811 51388 24823 51391
rect 25038 51388 25044 51400
rect 24811 51360 25044 51388
rect 24811 51357 24823 51360
rect 24765 51351 24823 51357
rect 25038 51348 25044 51360
rect 25096 51348 25102 51400
rect 6730 51320 6736 51332
rect 5460 51292 6736 51320
rect 6730 51280 6736 51292
rect 6788 51280 6794 51332
rect 7006 51280 7012 51332
rect 7064 51320 7070 51332
rect 7190 51320 7196 51332
rect 7064 51292 7196 51320
rect 7064 51280 7070 51292
rect 7190 51280 7196 51292
rect 7248 51280 7254 51332
rect 4246 51212 4252 51264
rect 4304 51252 4310 51264
rect 4617 51255 4675 51261
rect 4617 51252 4629 51255
rect 4304 51224 4629 51252
rect 4304 51212 4310 51224
rect 4617 51221 4629 51224
rect 4663 51221 4675 51255
rect 4617 51215 4675 51221
rect 25225 51255 25283 51261
rect 25225 51221 25237 51255
rect 25271 51252 25283 51255
rect 25866 51252 25872 51264
rect 25271 51224 25872 51252
rect 25271 51221 25283 51224
rect 25225 51215 25283 51221
rect 25866 51212 25872 51224
rect 25924 51212 25930 51264
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 1581 51051 1639 51057
rect 1581 51017 1593 51051
rect 1627 51048 1639 51051
rect 1670 51048 1676 51060
rect 1627 51020 1676 51048
rect 1627 51017 1639 51020
rect 1581 51011 1639 51017
rect 1670 51008 1676 51020
rect 1728 51008 1734 51060
rect 6914 51008 6920 51060
rect 6972 51008 6978 51060
rect 2314 50940 2320 50992
rect 2372 50980 2378 50992
rect 2372 50952 7788 50980
rect 2372 50940 2378 50952
rect 1762 50872 1768 50924
rect 1820 50872 1826 50924
rect 2501 50915 2559 50921
rect 2501 50881 2513 50915
rect 2547 50912 2559 50915
rect 4249 50915 4307 50921
rect 2547 50884 2912 50912
rect 2547 50881 2559 50884
rect 2501 50875 2559 50881
rect 2774 50804 2780 50856
rect 2832 50804 2838 50856
rect 2884 50776 2912 50884
rect 4249 50881 4261 50915
rect 4295 50912 4307 50915
rect 5442 50912 5448 50924
rect 4295 50884 5448 50912
rect 4295 50881 4307 50884
rect 4249 50875 4307 50881
rect 5442 50872 5448 50884
rect 5500 50872 5506 50924
rect 6825 50915 6883 50921
rect 6825 50881 6837 50915
rect 6871 50912 6883 50915
rect 7650 50912 7656 50924
rect 6871 50884 7656 50912
rect 6871 50881 6883 50884
rect 6825 50875 6883 50881
rect 7650 50872 7656 50884
rect 7708 50872 7714 50924
rect 7760 50921 7788 50952
rect 9582 50940 9588 50992
rect 9640 50940 9646 50992
rect 7745 50915 7803 50921
rect 7745 50881 7757 50915
rect 7791 50881 7803 50915
rect 7745 50875 7803 50881
rect 7834 50872 7840 50924
rect 7892 50912 7898 50924
rect 9401 50915 9459 50921
rect 9401 50912 9413 50915
rect 7892 50884 9413 50912
rect 7892 50872 7898 50884
rect 9401 50881 9413 50884
rect 9447 50881 9459 50915
rect 9401 50875 9459 50881
rect 24765 50915 24823 50921
rect 24765 50881 24777 50915
rect 24811 50912 24823 50915
rect 25038 50912 25044 50924
rect 24811 50884 25044 50912
rect 24811 50881 24823 50884
rect 24765 50875 24823 50881
rect 25038 50872 25044 50884
rect 25096 50872 25102 50924
rect 4338 50804 4344 50856
rect 4396 50844 4402 50856
rect 4617 50847 4675 50853
rect 4617 50844 4629 50847
rect 4396 50816 4629 50844
rect 4396 50804 4402 50816
rect 4617 50813 4629 50816
rect 4663 50813 4675 50847
rect 4617 50807 4675 50813
rect 7466 50804 7472 50856
rect 7524 50804 7530 50856
rect 4154 50776 4160 50788
rect 2884 50748 4160 50776
rect 4154 50736 4160 50748
rect 4212 50736 4218 50788
rect 25225 50711 25283 50717
rect 25225 50677 25237 50711
rect 25271 50708 25283 50711
rect 25682 50708 25688 50720
rect 25271 50680 25688 50708
rect 25271 50677 25283 50680
rect 25225 50671 25283 50677
rect 25682 50668 25688 50680
rect 25740 50668 25746 50720
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 6822 50464 6828 50516
rect 6880 50464 6886 50516
rect 8662 50464 8668 50516
rect 8720 50504 8726 50516
rect 9217 50507 9275 50513
rect 9217 50504 9229 50507
rect 8720 50476 9229 50504
rect 8720 50464 8726 50476
rect 9217 50473 9229 50476
rect 9263 50473 9275 50507
rect 9217 50467 9275 50473
rect 2746 50408 4016 50436
rect 1302 50328 1308 50380
rect 1360 50368 1366 50380
rect 2746 50368 2774 50408
rect 1360 50340 2774 50368
rect 3237 50371 3295 50377
rect 1360 50328 1366 50340
rect 3237 50337 3249 50371
rect 3283 50368 3295 50371
rect 3418 50368 3424 50380
rect 3283 50340 3424 50368
rect 3283 50337 3295 50340
rect 3237 50331 3295 50337
rect 3418 50328 3424 50340
rect 3476 50328 3482 50380
rect 3988 50377 4016 50408
rect 3973 50371 4031 50377
rect 3973 50337 3985 50371
rect 4019 50368 4031 50371
rect 5077 50371 5135 50377
rect 5077 50368 5089 50371
rect 4019 50340 5089 50368
rect 4019 50337 4031 50340
rect 3973 50331 4031 50337
rect 5077 50337 5089 50340
rect 5123 50337 5135 50371
rect 5077 50331 5135 50337
rect 2225 50303 2283 50309
rect 2225 50269 2237 50303
rect 2271 50269 2283 50303
rect 2225 50263 2283 50269
rect 4249 50303 4307 50309
rect 4249 50269 4261 50303
rect 4295 50300 4307 50303
rect 4430 50300 4436 50312
rect 4295 50272 4436 50300
rect 4295 50269 4307 50272
rect 4249 50263 4307 50269
rect 2240 50232 2268 50263
rect 4430 50260 4436 50272
rect 4488 50260 4494 50312
rect 5810 50260 5816 50312
rect 5868 50300 5874 50312
rect 7009 50303 7067 50309
rect 7009 50300 7021 50303
rect 5868 50272 7021 50300
rect 5868 50260 5874 50272
rect 7009 50269 7021 50272
rect 7055 50269 7067 50303
rect 7009 50263 7067 50269
rect 9398 50260 9404 50312
rect 9456 50260 9462 50312
rect 5074 50232 5080 50244
rect 2240 50204 5080 50232
rect 5074 50192 5080 50204
rect 5132 50192 5138 50244
rect 25314 50124 25320 50176
rect 25372 50164 25378 50176
rect 25409 50167 25467 50173
rect 25409 50164 25421 50167
rect 25372 50136 25421 50164
rect 25372 50124 25378 50136
rect 25409 50133 25421 50136
rect 25455 50133 25467 50167
rect 25409 50127 25467 50133
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 6549 49963 6607 49969
rect 6549 49960 6561 49963
rect 3988 49932 6561 49960
rect 3145 49895 3203 49901
rect 3145 49861 3157 49895
rect 3191 49892 3203 49895
rect 3510 49892 3516 49904
rect 3191 49864 3516 49892
rect 3191 49861 3203 49864
rect 3145 49855 3203 49861
rect 3510 49852 3516 49864
rect 3568 49852 3574 49904
rect 1946 49784 1952 49836
rect 2004 49784 2010 49836
rect 3988 49833 4016 49932
rect 6549 49929 6561 49932
rect 6595 49960 6607 49963
rect 9858 49960 9864 49972
rect 6595 49932 9864 49960
rect 6595 49929 6607 49932
rect 6549 49923 6607 49929
rect 9858 49920 9864 49932
rect 9916 49920 9922 49972
rect 20990 49920 20996 49972
rect 21048 49960 21054 49972
rect 25133 49963 25191 49969
rect 25133 49960 25145 49963
rect 21048 49932 25145 49960
rect 21048 49920 21054 49932
rect 25133 49929 25145 49932
rect 25179 49929 25191 49963
rect 25133 49923 25191 49929
rect 4246 49852 4252 49904
rect 4304 49852 4310 49904
rect 6365 49895 6423 49901
rect 6365 49892 6377 49895
rect 5474 49864 6377 49892
rect 6365 49861 6377 49864
rect 6411 49892 6423 49895
rect 9030 49892 9036 49904
rect 6411 49864 9036 49892
rect 6411 49861 6423 49864
rect 6365 49855 6423 49861
rect 9030 49852 9036 49864
rect 9088 49852 9094 49904
rect 9306 49852 9312 49904
rect 9364 49852 9370 49904
rect 3973 49827 4031 49833
rect 3973 49793 3985 49827
rect 4019 49793 4031 49827
rect 3973 49787 4031 49793
rect 7742 49784 7748 49836
rect 7800 49824 7806 49836
rect 9125 49827 9183 49833
rect 9125 49824 9137 49827
rect 7800 49796 9137 49824
rect 7800 49784 7806 49796
rect 9125 49793 9137 49796
rect 9171 49793 9183 49827
rect 9125 49787 9183 49793
rect 25314 49784 25320 49836
rect 25372 49784 25378 49836
rect 5997 49759 6055 49765
rect 5997 49725 6009 49759
rect 6043 49756 6055 49759
rect 8846 49756 8852 49768
rect 6043 49728 8852 49756
rect 6043 49725 6055 49728
rect 5997 49719 6055 49725
rect 8846 49716 8852 49728
rect 8904 49716 8910 49768
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 11609 49419 11667 49425
rect 11609 49385 11621 49419
rect 11655 49416 11667 49419
rect 11974 49416 11980 49428
rect 11655 49388 11980 49416
rect 11655 49385 11667 49388
rect 11609 49379 11667 49385
rect 11974 49376 11980 49388
rect 12032 49376 12038 49428
rect 1486 49240 1492 49292
rect 1544 49280 1550 49292
rect 2041 49283 2099 49289
rect 2041 49280 2053 49283
rect 1544 49252 2053 49280
rect 1544 49240 1550 49252
rect 2041 49249 2053 49252
rect 2087 49249 2099 49283
rect 2041 49243 2099 49249
rect 1765 49215 1823 49221
rect 1765 49181 1777 49215
rect 1811 49212 1823 49215
rect 1811 49184 2774 49212
rect 1811 49181 1823 49184
rect 1765 49175 1823 49181
rect 2746 49076 2774 49184
rect 10686 49172 10692 49224
rect 10744 49212 10750 49224
rect 11793 49215 11851 49221
rect 11793 49212 11805 49215
rect 10744 49184 11805 49212
rect 10744 49172 10750 49184
rect 11793 49181 11805 49184
rect 11839 49181 11851 49215
rect 11793 49175 11851 49181
rect 24857 49215 24915 49221
rect 24857 49181 24869 49215
rect 24903 49212 24915 49215
rect 25314 49212 25320 49224
rect 24903 49184 25320 49212
rect 24903 49181 24915 49184
rect 24857 49175 24915 49181
rect 25314 49172 25320 49184
rect 25372 49172 25378 49224
rect 3329 49079 3387 49085
rect 3329 49076 3341 49079
rect 2746 49048 3341 49076
rect 3329 49045 3341 49048
rect 3375 49076 3387 49079
rect 10778 49076 10784 49088
rect 3375 49048 10784 49076
rect 3375 49045 3387 49048
rect 3329 49039 3387 49045
rect 10778 49036 10784 49048
rect 10836 49036 10842 49088
rect 18322 49036 18328 49088
rect 18380 49076 18386 49088
rect 25133 49079 25191 49085
rect 25133 49076 25145 49079
rect 18380 49048 25145 49076
rect 18380 49036 18386 49048
rect 25133 49045 25145 49048
rect 25179 49045 25191 49079
rect 25133 49039 25191 49045
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 12713 48875 12771 48881
rect 12713 48841 12725 48875
rect 12759 48872 12771 48875
rect 12802 48872 12808 48884
rect 12759 48844 12808 48872
rect 12759 48841 12771 48844
rect 12713 48835 12771 48841
rect 12802 48832 12808 48844
rect 12860 48832 12866 48884
rect 12526 48696 12532 48748
rect 12584 48736 12590 48748
rect 12897 48739 12955 48745
rect 12897 48736 12909 48739
rect 12584 48708 12909 48736
rect 12584 48696 12590 48708
rect 12897 48705 12909 48708
rect 12943 48705 12955 48739
rect 12897 48699 12955 48705
rect 25498 48492 25504 48544
rect 25556 48492 25562 48544
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 17310 48220 17316 48272
rect 17368 48260 17374 48272
rect 17773 48263 17831 48269
rect 17773 48260 17785 48263
rect 17368 48232 17785 48260
rect 17368 48220 17374 48232
rect 17773 48229 17785 48232
rect 17819 48260 17831 48263
rect 19426 48260 19432 48272
rect 17819 48232 19432 48260
rect 17819 48229 17831 48232
rect 17773 48223 17831 48229
rect 19426 48220 19432 48232
rect 19484 48220 19490 48272
rect 24857 48127 24915 48133
rect 24857 48093 24869 48127
rect 24903 48124 24915 48127
rect 25314 48124 25320 48136
rect 24903 48096 25320 48124
rect 24903 48093 24915 48096
rect 24857 48087 24915 48093
rect 25314 48084 25320 48096
rect 25372 48084 25378 48136
rect 1302 48016 1308 48068
rect 1360 48056 1366 48068
rect 1673 48059 1731 48065
rect 1673 48056 1685 48059
rect 1360 48028 1685 48056
rect 1360 48016 1366 48028
rect 1673 48025 1685 48028
rect 1719 48056 1731 48059
rect 2133 48059 2191 48065
rect 2133 48056 2145 48059
rect 1719 48028 2145 48056
rect 1719 48025 1731 48028
rect 1673 48019 1731 48025
rect 2133 48025 2145 48028
rect 2179 48025 2191 48059
rect 2133 48019 2191 48025
rect 1765 47991 1823 47997
rect 1765 47957 1777 47991
rect 1811 47988 1823 47991
rect 4062 47988 4068 48000
rect 1811 47960 4068 47988
rect 1811 47957 1823 47960
rect 1765 47951 1823 47957
rect 4062 47948 4068 47960
rect 4120 47948 4126 48000
rect 7558 47948 7564 48000
rect 7616 47988 7622 48000
rect 11330 47988 11336 48000
rect 7616 47960 11336 47988
rect 7616 47948 7622 47960
rect 11330 47948 11336 47960
rect 11388 47948 11394 48000
rect 20254 47948 20260 48000
rect 20312 47988 20318 48000
rect 25133 47991 25191 47997
rect 25133 47988 25145 47991
rect 20312 47960 25145 47988
rect 20312 47948 20318 47960
rect 25133 47957 25145 47960
rect 25179 47957 25191 47991
rect 25133 47951 25191 47957
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 9122 47744 9128 47796
rect 9180 47744 9186 47796
rect 17218 47744 17224 47796
rect 17276 47744 17282 47796
rect 17310 47744 17316 47796
rect 17368 47744 17374 47796
rect 18414 47744 18420 47796
rect 18472 47744 18478 47796
rect 18506 47744 18512 47796
rect 18564 47784 18570 47796
rect 19061 47787 19119 47793
rect 19061 47784 19073 47787
rect 18564 47756 19073 47784
rect 18564 47744 18570 47756
rect 19061 47753 19073 47756
rect 19107 47753 19119 47787
rect 19061 47747 19119 47753
rect 9309 47651 9367 47657
rect 9309 47617 9321 47651
rect 9355 47648 9367 47651
rect 11422 47648 11428 47660
rect 9355 47620 11428 47648
rect 9355 47617 9367 47620
rect 9309 47611 9367 47617
rect 11422 47608 11428 47620
rect 11480 47608 11486 47660
rect 24394 47608 24400 47660
rect 24452 47648 24458 47660
rect 24765 47651 24823 47657
rect 24765 47648 24777 47651
rect 24452 47620 24777 47648
rect 24452 47608 24458 47620
rect 24765 47617 24777 47620
rect 24811 47617 24823 47651
rect 24765 47611 24823 47617
rect 17405 47583 17463 47589
rect 17405 47549 17417 47583
rect 17451 47549 17463 47583
rect 17405 47543 17463 47549
rect 16298 47472 16304 47524
rect 16356 47512 16362 47524
rect 17420 47512 17448 47543
rect 18414 47540 18420 47592
rect 18472 47580 18478 47592
rect 18601 47583 18659 47589
rect 18601 47580 18613 47583
rect 18472 47552 18613 47580
rect 18472 47540 18478 47552
rect 18601 47549 18613 47552
rect 18647 47549 18659 47583
rect 18601 47543 18659 47549
rect 24489 47583 24547 47589
rect 24489 47549 24501 47583
rect 24535 47580 24547 47583
rect 25498 47580 25504 47592
rect 24535 47552 25504 47580
rect 24535 47549 24547 47552
rect 24489 47543 24547 47549
rect 25498 47540 25504 47552
rect 25556 47540 25562 47592
rect 16356 47484 17448 47512
rect 16356 47472 16362 47484
rect 16574 47404 16580 47456
rect 16632 47444 16638 47456
rect 16853 47447 16911 47453
rect 16853 47444 16865 47447
rect 16632 47416 16865 47444
rect 16632 47404 16638 47416
rect 16853 47413 16865 47416
rect 16899 47413 16911 47447
rect 16853 47407 16911 47413
rect 17494 47404 17500 47456
rect 17552 47444 17558 47456
rect 18049 47447 18107 47453
rect 18049 47444 18061 47447
rect 17552 47416 18061 47444
rect 17552 47404 17558 47416
rect 18049 47413 18061 47416
rect 18095 47413 18107 47447
rect 18049 47407 18107 47413
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 9858 47200 9864 47252
rect 9916 47200 9922 47252
rect 15920 47243 15978 47249
rect 15920 47209 15932 47243
rect 15966 47240 15978 47243
rect 18414 47240 18420 47252
rect 15966 47212 18420 47240
rect 15966 47209 15978 47212
rect 15920 47203 15978 47209
rect 18414 47200 18420 47212
rect 18472 47200 18478 47252
rect 19337 47243 19395 47249
rect 19337 47209 19349 47243
rect 19383 47240 19395 47243
rect 20346 47240 20352 47252
rect 19383 47212 20352 47240
rect 19383 47209 19395 47212
rect 19337 47203 19395 47209
rect 9876 47104 9904 47200
rect 18141 47175 18199 47181
rect 18141 47141 18153 47175
rect 18187 47172 18199 47175
rect 18506 47172 18512 47184
rect 18187 47144 18512 47172
rect 18187 47141 18199 47144
rect 18141 47135 18199 47141
rect 18506 47132 18512 47144
rect 18564 47132 18570 47184
rect 19352 47172 19380 47203
rect 20346 47200 20352 47212
rect 20404 47200 20410 47252
rect 21634 47200 21640 47252
rect 21692 47200 21698 47252
rect 18708 47144 19380 47172
rect 10229 47107 10287 47113
rect 10229 47104 10241 47107
rect 9876 47076 10241 47104
rect 10229 47073 10241 47076
rect 10275 47073 10287 47107
rect 10229 47067 10287 47073
rect 15657 47107 15715 47113
rect 15657 47073 15669 47107
rect 15703 47104 15715 47107
rect 16666 47104 16672 47116
rect 15703 47076 16672 47104
rect 15703 47073 15715 47076
rect 15657 47067 15715 47073
rect 16666 47064 16672 47076
rect 16724 47064 16730 47116
rect 16942 47064 16948 47116
rect 17000 47104 17006 47116
rect 17000 47076 17172 47104
rect 17000 47064 17006 47076
rect 17144 47036 17172 47076
rect 17310 47064 17316 47116
rect 17368 47104 17374 47116
rect 17405 47107 17463 47113
rect 17405 47104 17417 47107
rect 17368 47076 17417 47104
rect 17368 47064 17374 47076
rect 17405 47073 17417 47076
rect 17451 47073 17463 47107
rect 17405 47067 17463 47073
rect 18598 47064 18604 47116
rect 18656 47064 18662 47116
rect 18509 47039 18567 47045
rect 18509 47036 18521 47039
rect 17144 47008 18521 47036
rect 18509 47005 18521 47008
rect 18555 47036 18567 47039
rect 18708 47036 18736 47144
rect 21818 47132 21824 47184
rect 21876 47172 21882 47184
rect 25133 47175 25191 47181
rect 25133 47172 25145 47175
rect 21876 47144 25145 47172
rect 21876 47132 21882 47144
rect 25133 47141 25145 47144
rect 25179 47141 25191 47175
rect 25133 47135 25191 47141
rect 18785 47107 18843 47113
rect 18785 47073 18797 47107
rect 18831 47104 18843 47107
rect 19334 47104 19340 47116
rect 18831 47076 19340 47104
rect 18831 47073 18843 47076
rect 18785 47067 18843 47073
rect 19334 47064 19340 47076
rect 19392 47064 19398 47116
rect 22557 47107 22615 47113
rect 22557 47073 22569 47107
rect 22603 47104 22615 47107
rect 22603 47076 22784 47104
rect 22603 47073 22615 47076
rect 22557 47067 22615 47073
rect 18555 47008 18736 47036
rect 18555 47005 18567 47008
rect 18509 46999 18567 47005
rect 21634 46996 21640 47048
rect 21692 47036 21698 47048
rect 22373 47039 22431 47045
rect 22373 47036 22385 47039
rect 21692 47008 22385 47036
rect 21692 46996 21698 47008
rect 22373 47005 22385 47008
rect 22419 47005 22431 47039
rect 22373 46999 22431 47005
rect 22465 47039 22523 47045
rect 22465 47005 22477 47039
rect 22511 47036 22523 47039
rect 22646 47036 22652 47048
rect 22511 47008 22652 47036
rect 22511 47005 22523 47008
rect 22465 46999 22523 47005
rect 22646 46996 22652 47008
rect 22704 46996 22710 47048
rect 9030 46928 9036 46980
rect 9088 46968 9094 46980
rect 9088 46940 9674 46968
rect 9088 46928 9094 46940
rect 9646 46900 9674 46940
rect 10502 46928 10508 46980
rect 10560 46928 10566 46980
rect 12253 46971 12311 46977
rect 12253 46968 12265 46971
rect 10888 46940 10994 46968
rect 11900 46940 12265 46968
rect 10042 46900 10048 46912
rect 9646 46872 10048 46900
rect 10042 46860 10048 46872
rect 10100 46900 10106 46912
rect 10888 46900 10916 46940
rect 11900 46900 11928 46940
rect 12253 46937 12265 46940
rect 12299 46968 12311 46971
rect 12618 46968 12624 46980
rect 12299 46940 12624 46968
rect 12299 46937 12311 46940
rect 12253 46931 12311 46937
rect 12618 46928 12624 46940
rect 12676 46968 12682 46980
rect 13078 46968 13084 46980
rect 12676 46940 13084 46968
rect 12676 46928 12682 46940
rect 13078 46928 13084 46940
rect 13136 46968 13142 46980
rect 14185 46971 14243 46977
rect 14185 46968 14197 46971
rect 13136 46940 14197 46968
rect 13136 46928 13142 46940
rect 14185 46937 14197 46940
rect 14231 46937 14243 46971
rect 14185 46931 14243 46937
rect 16390 46928 16396 46980
rect 16448 46928 16454 46980
rect 10100 46872 11928 46900
rect 11977 46903 12035 46909
rect 10100 46860 10106 46872
rect 11977 46869 11989 46903
rect 12023 46900 12035 46903
rect 12158 46900 12164 46912
rect 12023 46872 12164 46900
rect 12023 46869 12035 46872
rect 11977 46863 12035 46869
rect 12158 46860 12164 46872
rect 12216 46860 12222 46912
rect 17586 46860 17592 46912
rect 17644 46900 17650 46912
rect 17681 46903 17739 46909
rect 17681 46900 17693 46903
rect 17644 46872 17693 46900
rect 17644 46860 17650 46872
rect 17681 46869 17693 46872
rect 17727 46869 17739 46903
rect 17681 46863 17739 46869
rect 22002 46860 22008 46912
rect 22060 46860 22066 46912
rect 22646 46860 22652 46912
rect 22704 46900 22710 46912
rect 22756 46900 22784 47076
rect 25317 47039 25375 47045
rect 25317 47036 25329 47039
rect 24872 47008 25329 47036
rect 24762 46928 24768 46980
rect 24820 46968 24826 46980
rect 24872 46977 24900 47008
rect 25317 47005 25329 47008
rect 25363 47005 25375 47039
rect 25317 46999 25375 47005
rect 24857 46971 24915 46977
rect 24857 46968 24869 46971
rect 24820 46940 24869 46968
rect 24820 46928 24826 46940
rect 24857 46937 24869 46940
rect 24903 46937 24915 46971
rect 24857 46931 24915 46937
rect 22704 46872 22784 46900
rect 22704 46860 22710 46872
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 7193 46699 7251 46705
rect 7193 46665 7205 46699
rect 7239 46696 7251 46699
rect 7466 46696 7472 46708
rect 7239 46668 7472 46696
rect 7239 46665 7251 46668
rect 7193 46659 7251 46665
rect 7466 46656 7472 46668
rect 7524 46656 7530 46708
rect 10870 46656 10876 46708
rect 10928 46656 10934 46708
rect 14182 46696 14188 46708
rect 12636 46668 14188 46696
rect 12636 46637 12664 46668
rect 14182 46656 14188 46668
rect 14240 46656 14246 46708
rect 18414 46656 18420 46708
rect 18472 46696 18478 46708
rect 18601 46699 18659 46705
rect 18601 46696 18613 46699
rect 18472 46668 18613 46696
rect 18472 46656 18478 46668
rect 18601 46665 18613 46668
rect 18647 46665 18659 46699
rect 18601 46659 18659 46665
rect 18966 46656 18972 46708
rect 19024 46696 19030 46708
rect 20809 46699 20867 46705
rect 20809 46696 20821 46699
rect 19024 46668 20821 46696
rect 19024 46656 19030 46668
rect 20809 46665 20821 46668
rect 20855 46665 20867 46699
rect 20809 46659 20867 46665
rect 22554 46656 22560 46708
rect 22612 46696 22618 46708
rect 22649 46699 22707 46705
rect 22649 46696 22661 46699
rect 22612 46668 22661 46696
rect 22612 46656 22618 46668
rect 22649 46665 22661 46668
rect 22695 46665 22707 46699
rect 22649 46659 22707 46665
rect 12621 46631 12679 46637
rect 12621 46597 12633 46631
rect 12667 46597 12679 46631
rect 12621 46591 12679 46597
rect 13078 46588 13084 46640
rect 13136 46588 13142 46640
rect 15102 46588 15108 46640
rect 15160 46628 15166 46640
rect 15160 46600 15318 46628
rect 15160 46588 15166 46600
rect 16390 46588 16396 46640
rect 16448 46628 16454 46640
rect 17586 46628 17592 46640
rect 16448 46600 17592 46628
rect 16448 46588 16454 46600
rect 17586 46588 17592 46600
rect 17644 46588 17650 46640
rect 20898 46628 20904 46640
rect 20562 46600 20904 46628
rect 20898 46588 20904 46600
rect 20956 46628 20962 46640
rect 21085 46631 21143 46637
rect 21085 46628 21097 46631
rect 20956 46600 21097 46628
rect 20956 46588 20962 46600
rect 21085 46597 21097 46600
rect 21131 46597 21143 46631
rect 22664 46628 22692 46659
rect 22738 46656 22744 46708
rect 22796 46656 22802 46708
rect 23477 46631 23535 46637
rect 23477 46628 23489 46631
rect 22664 46600 23489 46628
rect 21085 46591 21143 46597
rect 23477 46597 23489 46600
rect 23523 46597 23535 46631
rect 23477 46591 23535 46597
rect 7377 46563 7435 46569
rect 7377 46529 7389 46563
rect 7423 46560 7435 46563
rect 7558 46560 7564 46572
rect 7423 46532 7564 46560
rect 7423 46529 7435 46532
rect 7377 46523 7435 46529
rect 7558 46520 7564 46532
rect 7616 46520 7622 46572
rect 11054 46520 11060 46572
rect 11112 46520 11118 46572
rect 24210 46520 24216 46572
rect 24268 46560 24274 46572
rect 24765 46563 24823 46569
rect 24765 46560 24777 46563
rect 24268 46532 24777 46560
rect 24268 46520 24274 46532
rect 24765 46529 24777 46532
rect 24811 46529 24823 46563
rect 24765 46523 24823 46529
rect 11882 46452 11888 46504
rect 11940 46492 11946 46504
rect 12345 46495 12403 46501
rect 12345 46492 12357 46495
rect 11940 46464 12357 46492
rect 11940 46452 11946 46464
rect 12345 46461 12357 46464
rect 12391 46492 12403 46495
rect 13354 46492 13360 46504
rect 12391 46464 13360 46492
rect 12391 46461 12403 46464
rect 12345 46455 12403 46461
rect 13354 46452 13360 46464
rect 13412 46492 13418 46504
rect 14553 46495 14611 46501
rect 14553 46492 14565 46495
rect 13412 46464 14565 46492
rect 13412 46452 13418 46464
rect 14553 46461 14565 46464
rect 14599 46461 14611 46495
rect 14553 46455 14611 46461
rect 14829 46495 14887 46501
rect 14829 46461 14841 46495
rect 14875 46492 14887 46495
rect 14875 46464 16574 46492
rect 14875 46461 14887 46464
rect 14829 46455 14887 46461
rect 13722 46316 13728 46368
rect 13780 46356 13786 46368
rect 14093 46359 14151 46365
rect 14093 46356 14105 46359
rect 13780 46328 14105 46356
rect 13780 46316 13786 46328
rect 14093 46325 14105 46328
rect 14139 46325 14151 46359
rect 14093 46319 14151 46325
rect 16298 46316 16304 46368
rect 16356 46316 16362 46368
rect 16546 46356 16574 46464
rect 16850 46452 16856 46504
rect 16908 46452 16914 46504
rect 17129 46495 17187 46501
rect 17129 46461 17141 46495
rect 17175 46492 17187 46495
rect 18598 46492 18604 46504
rect 17175 46464 18604 46492
rect 17175 46461 17187 46464
rect 17129 46455 17187 46461
rect 18598 46452 18604 46464
rect 18656 46452 18662 46504
rect 19061 46495 19119 46501
rect 19061 46461 19073 46495
rect 19107 46461 19119 46495
rect 19061 46455 19119 46461
rect 17218 46356 17224 46368
rect 16546 46328 17224 46356
rect 17218 46316 17224 46328
rect 17276 46316 17282 46368
rect 19076 46356 19104 46455
rect 19334 46452 19340 46504
rect 19392 46452 19398 46504
rect 22186 46452 22192 46504
rect 22244 46492 22250 46504
rect 22833 46495 22891 46501
rect 22833 46492 22845 46495
rect 22244 46464 22845 46492
rect 22244 46452 22250 46464
rect 22833 46461 22845 46464
rect 22879 46492 22891 46495
rect 23293 46495 23351 46501
rect 23293 46492 23305 46495
rect 22879 46464 23305 46492
rect 22879 46461 22891 46464
rect 22833 46455 22891 46461
rect 23293 46461 23305 46464
rect 23339 46461 23351 46495
rect 23293 46455 23351 46461
rect 24486 46452 24492 46504
rect 24544 46452 24550 46504
rect 19426 46356 19432 46368
rect 19076 46328 19432 46356
rect 19426 46316 19432 46328
rect 19484 46316 19490 46368
rect 22281 46359 22339 46365
rect 22281 46325 22293 46359
rect 22327 46356 22339 46359
rect 22738 46356 22744 46368
rect 22327 46328 22744 46356
rect 22327 46325 22339 46328
rect 22281 46319 22339 46325
rect 22738 46316 22744 46328
rect 22796 46316 22802 46368
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 5902 46112 5908 46164
rect 5960 46152 5966 46164
rect 8113 46155 8171 46161
rect 8113 46152 8125 46155
rect 5960 46124 8125 46152
rect 5960 46112 5966 46124
rect 8113 46121 8125 46124
rect 8159 46121 8171 46155
rect 8113 46115 8171 46121
rect 9125 46155 9183 46161
rect 9125 46121 9137 46155
rect 9171 46152 9183 46155
rect 9214 46152 9220 46164
rect 9171 46124 9220 46152
rect 9171 46121 9183 46124
rect 9125 46115 9183 46121
rect 9214 46112 9220 46124
rect 9272 46112 9278 46164
rect 10686 46112 10692 46164
rect 10744 46112 10750 46164
rect 17586 46112 17592 46164
rect 17644 46152 17650 46164
rect 18693 46155 18751 46161
rect 18693 46152 18705 46155
rect 17644 46124 18705 46152
rect 17644 46112 17650 46124
rect 18693 46121 18705 46124
rect 18739 46121 18751 46155
rect 18693 46115 18751 46121
rect 19429 46155 19487 46161
rect 19429 46121 19441 46155
rect 19475 46152 19487 46155
rect 19610 46152 19616 46164
rect 19475 46124 19616 46152
rect 19475 46121 19487 46124
rect 19429 46115 19487 46121
rect 19610 46112 19616 46124
rect 19668 46112 19674 46164
rect 24486 46112 24492 46164
rect 24544 46152 24550 46164
rect 25409 46155 25467 46161
rect 25409 46152 25421 46155
rect 24544 46124 25421 46152
rect 24544 46112 24550 46124
rect 25409 46121 25421 46124
rect 25455 46152 25467 46155
rect 25498 46152 25504 46164
rect 25455 46124 25504 46152
rect 25455 46121 25467 46124
rect 25409 46115 25467 46121
rect 25498 46112 25504 46124
rect 25556 46112 25562 46164
rect 7650 46044 7656 46096
rect 7708 46084 7714 46096
rect 10045 46087 10103 46093
rect 10045 46084 10057 46087
rect 7708 46056 10057 46084
rect 7708 46044 7714 46056
rect 10045 46053 10057 46056
rect 10091 46053 10103 46087
rect 10045 46047 10103 46053
rect 11348 46056 12020 46084
rect 1857 46019 1915 46025
rect 1857 45985 1869 46019
rect 1903 46016 1915 46019
rect 9490 46016 9496 46028
rect 1903 45988 9496 46016
rect 1903 45985 1915 45988
rect 1857 45979 1915 45985
rect 9490 45976 9496 45988
rect 9548 45976 9554 46028
rect 11348 46025 11376 46056
rect 11333 46019 11391 46025
rect 11333 45985 11345 46019
rect 11379 45985 11391 46019
rect 11333 45979 11391 45985
rect 11882 45976 11888 46028
rect 11940 45976 11946 46028
rect 11992 46016 12020 46056
rect 12158 46016 12164 46028
rect 11992 45988 12164 46016
rect 12158 45976 12164 45988
rect 12216 45976 12222 46028
rect 12618 45976 12624 46028
rect 12676 46016 12682 46028
rect 13998 46016 14004 46028
rect 12676 45988 14004 46016
rect 12676 45976 12682 45988
rect 13998 45976 14004 45988
rect 14056 46016 14062 46028
rect 14093 46019 14151 46025
rect 14093 46016 14105 46019
rect 14056 45988 14105 46016
rect 14056 45976 14062 45988
rect 14093 45985 14105 45988
rect 14139 45985 14151 46019
rect 14093 45979 14151 45985
rect 20162 45976 20168 46028
rect 20220 45976 20226 46028
rect 20349 46019 20407 46025
rect 20349 45985 20361 46019
rect 20395 46016 20407 46019
rect 20438 46016 20444 46028
rect 20395 45988 20444 46016
rect 20395 45985 20407 45988
rect 20349 45979 20407 45985
rect 20438 45976 20444 45988
rect 20496 45976 20502 46028
rect 21358 45976 21364 46028
rect 21416 45976 21422 46028
rect 21545 46019 21603 46025
rect 21545 45985 21557 46019
rect 21591 46016 21603 46019
rect 21726 46016 21732 46028
rect 21591 45988 21732 46016
rect 21591 45985 21603 45988
rect 21545 45979 21603 45985
rect 21726 45976 21732 45988
rect 21784 45976 21790 46028
rect 1302 45908 1308 45960
rect 1360 45948 1366 45960
rect 1581 45951 1639 45957
rect 1581 45948 1593 45951
rect 1360 45920 1593 45948
rect 1360 45908 1366 45920
rect 1581 45917 1593 45920
rect 1627 45917 1639 45951
rect 1581 45911 1639 45917
rect 7190 45908 7196 45960
rect 7248 45948 7254 45960
rect 9309 45951 9367 45957
rect 9309 45948 9321 45951
rect 7248 45920 9321 45948
rect 7248 45908 7254 45920
rect 9309 45917 9321 45920
rect 9355 45917 9367 45951
rect 9309 45911 9367 45917
rect 10229 45951 10287 45957
rect 10229 45917 10241 45951
rect 10275 45917 10287 45951
rect 10229 45911 10287 45917
rect 11057 45951 11115 45957
rect 11057 45917 11069 45951
rect 11103 45948 11115 45951
rect 11790 45948 11796 45960
rect 11103 45920 11796 45948
rect 11103 45917 11115 45920
rect 11057 45911 11115 45917
rect 6914 45840 6920 45892
rect 6972 45880 6978 45892
rect 8021 45883 8079 45889
rect 8021 45880 8033 45883
rect 6972 45852 8033 45880
rect 6972 45840 6978 45852
rect 8021 45849 8033 45852
rect 8067 45880 8079 45883
rect 8481 45883 8539 45889
rect 8481 45880 8493 45883
rect 8067 45852 8493 45880
rect 8067 45849 8079 45852
rect 8021 45843 8079 45849
rect 8481 45849 8493 45852
rect 8527 45849 8539 45883
rect 10244 45880 10272 45911
rect 11790 45908 11796 45920
rect 11848 45908 11854 45960
rect 19610 45908 19616 45960
rect 19668 45948 19674 45960
rect 20070 45948 20076 45960
rect 19668 45920 20076 45948
rect 19668 45908 19674 45920
rect 20070 45908 20076 45920
rect 20128 45908 20134 45960
rect 21082 45908 21088 45960
rect 21140 45948 21146 45960
rect 21269 45951 21327 45957
rect 21269 45948 21281 45951
rect 21140 45920 21281 45948
rect 21140 45908 21146 45920
rect 21269 45917 21281 45920
rect 21315 45948 21327 45951
rect 21910 45948 21916 45960
rect 21315 45920 21916 45948
rect 21315 45917 21327 45920
rect 21269 45911 21327 45917
rect 21910 45908 21916 45920
rect 21968 45908 21974 45960
rect 23201 45951 23259 45957
rect 23201 45917 23213 45951
rect 23247 45917 23259 45951
rect 23201 45911 23259 45917
rect 23477 45951 23535 45957
rect 23477 45917 23489 45951
rect 23523 45948 23535 45951
rect 24026 45948 24032 45960
rect 23523 45920 24032 45948
rect 23523 45917 23535 45920
rect 23477 45911 23535 45917
rect 10244 45852 12434 45880
rect 8481 45843 8539 45849
rect 11146 45772 11152 45824
rect 11204 45772 11210 45824
rect 12406 45812 12434 45852
rect 12618 45840 12624 45892
rect 12676 45840 12682 45892
rect 14734 45880 14740 45892
rect 13556 45852 14740 45880
rect 13556 45812 13584 45852
rect 14734 45840 14740 45852
rect 14792 45840 14798 45892
rect 12406 45784 13584 45812
rect 13630 45772 13636 45824
rect 13688 45772 13694 45824
rect 16390 45772 16396 45824
rect 16448 45772 16454 45824
rect 19705 45815 19763 45821
rect 19705 45781 19717 45815
rect 19751 45812 19763 45815
rect 19886 45812 19892 45824
rect 19751 45784 19892 45812
rect 19751 45781 19763 45784
rect 19705 45775 19763 45781
rect 19886 45772 19892 45784
rect 19944 45772 19950 45824
rect 20714 45772 20720 45824
rect 20772 45812 20778 45824
rect 20901 45815 20959 45821
rect 20901 45812 20913 45815
rect 20772 45784 20913 45812
rect 20772 45772 20778 45784
rect 20901 45781 20913 45784
rect 20947 45781 20959 45815
rect 23216 45812 23244 45911
rect 24026 45908 24032 45920
rect 24084 45908 24090 45960
rect 24489 45815 24547 45821
rect 24489 45812 24501 45815
rect 23216 45784 24501 45812
rect 20901 45775 20959 45781
rect 24489 45781 24501 45784
rect 24535 45812 24547 45815
rect 24854 45812 24860 45824
rect 24535 45784 24860 45812
rect 24535 45781 24547 45784
rect 24489 45775 24547 45781
rect 24854 45772 24860 45784
rect 24912 45772 24918 45824
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 1302 45568 1308 45620
rect 1360 45608 1366 45620
rect 1397 45611 1455 45617
rect 1397 45608 1409 45611
rect 1360 45580 1409 45608
rect 1360 45568 1366 45580
rect 1397 45577 1409 45580
rect 1443 45577 1455 45611
rect 1397 45571 1455 45577
rect 19334 45568 19340 45620
rect 19392 45608 19398 45620
rect 20165 45611 20223 45617
rect 20165 45608 20177 45611
rect 19392 45580 20177 45608
rect 19392 45568 19398 45580
rect 20165 45577 20177 45580
rect 20211 45577 20223 45611
rect 23753 45611 23811 45617
rect 23753 45608 23765 45611
rect 20165 45571 20223 45577
rect 22664 45580 23765 45608
rect 8846 45500 8852 45552
rect 8904 45500 8910 45552
rect 9766 45540 9772 45552
rect 9232 45512 9772 45540
rect 8864 45404 8892 45500
rect 9232 45484 9260 45512
rect 9766 45500 9772 45512
rect 9824 45500 9830 45552
rect 10042 45500 10048 45552
rect 10100 45500 10106 45552
rect 13998 45500 14004 45552
rect 14056 45540 14062 45552
rect 15102 45540 15108 45552
rect 14056 45512 15108 45540
rect 14056 45500 14062 45512
rect 15102 45500 15108 45512
rect 15160 45500 15166 45552
rect 21726 45500 21732 45552
rect 21784 45540 21790 45552
rect 22664 45540 22692 45580
rect 23753 45577 23765 45580
rect 23799 45577 23811 45611
rect 23753 45571 23811 45577
rect 21784 45512 22692 45540
rect 21784 45500 21790 45512
rect 9214 45432 9220 45484
rect 9272 45432 9278 45484
rect 19826 45444 20576 45472
rect 23414 45444 24164 45472
rect 9493 45407 9551 45413
rect 9493 45404 9505 45407
rect 8864 45376 9505 45404
rect 9493 45373 9505 45376
rect 9539 45373 9551 45407
rect 9493 45367 9551 45373
rect 9858 45364 9864 45416
rect 9916 45404 9922 45416
rect 11517 45407 11575 45413
rect 11517 45404 11529 45407
rect 9916 45376 11529 45404
rect 9916 45364 9922 45376
rect 11517 45373 11529 45376
rect 11563 45373 11575 45407
rect 11517 45367 11575 45373
rect 14369 45407 14427 45413
rect 14369 45373 14381 45407
rect 14415 45373 14427 45407
rect 14369 45367 14427 45373
rect 14645 45407 14703 45413
rect 14645 45373 14657 45407
rect 14691 45404 14703 45407
rect 16298 45404 16304 45416
rect 14691 45376 16304 45404
rect 14691 45373 14703 45376
rect 14645 45367 14703 45373
rect 10502 45296 10508 45348
rect 10560 45336 10566 45348
rect 10965 45339 11023 45345
rect 10965 45336 10977 45339
rect 10560 45308 10977 45336
rect 10560 45296 10566 45308
rect 10965 45305 10977 45308
rect 11011 45336 11023 45339
rect 12250 45336 12256 45348
rect 11011 45308 12256 45336
rect 11011 45305 11023 45308
rect 10965 45299 11023 45305
rect 12250 45296 12256 45308
rect 12308 45296 12314 45348
rect 10042 45228 10048 45280
rect 10100 45268 10106 45280
rect 11241 45271 11299 45277
rect 11241 45268 11253 45271
rect 10100 45240 11253 45268
rect 10100 45228 10106 45240
rect 11241 45237 11253 45240
rect 11287 45237 11299 45271
rect 11241 45231 11299 45237
rect 12161 45271 12219 45277
rect 12161 45237 12173 45271
rect 12207 45268 12219 45271
rect 12434 45268 12440 45280
rect 12207 45240 12440 45268
rect 12207 45237 12219 45240
rect 12161 45231 12219 45237
rect 12434 45228 12440 45240
rect 12492 45228 12498 45280
rect 14384 45268 14412 45367
rect 16298 45364 16304 45376
rect 16356 45364 16362 45416
rect 18322 45364 18328 45416
rect 18380 45404 18386 45416
rect 18417 45407 18475 45413
rect 18417 45404 18429 45407
rect 18380 45376 18429 45404
rect 18380 45364 18386 45376
rect 18417 45373 18429 45376
rect 18463 45373 18475 45407
rect 18417 45367 18475 45373
rect 18693 45407 18751 45413
rect 18693 45373 18705 45407
rect 18739 45404 18751 45407
rect 20070 45404 20076 45416
rect 18739 45376 20076 45404
rect 18739 45373 18751 45376
rect 18693 45367 18751 45373
rect 20070 45364 20076 45376
rect 20128 45364 20134 45416
rect 15838 45296 15844 45348
rect 15896 45336 15902 45348
rect 16390 45336 16396 45348
rect 15896 45308 16396 45336
rect 15896 45296 15902 45308
rect 16390 45296 16396 45308
rect 16448 45296 16454 45348
rect 14826 45268 14832 45280
rect 14384 45240 14832 45268
rect 14826 45228 14832 45240
rect 14884 45228 14890 45280
rect 16114 45228 16120 45280
rect 16172 45228 16178 45280
rect 18874 45228 18880 45280
rect 18932 45268 18938 45280
rect 20548 45277 20576 45444
rect 22005 45407 22063 45413
rect 22005 45373 22017 45407
rect 22051 45373 22063 45407
rect 22005 45367 22063 45373
rect 22281 45407 22339 45413
rect 22281 45373 22293 45407
rect 22327 45404 22339 45407
rect 22327 45376 23428 45404
rect 22327 45373 22339 45376
rect 22281 45367 22339 45373
rect 20533 45271 20591 45277
rect 20533 45268 20545 45271
rect 18932 45240 20545 45268
rect 18932 45228 18938 45240
rect 20533 45237 20545 45240
rect 20579 45268 20591 45271
rect 20898 45268 20904 45280
rect 20579 45240 20904 45268
rect 20579 45237 20591 45240
rect 20533 45231 20591 45237
rect 20898 45228 20904 45240
rect 20956 45228 20962 45280
rect 22020 45268 22048 45367
rect 23400 45348 23428 45376
rect 23382 45296 23388 45348
rect 23440 45296 23446 45348
rect 22278 45268 22284 45280
rect 22020 45240 22284 45268
rect 22278 45228 22284 45240
rect 22336 45228 22342 45280
rect 24136 45277 24164 45444
rect 24486 45364 24492 45416
rect 24544 45364 24550 45416
rect 24670 45364 24676 45416
rect 24728 45404 24734 45416
rect 24765 45407 24823 45413
rect 24765 45404 24777 45407
rect 24728 45376 24777 45404
rect 24728 45364 24734 45376
rect 24765 45373 24777 45376
rect 24811 45373 24823 45407
rect 24765 45367 24823 45373
rect 24121 45271 24179 45277
rect 24121 45237 24133 45271
rect 24167 45268 24179 45271
rect 24302 45268 24308 45280
rect 24167 45240 24308 45268
rect 24167 45237 24179 45240
rect 24121 45231 24179 45237
rect 24302 45228 24308 45240
rect 24360 45228 24366 45280
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 7282 45024 7288 45076
rect 7340 45064 7346 45076
rect 9309 45067 9367 45073
rect 9309 45064 9321 45067
rect 7340 45036 9321 45064
rect 7340 45024 7346 45036
rect 9309 45033 9321 45036
rect 9355 45033 9367 45067
rect 9309 45027 9367 45033
rect 11238 45024 11244 45076
rect 11296 45064 11302 45076
rect 11609 45067 11667 45073
rect 11609 45064 11621 45067
rect 11296 45036 11621 45064
rect 11296 45024 11302 45036
rect 11609 45033 11621 45036
rect 11655 45033 11667 45067
rect 11609 45027 11667 45033
rect 12066 45024 12072 45076
rect 12124 45064 12130 45076
rect 12437 45067 12495 45073
rect 12437 45064 12449 45067
rect 12124 45036 12449 45064
rect 12124 45024 12130 45036
rect 12437 45033 12449 45036
rect 12483 45033 12495 45067
rect 12437 45027 12495 45033
rect 12526 45024 12532 45076
rect 12584 45064 12590 45076
rect 12989 45067 13047 45073
rect 12989 45064 13001 45067
rect 12584 45036 13001 45064
rect 12584 45024 12590 45036
rect 12989 45033 13001 45036
rect 13035 45033 13047 45067
rect 12989 45027 13047 45033
rect 16390 45024 16396 45076
rect 16448 45064 16454 45076
rect 17129 45067 17187 45073
rect 17129 45064 17141 45067
rect 16448 45036 17141 45064
rect 16448 45024 16454 45036
rect 17129 45033 17141 45036
rect 17175 45033 17187 45067
rect 17129 45027 17187 45033
rect 4706 44956 4712 45008
rect 4764 44996 4770 45008
rect 7929 44999 7987 45005
rect 7929 44996 7941 44999
rect 4764 44968 7941 44996
rect 4764 44956 4770 44968
rect 7929 44965 7941 44968
rect 7975 44965 7987 44999
rect 7929 44959 7987 44965
rect 12618 44888 12624 44940
rect 12676 44928 12682 44940
rect 13541 44931 13599 44937
rect 13541 44928 13553 44931
rect 12676 44900 13553 44928
rect 12676 44888 12682 44900
rect 13541 44897 13553 44900
rect 13587 44928 13599 44931
rect 13722 44928 13728 44940
rect 13587 44900 13728 44928
rect 13587 44897 13599 44900
rect 13541 44891 13599 44897
rect 13722 44888 13728 44900
rect 13780 44888 13786 44940
rect 16850 44928 16856 44940
rect 15120 44900 16856 44928
rect 13357 44863 13415 44869
rect 13357 44829 13369 44863
rect 13403 44860 13415 44863
rect 13446 44860 13452 44872
rect 13403 44832 13452 44860
rect 13403 44829 13415 44832
rect 13357 44823 13415 44829
rect 13446 44820 13452 44832
rect 13504 44820 13510 44872
rect 14826 44820 14832 44872
rect 14884 44860 14890 44872
rect 15120 44869 15148 44900
rect 16850 44888 16856 44900
rect 16908 44888 16914 44940
rect 21634 44888 21640 44940
rect 21692 44928 21698 44940
rect 21692 44900 23796 44928
rect 21692 44888 21698 44900
rect 15105 44863 15163 44869
rect 15105 44860 15117 44863
rect 14884 44832 15117 44860
rect 14884 44820 14890 44832
rect 15105 44829 15117 44832
rect 15151 44829 15163 44863
rect 15105 44823 15163 44829
rect 16758 44820 16764 44872
rect 16816 44860 16822 44872
rect 16942 44860 16948 44872
rect 16816 44832 16948 44860
rect 16816 44820 16822 44832
rect 16942 44820 16948 44832
rect 17000 44820 17006 44872
rect 19518 44820 19524 44872
rect 19576 44820 19582 44872
rect 20898 44820 20904 44872
rect 20956 44860 20962 44872
rect 21652 44860 21680 44888
rect 20956 44832 21680 44860
rect 20956 44820 20962 44832
rect 22278 44820 22284 44872
rect 22336 44820 22342 44872
rect 7745 44795 7803 44801
rect 7745 44761 7757 44795
rect 7791 44792 7803 44795
rect 9217 44795 9275 44801
rect 7791 44764 8340 44792
rect 7791 44761 7803 44764
rect 7745 44755 7803 44761
rect 6457 44727 6515 44733
rect 6457 44693 6469 44727
rect 6503 44724 6515 44727
rect 6638 44724 6644 44736
rect 6503 44696 6644 44724
rect 6503 44693 6515 44696
rect 6457 44687 6515 44693
rect 6638 44684 6644 44696
rect 6696 44684 6702 44736
rect 7193 44727 7251 44733
rect 7193 44693 7205 44727
rect 7239 44724 7251 44727
rect 7282 44724 7288 44736
rect 7239 44696 7288 44724
rect 7239 44693 7251 44696
rect 7193 44687 7251 44693
rect 7282 44684 7288 44696
rect 7340 44684 7346 44736
rect 8312 44733 8340 44764
rect 9217 44761 9229 44795
rect 9263 44792 9275 44795
rect 11149 44795 11207 44801
rect 9263 44764 9812 44792
rect 9263 44761 9275 44764
rect 9217 44755 9275 44761
rect 9784 44736 9812 44764
rect 11149 44761 11161 44795
rect 11195 44792 11207 44795
rect 11517 44795 11575 44801
rect 11517 44792 11529 44795
rect 11195 44764 11529 44792
rect 11195 44761 11207 44764
rect 11149 44755 11207 44761
rect 11517 44761 11529 44764
rect 11563 44792 11575 44795
rect 12345 44795 12403 44801
rect 11563 44764 12112 44792
rect 11563 44761 11575 44764
rect 11517 44755 11575 44761
rect 8297 44727 8355 44733
rect 8297 44693 8309 44727
rect 8343 44724 8355 44727
rect 8662 44724 8668 44736
rect 8343 44696 8668 44724
rect 8343 44693 8355 44696
rect 8297 44687 8355 44693
rect 8662 44684 8668 44696
rect 8720 44684 8726 44736
rect 9766 44684 9772 44736
rect 9824 44684 9830 44736
rect 12084 44724 12112 44764
rect 12345 44761 12357 44795
rect 12391 44792 12403 44795
rect 12434 44792 12440 44804
rect 12391 44764 12440 44792
rect 12391 44761 12403 44764
rect 12345 44755 12403 44761
rect 12434 44752 12440 44764
rect 12492 44752 12498 44804
rect 15381 44795 15439 44801
rect 15381 44761 15393 44795
rect 15427 44792 15439 44795
rect 15654 44792 15660 44804
rect 15427 44764 15660 44792
rect 15427 44761 15439 44764
rect 15381 44755 15439 44761
rect 15654 44752 15660 44764
rect 15712 44752 15718 44804
rect 15838 44752 15844 44804
rect 15896 44752 15902 44804
rect 19794 44752 19800 44804
rect 19852 44752 19858 44804
rect 22554 44752 22560 44804
rect 22612 44752 22618 44804
rect 23768 44792 23796 44900
rect 23768 44778 24348 44792
rect 23782 44764 24348 44778
rect 24320 44736 24348 44764
rect 12526 44724 12532 44736
rect 12084 44696 12532 44724
rect 12526 44684 12532 44696
rect 12584 44684 12590 44736
rect 13449 44727 13507 44733
rect 13449 44693 13461 44727
rect 13495 44724 13507 44727
rect 15194 44724 15200 44736
rect 13495 44696 15200 44724
rect 13495 44693 13507 44696
rect 13449 44687 13507 44693
rect 15194 44684 15200 44696
rect 15252 44684 15258 44736
rect 16853 44727 16911 44733
rect 16853 44693 16865 44727
rect 16899 44724 16911 44727
rect 17218 44724 17224 44736
rect 16899 44696 17224 44724
rect 16899 44693 16911 44696
rect 16853 44687 16911 44693
rect 17218 44684 17224 44696
rect 17276 44684 17282 44736
rect 19978 44684 19984 44736
rect 20036 44724 20042 44736
rect 21269 44727 21327 44733
rect 21269 44724 21281 44727
rect 20036 44696 21281 44724
rect 20036 44684 20042 44696
rect 21269 44693 21281 44696
rect 21315 44693 21327 44727
rect 21269 44687 21327 44693
rect 23382 44684 23388 44736
rect 23440 44724 23446 44736
rect 24029 44727 24087 44733
rect 24029 44724 24041 44727
rect 23440 44696 24041 44724
rect 23440 44684 23446 44696
rect 24029 44693 24041 44696
rect 24075 44693 24087 44727
rect 24029 44687 24087 44693
rect 24302 44684 24308 44736
rect 24360 44724 24366 44736
rect 24397 44727 24455 44733
rect 24397 44724 24409 44727
rect 24360 44696 24409 44724
rect 24360 44684 24366 44696
rect 24397 44693 24409 44696
rect 24443 44693 24455 44727
rect 24397 44687 24455 44693
rect 24486 44684 24492 44736
rect 24544 44724 24550 44736
rect 25498 44724 25504 44736
rect 24544 44696 25504 44724
rect 24544 44684 24550 44696
rect 25498 44684 25504 44696
rect 25556 44684 25562 44736
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 5810 44480 5816 44532
rect 5868 44480 5874 44532
rect 6730 44480 6736 44532
rect 6788 44480 6794 44532
rect 7374 44480 7380 44532
rect 7432 44520 7438 44532
rect 7469 44523 7527 44529
rect 7469 44520 7481 44523
rect 7432 44492 7481 44520
rect 7432 44480 7438 44492
rect 7469 44489 7481 44492
rect 7515 44489 7527 44523
rect 7469 44483 7527 44489
rect 7834 44480 7840 44532
rect 7892 44520 7898 44532
rect 8021 44523 8079 44529
rect 8021 44520 8033 44523
rect 7892 44492 8033 44520
rect 7892 44480 7898 44492
rect 8021 44489 8033 44492
rect 8067 44489 8079 44523
rect 8021 44483 8079 44489
rect 9674 44480 9680 44532
rect 9732 44520 9738 44532
rect 11057 44523 11115 44529
rect 11057 44520 11069 44523
rect 9732 44492 11069 44520
rect 9732 44480 9738 44492
rect 11057 44489 11069 44492
rect 11103 44489 11115 44523
rect 11057 44483 11115 44489
rect 11146 44480 11152 44532
rect 11204 44520 11210 44532
rect 11885 44523 11943 44529
rect 11885 44520 11897 44523
rect 11204 44492 11897 44520
rect 11204 44480 11210 44492
rect 11885 44489 11897 44492
rect 11931 44489 11943 44523
rect 11885 44483 11943 44489
rect 12253 44523 12311 44529
rect 12253 44489 12265 44523
rect 12299 44520 12311 44523
rect 16390 44520 16396 44532
rect 12299 44492 16396 44520
rect 12299 44489 12311 44492
rect 12253 44483 12311 44489
rect 16390 44480 16396 44492
rect 16448 44480 16454 44532
rect 18874 44520 18880 44532
rect 17512 44492 18880 44520
rect 7098 44412 7104 44464
rect 7156 44452 7162 44464
rect 9125 44455 9183 44461
rect 9125 44452 9137 44455
rect 7156 44424 9137 44452
rect 7156 44412 7162 44424
rect 9125 44421 9137 44424
rect 9171 44421 9183 44455
rect 9125 44415 9183 44421
rect 12342 44412 12348 44464
rect 12400 44452 12406 44464
rect 13354 44452 13360 44464
rect 12400 44424 13360 44452
rect 12400 44412 12406 44424
rect 5258 44344 5264 44396
rect 5316 44384 5322 44396
rect 5997 44387 6055 44393
rect 5997 44384 6009 44387
rect 5316 44356 6009 44384
rect 5316 44344 5322 44356
rect 5997 44353 6009 44356
rect 6043 44353 6055 44387
rect 5997 44347 6055 44353
rect 6641 44387 6699 44393
rect 6641 44353 6653 44387
rect 6687 44384 6699 44387
rect 6730 44384 6736 44396
rect 6687 44356 6736 44384
rect 6687 44353 6699 44356
rect 6641 44347 6699 44353
rect 6730 44344 6736 44356
rect 6788 44344 6794 44396
rect 7374 44344 7380 44396
rect 7432 44344 7438 44396
rect 7466 44344 7472 44396
rect 7524 44384 7530 44396
rect 8205 44387 8263 44393
rect 8205 44384 8217 44387
rect 7524 44356 8217 44384
rect 7524 44344 7530 44356
rect 8205 44353 8217 44356
rect 8251 44353 8263 44387
rect 8205 44347 8263 44353
rect 8938 44344 8944 44396
rect 8996 44384 9002 44396
rect 13188 44393 13216 44424
rect 13354 44412 13360 44424
rect 13412 44412 13418 44464
rect 13998 44412 14004 44464
rect 14056 44412 14062 44464
rect 15102 44412 15108 44464
rect 15160 44452 15166 44464
rect 15381 44455 15439 44461
rect 15381 44452 15393 44455
rect 15160 44424 15393 44452
rect 15160 44412 15166 44424
rect 15381 44421 15393 44424
rect 15427 44452 15439 44455
rect 15838 44452 15844 44464
rect 15427 44424 15844 44452
rect 15427 44421 15439 44424
rect 15381 44415 15439 44421
rect 15838 44412 15844 44424
rect 15896 44452 15902 44464
rect 17512 44452 17540 44492
rect 18874 44480 18880 44492
rect 18932 44480 18938 44532
rect 19794 44480 19800 44532
rect 19852 44520 19858 44532
rect 20438 44520 20444 44532
rect 19852 44492 20444 44520
rect 19852 44480 19858 44492
rect 20438 44480 20444 44492
rect 20496 44520 20502 44532
rect 21269 44523 21327 44529
rect 21269 44520 21281 44523
rect 20496 44492 21281 44520
rect 20496 44480 20502 44492
rect 21269 44489 21281 44492
rect 21315 44489 21327 44523
rect 21269 44483 21327 44489
rect 21634 44480 21640 44532
rect 21692 44480 21698 44532
rect 22554 44480 22560 44532
rect 22612 44520 22618 44532
rect 24029 44523 24087 44529
rect 24029 44520 24041 44523
rect 22612 44492 24041 44520
rect 22612 44480 22618 44492
rect 24029 44489 24041 44492
rect 24075 44489 24087 44523
rect 24029 44483 24087 44489
rect 21652 44452 21680 44480
rect 24302 44452 24308 44464
rect 15896 44424 17618 44452
rect 21022 44424 21680 44452
rect 23782 44424 24308 44452
rect 15896 44412 15902 44424
rect 24302 44412 24308 44424
rect 24360 44412 24366 44464
rect 9401 44387 9459 44393
rect 9401 44384 9413 44387
rect 8996 44356 9413 44384
rect 8996 44344 9002 44356
rect 9401 44353 9413 44356
rect 9447 44353 9459 44387
rect 9401 44347 9459 44353
rect 10965 44387 11023 44393
rect 10965 44353 10977 44387
rect 11011 44384 11023 44387
rect 13173 44387 13231 44393
rect 11011 44356 11652 44384
rect 11011 44353 11023 44356
rect 10965 44347 11023 44353
rect 11624 44260 11652 44356
rect 13173 44353 13185 44387
rect 13219 44353 13231 44387
rect 13173 44347 13231 44353
rect 24489 44387 24547 44393
rect 24489 44353 24501 44387
rect 24535 44384 24547 44387
rect 25314 44384 25320 44396
rect 24535 44356 25320 44384
rect 24535 44353 24547 44356
rect 24489 44347 24547 44353
rect 25314 44344 25320 44356
rect 25372 44344 25378 44396
rect 11698 44276 11704 44328
rect 11756 44316 11762 44328
rect 12345 44319 12403 44325
rect 12345 44316 12357 44319
rect 11756 44288 12357 44316
rect 11756 44276 11762 44288
rect 12345 44285 12357 44288
rect 12391 44285 12403 44319
rect 12345 44279 12403 44285
rect 12437 44319 12495 44325
rect 12437 44285 12449 44319
rect 12483 44285 12495 44319
rect 12437 44279 12495 44285
rect 11606 44208 11612 44260
rect 11664 44208 11670 44260
rect 12250 44208 12256 44260
rect 12308 44248 12314 44260
rect 12452 44248 12480 44279
rect 14182 44276 14188 44328
rect 14240 44316 14246 44328
rect 14921 44319 14979 44325
rect 14921 44316 14933 44319
rect 14240 44288 14933 44316
rect 14240 44276 14246 44288
rect 14921 44285 14933 44288
rect 14967 44285 14979 44319
rect 14921 44279 14979 44285
rect 16850 44276 16856 44328
rect 16908 44276 16914 44328
rect 17129 44319 17187 44325
rect 17129 44285 17141 44319
rect 17175 44316 17187 44319
rect 18966 44316 18972 44328
rect 17175 44288 18972 44316
rect 17175 44285 17187 44288
rect 17129 44279 17187 44285
rect 18966 44276 18972 44288
rect 19024 44276 19030 44328
rect 19518 44276 19524 44328
rect 19576 44316 19582 44328
rect 19797 44319 19855 44325
rect 19576 44288 19656 44316
rect 19576 44276 19582 44288
rect 12308 44220 12480 44248
rect 12308 44208 12314 44220
rect 13436 44183 13494 44189
rect 13436 44149 13448 44183
rect 13482 44180 13494 44183
rect 13630 44180 13636 44192
rect 13482 44152 13636 44180
rect 13482 44149 13494 44152
rect 13436 44143 13494 44149
rect 13630 44140 13636 44152
rect 13688 44180 13694 44192
rect 15197 44183 15255 44189
rect 15197 44180 15209 44183
rect 13688 44152 15209 44180
rect 13688 44140 13694 44152
rect 15197 44149 15209 44152
rect 15243 44180 15255 44183
rect 16482 44180 16488 44192
rect 15243 44152 16488 44180
rect 15243 44149 15255 44152
rect 15197 44143 15255 44149
rect 16482 44140 16488 44152
rect 16540 44140 16546 44192
rect 16868 44180 16896 44276
rect 18322 44180 18328 44192
rect 16868 44152 18328 44180
rect 18322 44140 18328 44152
rect 18380 44140 18386 44192
rect 18598 44140 18604 44192
rect 18656 44180 18662 44192
rect 18782 44180 18788 44192
rect 18656 44152 18788 44180
rect 18656 44140 18662 44152
rect 18782 44140 18788 44152
rect 18840 44140 18846 44192
rect 19628 44180 19656 44288
rect 19797 44285 19809 44319
rect 19843 44316 19855 44319
rect 20806 44316 20812 44328
rect 19843 44288 20812 44316
rect 19843 44285 19855 44288
rect 19797 44279 19855 44285
rect 20806 44276 20812 44288
rect 20864 44276 20870 44328
rect 22278 44276 22284 44328
rect 22336 44316 22342 44328
rect 22557 44319 22615 44325
rect 22336 44288 22416 44316
rect 22336 44276 22342 44288
rect 22388 44180 22416 44288
rect 22557 44285 22569 44319
rect 22603 44316 22615 44319
rect 22646 44316 22652 44328
rect 22603 44288 22652 44316
rect 22603 44285 22615 44288
rect 22557 44279 22615 44285
rect 22646 44276 22652 44288
rect 22704 44276 22710 44328
rect 24762 44276 24768 44328
rect 24820 44276 24826 44328
rect 23290 44180 23296 44192
rect 19628 44152 23296 44180
rect 23290 44140 23296 44152
rect 23348 44140 23354 44192
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 8389 43979 8447 43985
rect 8389 43945 8401 43979
rect 8435 43976 8447 43979
rect 9398 43976 9404 43988
rect 8435 43948 9404 43976
rect 8435 43945 8447 43948
rect 8389 43939 8447 43945
rect 9398 43936 9404 43948
rect 9456 43936 9462 43988
rect 11330 43936 11336 43988
rect 11388 43976 11394 43988
rect 11609 43979 11667 43985
rect 11609 43976 11621 43979
rect 11388 43948 11621 43976
rect 11388 43936 11394 43948
rect 11609 43945 11621 43948
rect 11655 43945 11667 43979
rect 11609 43939 11667 43945
rect 23290 43936 23296 43988
rect 23348 43976 23354 43988
rect 23474 43976 23480 43988
rect 23348 43948 23480 43976
rect 23348 43936 23354 43948
rect 23474 43936 23480 43948
rect 23532 43936 23538 43988
rect 6917 43911 6975 43917
rect 6917 43877 6929 43911
rect 6963 43908 6975 43911
rect 7006 43908 7012 43920
rect 6963 43880 7012 43908
rect 6963 43877 6975 43880
rect 6917 43871 6975 43877
rect 7006 43868 7012 43880
rect 7064 43868 7070 43920
rect 9125 43843 9183 43849
rect 9125 43809 9137 43843
rect 9171 43840 9183 43843
rect 9398 43840 9404 43852
rect 9171 43812 9404 43840
rect 9171 43809 9183 43812
rect 9125 43803 9183 43809
rect 9398 43800 9404 43812
rect 9456 43800 9462 43852
rect 22462 43800 22468 43852
rect 22520 43800 22526 43852
rect 22649 43843 22707 43849
rect 22649 43809 22661 43843
rect 22695 43840 22707 43843
rect 23290 43840 23296 43852
rect 22695 43812 23296 43840
rect 22695 43809 22707 43812
rect 22649 43803 22707 43809
rect 23290 43800 23296 43812
rect 23348 43800 23354 43852
rect 8478 43732 8484 43784
rect 8536 43772 8542 43784
rect 8573 43775 8631 43781
rect 8573 43772 8585 43775
rect 8536 43744 8585 43772
rect 8536 43732 8542 43744
rect 8573 43741 8585 43744
rect 8619 43741 8631 43775
rect 15470 43772 15476 43784
rect 8573 43735 8631 43741
rect 10796 43744 15476 43772
rect 6733 43707 6791 43713
rect 6733 43673 6745 43707
rect 6779 43704 6791 43707
rect 9401 43707 9459 43713
rect 6779 43676 7144 43704
rect 6779 43673 6791 43676
rect 6733 43667 6791 43673
rect 7116 43648 7144 43676
rect 9401 43673 9413 43707
rect 9447 43673 9459 43707
rect 9401 43667 9459 43673
rect 1210 43596 1216 43648
rect 1268 43636 1274 43648
rect 1397 43639 1455 43645
rect 1397 43636 1409 43639
rect 1268 43608 1409 43636
rect 1268 43596 1274 43608
rect 1397 43605 1409 43608
rect 1443 43605 1455 43639
rect 1397 43599 1455 43605
rect 7098 43596 7104 43648
rect 7156 43636 7162 43648
rect 7193 43639 7251 43645
rect 7193 43636 7205 43639
rect 7156 43608 7205 43636
rect 7156 43596 7162 43608
rect 7193 43605 7205 43608
rect 7239 43605 7251 43639
rect 9416 43636 9444 43667
rect 10042 43664 10048 43716
rect 10100 43664 10106 43716
rect 10796 43636 10824 43744
rect 15470 43732 15476 43744
rect 15528 43732 15534 43784
rect 11517 43707 11575 43713
rect 11517 43673 11529 43707
rect 11563 43704 11575 43707
rect 25409 43707 25467 43713
rect 25409 43704 25421 43707
rect 11563 43676 12112 43704
rect 11563 43673 11575 43676
rect 11517 43667 11575 43673
rect 12084 43648 12112 43676
rect 24320 43676 25421 43704
rect 24320 43648 24348 43676
rect 25409 43673 25421 43676
rect 25455 43673 25467 43707
rect 25409 43667 25467 43673
rect 9416 43608 10824 43636
rect 10873 43639 10931 43645
rect 7193 43599 7251 43605
rect 10873 43605 10885 43639
rect 10919 43636 10931 43639
rect 10962 43636 10968 43648
rect 10919 43608 10968 43636
rect 10919 43605 10931 43608
rect 10873 43599 10931 43605
rect 10962 43596 10968 43608
rect 11020 43596 11026 43648
rect 12066 43596 12072 43648
rect 12124 43596 12130 43648
rect 17402 43596 17408 43648
rect 17460 43636 17466 43648
rect 17957 43639 18015 43645
rect 17957 43636 17969 43639
rect 17460 43608 17969 43636
rect 17460 43596 17466 43608
rect 17957 43605 17969 43608
rect 18003 43636 18015 43639
rect 20254 43636 20260 43648
rect 18003 43608 20260 43636
rect 18003 43605 18015 43608
rect 17957 43599 18015 43605
rect 20254 43596 20260 43608
rect 20312 43596 20318 43648
rect 21910 43596 21916 43648
rect 21968 43636 21974 43648
rect 22005 43639 22063 43645
rect 22005 43636 22017 43639
rect 21968 43608 22017 43636
rect 21968 43596 21974 43608
rect 22005 43605 22017 43608
rect 22051 43605 22063 43639
rect 22005 43599 22063 43605
rect 22373 43639 22431 43645
rect 22373 43605 22385 43639
rect 22419 43636 22431 43639
rect 22462 43636 22468 43648
rect 22419 43608 22468 43636
rect 22419 43605 22431 43608
rect 22373 43599 22431 43605
rect 22462 43596 22468 43608
rect 22520 43636 22526 43648
rect 22830 43636 22836 43648
rect 22520 43608 22836 43636
rect 22520 43596 22526 43608
rect 22830 43596 22836 43608
rect 22888 43636 22894 43648
rect 23017 43639 23075 43645
rect 23017 43636 23029 43639
rect 22888 43608 23029 43636
rect 22888 43596 22894 43608
rect 23017 43605 23029 43608
rect 23063 43605 23075 43639
rect 23017 43599 23075 43605
rect 24213 43639 24271 43645
rect 24213 43605 24225 43639
rect 24259 43636 24271 43639
rect 24302 43636 24308 43648
rect 24259 43608 24308 43636
rect 24259 43605 24271 43608
rect 24213 43599 24271 43605
rect 24302 43596 24308 43608
rect 24360 43596 24366 43648
rect 25314 43596 25320 43648
rect 25372 43596 25378 43648
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 7742 43392 7748 43444
rect 7800 43392 7806 43444
rect 8570 43392 8576 43444
rect 8628 43432 8634 43444
rect 9493 43435 9551 43441
rect 9493 43432 9505 43435
rect 8628 43404 9505 43432
rect 8628 43392 8634 43404
rect 9493 43401 9505 43404
rect 9539 43432 9551 43435
rect 9582 43432 9588 43444
rect 9539 43404 9588 43432
rect 9539 43401 9551 43404
rect 9493 43395 9551 43401
rect 9582 43392 9588 43404
rect 9640 43392 9646 43444
rect 10410 43392 10416 43444
rect 10468 43432 10474 43444
rect 10597 43435 10655 43441
rect 10597 43432 10609 43435
rect 10468 43404 10609 43432
rect 10468 43392 10474 43404
rect 10597 43401 10609 43404
rect 10643 43401 10655 43435
rect 10597 43395 10655 43401
rect 15010 43392 15016 43444
rect 15068 43392 15074 43444
rect 17402 43392 17408 43444
rect 17460 43392 17466 43444
rect 17494 43392 17500 43444
rect 17552 43392 17558 43444
rect 20070 43392 20076 43444
rect 20128 43392 20134 43444
rect 20441 43435 20499 43441
rect 20441 43401 20453 43435
rect 20487 43432 20499 43435
rect 21358 43432 21364 43444
rect 20487 43404 21364 43432
rect 20487 43401 20499 43404
rect 20441 43395 20499 43401
rect 4614 43324 4620 43376
rect 4672 43364 4678 43376
rect 8665 43367 8723 43373
rect 8665 43364 8677 43367
rect 4672 43336 8677 43364
rect 4672 43324 4678 43336
rect 8665 43333 8677 43336
rect 8711 43333 8723 43367
rect 8665 43327 8723 43333
rect 10042 43324 10048 43376
rect 10100 43364 10106 43376
rect 11057 43367 11115 43373
rect 11057 43364 11069 43367
rect 10100 43336 11069 43364
rect 10100 43324 10106 43336
rect 11057 43333 11069 43336
rect 11103 43333 11115 43367
rect 11057 43327 11115 43333
rect 12618 43324 12624 43376
rect 12676 43324 12682 43376
rect 13998 43364 14004 43376
rect 13846 43336 14004 43364
rect 13998 43324 14004 43336
rect 14056 43324 14062 43376
rect 20456 43364 20484 43395
rect 21358 43392 21364 43404
rect 21416 43432 21422 43444
rect 21453 43435 21511 43441
rect 21453 43432 21465 43435
rect 21416 43404 21465 43432
rect 21416 43392 21422 43404
rect 21453 43401 21465 43404
rect 21499 43432 21511 43435
rect 21634 43432 21640 43444
rect 21499 43404 21640 43432
rect 21499 43401 21511 43404
rect 21453 43395 21511 43401
rect 21634 43392 21640 43404
rect 21692 43392 21698 43444
rect 22370 43392 22376 43444
rect 22428 43432 22434 43444
rect 22465 43435 22523 43441
rect 22465 43432 22477 43435
rect 22428 43404 22477 43432
rect 22428 43392 22434 43404
rect 22465 43401 22477 43404
rect 22511 43401 22523 43435
rect 22465 43395 22523 43401
rect 15028 43336 15424 43364
rect 19826 43336 20484 43364
rect 1210 43256 1216 43308
rect 1268 43296 1274 43308
rect 1581 43299 1639 43305
rect 1581 43296 1593 43299
rect 1268 43268 1593 43296
rect 1268 43256 1274 43268
rect 1581 43265 1593 43268
rect 1627 43265 1639 43299
rect 1581 43259 1639 43265
rect 7650 43256 7656 43308
rect 7708 43296 7714 43308
rect 7929 43299 7987 43305
rect 7929 43296 7941 43299
rect 7708 43268 7941 43296
rect 7708 43256 7714 43268
rect 7929 43265 7941 43268
rect 7975 43265 7987 43299
rect 7929 43259 7987 43265
rect 8386 43256 8392 43308
rect 8444 43296 8450 43308
rect 8481 43299 8539 43305
rect 8481 43296 8493 43299
rect 8444 43268 8493 43296
rect 8444 43256 8450 43268
rect 8481 43265 8493 43268
rect 8527 43265 8539 43299
rect 8481 43259 8539 43265
rect 9490 43256 9496 43308
rect 9548 43296 9554 43308
rect 9585 43299 9643 43305
rect 9585 43296 9597 43299
rect 9548 43268 9597 43296
rect 9548 43256 9554 43268
rect 9585 43265 9597 43268
rect 9631 43265 9643 43299
rect 9585 43259 9643 43265
rect 10318 43256 10324 43308
rect 10376 43296 10382 43308
rect 10505 43299 10563 43305
rect 10505 43296 10517 43299
rect 10376 43268 10517 43296
rect 10376 43256 10382 43268
rect 10505 43265 10517 43268
rect 10551 43265 10563 43299
rect 10505 43259 10563 43265
rect 12342 43256 12348 43308
rect 12400 43256 12406 43308
rect 8846 43188 8852 43240
rect 8904 43228 8910 43240
rect 9677 43231 9735 43237
rect 9677 43228 9689 43231
rect 8904 43200 9689 43228
rect 8904 43188 8910 43200
rect 9677 43197 9689 43200
rect 9723 43228 9735 43231
rect 15028 43228 15056 43336
rect 15105 43299 15163 43305
rect 15105 43265 15117 43299
rect 15151 43296 15163 43299
rect 15151 43268 15332 43296
rect 15151 43265 15163 43268
rect 15105 43259 15163 43265
rect 9723 43200 15056 43228
rect 15197 43231 15255 43237
rect 9723 43197 9735 43200
rect 9677 43191 9735 43197
rect 15197 43197 15209 43231
rect 15243 43197 15255 43231
rect 15197 43191 15255 43197
rect 9125 43163 9183 43169
rect 9125 43129 9137 43163
rect 9171 43160 9183 43163
rect 11698 43160 11704 43172
rect 9171 43132 11704 43160
rect 9171 43129 9183 43132
rect 9125 43123 9183 43129
rect 11698 43120 11704 43132
rect 11756 43120 11762 43172
rect 14918 43120 14924 43172
rect 14976 43160 14982 43172
rect 15212 43160 15240 43191
rect 14976 43132 15240 43160
rect 14976 43120 14982 43132
rect 2222 43052 2228 43104
rect 2280 43052 2286 43104
rect 13998 43052 14004 43104
rect 14056 43092 14062 43104
rect 14093 43095 14151 43101
rect 14093 43092 14105 43095
rect 14056 43064 14105 43092
rect 14056 43052 14062 43064
rect 14093 43061 14105 43064
rect 14139 43061 14151 43095
rect 14093 43055 14151 43061
rect 14182 43052 14188 43104
rect 14240 43092 14246 43104
rect 14645 43095 14703 43101
rect 14645 43092 14657 43095
rect 14240 43064 14657 43092
rect 14240 43052 14246 43064
rect 14645 43061 14657 43064
rect 14691 43061 14703 43095
rect 15304 43092 15332 43268
rect 15396 43160 15424 43336
rect 24302 43324 24308 43376
rect 24360 43324 24366 43376
rect 21634 43256 21640 43308
rect 21692 43296 21698 43308
rect 22373 43299 22431 43305
rect 22373 43296 22385 43299
rect 21692 43268 22385 43296
rect 21692 43256 21698 43268
rect 22373 43265 22385 43268
rect 22419 43265 22431 43299
rect 22373 43259 22431 43265
rect 15654 43188 15660 43240
rect 15712 43228 15718 43240
rect 17310 43228 17316 43240
rect 15712 43200 17316 43228
rect 15712 43188 15718 43200
rect 17310 43188 17316 43200
rect 17368 43228 17374 43240
rect 17589 43231 17647 43237
rect 17589 43228 17601 43231
rect 17368 43200 17601 43228
rect 17368 43188 17374 43200
rect 17589 43197 17601 43200
rect 17635 43197 17647 43231
rect 17589 43191 17647 43197
rect 18322 43188 18328 43240
rect 18380 43188 18386 43240
rect 18601 43231 18659 43237
rect 18601 43197 18613 43231
rect 18647 43228 18659 43231
rect 19978 43228 19984 43240
rect 18647 43200 19984 43228
rect 18647 43197 18659 43200
rect 18601 43191 18659 43197
rect 19978 43188 19984 43200
rect 20036 43188 20042 43240
rect 22646 43188 22652 43240
rect 22704 43188 22710 43240
rect 23474 43188 23480 43240
rect 23532 43228 23538 43240
rect 23569 43231 23627 43237
rect 23569 43228 23581 43231
rect 23532 43200 23581 43228
rect 23532 43188 23538 43200
rect 23569 43197 23581 43200
rect 23615 43197 23627 43231
rect 23569 43191 23627 43197
rect 23842 43188 23848 43240
rect 23900 43188 23906 43240
rect 18138 43160 18144 43172
rect 15396 43132 18144 43160
rect 18138 43120 18144 43132
rect 18196 43120 18202 43172
rect 15562 43092 15568 43104
rect 15304 43064 15568 43092
rect 14645 43055 14703 43061
rect 15562 43052 15568 43064
rect 15620 43092 15626 43104
rect 15749 43095 15807 43101
rect 15749 43092 15761 43095
rect 15620 43064 15761 43092
rect 15620 43052 15626 43064
rect 15749 43061 15761 43064
rect 15795 43092 15807 43095
rect 15838 43092 15844 43104
rect 15795 43064 15844 43092
rect 15795 43061 15807 43064
rect 15749 43055 15807 43061
rect 15838 43052 15844 43064
rect 15896 43052 15902 43104
rect 16666 43052 16672 43104
rect 16724 43052 16730 43104
rect 17034 43052 17040 43104
rect 17092 43052 17098 43104
rect 18340 43092 18368 43188
rect 19242 43092 19248 43104
rect 18340 43064 19248 43092
rect 19242 43052 19248 43064
rect 19300 43052 19306 43104
rect 21634 43052 21640 43104
rect 21692 43052 21698 43104
rect 22005 43095 22063 43101
rect 22005 43061 22017 43095
rect 22051 43092 22063 43095
rect 24946 43092 24952 43104
rect 22051 43064 24952 43092
rect 22051 43061 22063 43064
rect 22005 43055 22063 43061
rect 24946 43052 24952 43064
rect 25004 43052 25010 43104
rect 25222 43052 25228 43104
rect 25280 43092 25286 43104
rect 25317 43095 25375 43101
rect 25317 43092 25329 43095
rect 25280 43064 25329 43092
rect 25280 43052 25286 43064
rect 25317 43061 25329 43064
rect 25363 43061 25375 43095
rect 25317 43055 25375 43061
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 8570 42848 8576 42900
rect 8628 42848 8634 42900
rect 8846 42888 8852 42900
rect 8680 42860 8852 42888
rect 4890 42712 4896 42764
rect 4948 42752 4954 42764
rect 4985 42755 5043 42761
rect 4985 42752 4997 42755
rect 4948 42724 4997 42752
rect 4948 42712 4954 42724
rect 4985 42721 4997 42724
rect 5031 42721 5043 42755
rect 4985 42715 5043 42721
rect 8570 42712 8576 42764
rect 8628 42752 8634 42764
rect 8680 42752 8708 42860
rect 8846 42848 8852 42860
rect 8904 42888 8910 42900
rect 8941 42891 8999 42897
rect 8941 42888 8953 42891
rect 8904 42860 8953 42888
rect 8904 42848 8910 42860
rect 8941 42857 8953 42860
rect 8987 42857 8999 42891
rect 8941 42851 8999 42857
rect 9217 42891 9275 42897
rect 9217 42857 9229 42891
rect 9263 42888 9275 42891
rect 9306 42888 9312 42900
rect 9263 42860 9312 42888
rect 9263 42857 9275 42860
rect 9217 42851 9275 42857
rect 9306 42848 9312 42860
rect 9364 42888 9370 42900
rect 9490 42888 9496 42900
rect 9364 42860 9496 42888
rect 9364 42848 9370 42860
rect 9490 42848 9496 42860
rect 9548 42848 9554 42900
rect 12158 42848 12164 42900
rect 12216 42888 12222 42900
rect 12897 42891 12955 42897
rect 12897 42888 12909 42891
rect 12216 42860 12909 42888
rect 12216 42848 12222 42860
rect 12897 42857 12909 42860
rect 12943 42888 12955 42891
rect 13906 42888 13912 42900
rect 12943 42860 13912 42888
rect 12943 42857 12955 42860
rect 12897 42851 12955 42857
rect 13906 42848 13912 42860
rect 13964 42888 13970 42900
rect 14277 42891 14335 42897
rect 14277 42888 14289 42891
rect 13964 42860 14289 42888
rect 13964 42848 13970 42860
rect 14277 42857 14289 42860
rect 14323 42888 14335 42891
rect 15562 42888 15568 42900
rect 14323 42860 15568 42888
rect 14323 42857 14335 42860
rect 14277 42851 14335 42857
rect 15562 42848 15568 42860
rect 15620 42888 15626 42900
rect 15838 42888 15844 42900
rect 15620 42860 15844 42888
rect 15620 42848 15626 42860
rect 15838 42848 15844 42860
rect 15896 42888 15902 42900
rect 16666 42888 16672 42900
rect 15896 42860 16672 42888
rect 15896 42848 15902 42860
rect 16666 42848 16672 42860
rect 16724 42848 16730 42900
rect 19784 42891 19842 42897
rect 19784 42857 19796 42891
rect 19830 42888 19842 42891
rect 20346 42888 20352 42900
rect 19830 42860 20352 42888
rect 19830 42857 19842 42860
rect 19784 42851 19842 42857
rect 20346 42848 20352 42860
rect 20404 42888 20410 42900
rect 21726 42888 21732 42900
rect 20404 42860 21732 42888
rect 20404 42848 20410 42860
rect 21726 42848 21732 42860
rect 21784 42848 21790 42900
rect 8628 42724 8708 42752
rect 8628 42712 8634 42724
rect 9214 42712 9220 42764
rect 9272 42752 9278 42764
rect 9309 42755 9367 42761
rect 9309 42752 9321 42755
rect 9272 42724 9321 42752
rect 9272 42712 9278 42724
rect 9309 42721 9321 42724
rect 9355 42721 9367 42755
rect 9309 42715 9367 42721
rect 9398 42712 9404 42764
rect 9456 42752 9462 42764
rect 10781 42755 10839 42761
rect 10781 42752 10793 42755
rect 9456 42724 10793 42752
rect 9456 42712 9462 42724
rect 10781 42721 10793 42724
rect 10827 42752 10839 42755
rect 12342 42752 12348 42764
rect 10827 42724 12348 42752
rect 10827 42721 10839 42724
rect 10781 42715 10839 42721
rect 12342 42712 12348 42724
rect 12400 42712 12406 42764
rect 14826 42712 14832 42764
rect 14884 42712 14890 42764
rect 17773 42755 17831 42761
rect 17773 42721 17785 42755
rect 17819 42752 17831 42755
rect 18138 42752 18144 42764
rect 17819 42724 18144 42752
rect 17819 42721 17831 42724
rect 17773 42715 17831 42721
rect 18138 42712 18144 42724
rect 18196 42712 18202 42764
rect 18414 42712 18420 42764
rect 18472 42712 18478 42764
rect 19521 42755 19579 42761
rect 19521 42721 19533 42755
rect 19567 42752 19579 42755
rect 19567 42724 21772 42752
rect 19567 42721 19579 42724
rect 19521 42715 19579 42721
rect 1673 42687 1731 42693
rect 1673 42653 1685 42687
rect 1719 42684 1731 42687
rect 2222 42684 2228 42696
rect 1719 42656 2228 42684
rect 1719 42653 1731 42656
rect 1673 42647 1731 42653
rect 2222 42644 2228 42656
rect 2280 42644 2286 42696
rect 12158 42644 12164 42696
rect 12216 42644 12222 42696
rect 12434 42644 12440 42696
rect 12492 42684 12498 42696
rect 14366 42684 14372 42696
rect 12492 42656 14372 42684
rect 12492 42644 12498 42656
rect 14366 42644 14372 42656
rect 14424 42644 14430 42696
rect 17589 42687 17647 42693
rect 17589 42653 17601 42687
rect 17635 42684 17647 42687
rect 18432 42684 18460 42712
rect 21358 42684 21364 42696
rect 17635 42656 18460 42684
rect 20930 42656 21364 42684
rect 17635 42653 17647 42656
rect 17589 42647 17647 42653
rect 21358 42644 21364 42656
rect 21416 42644 21422 42696
rect 21744 42684 21772 42724
rect 22002 42712 22008 42764
rect 22060 42752 22066 42764
rect 22281 42755 22339 42761
rect 22281 42752 22293 42755
rect 22060 42724 22293 42752
rect 22060 42712 22066 42724
rect 22281 42721 22293 42724
rect 22327 42721 22339 42755
rect 22281 42715 22339 42721
rect 22465 42755 22523 42761
rect 22465 42721 22477 42755
rect 22511 42752 22523 42755
rect 22554 42752 22560 42764
rect 22511 42724 22560 42752
rect 22511 42721 22523 42724
rect 22465 42715 22523 42721
rect 22554 42712 22560 42724
rect 22612 42712 22618 42764
rect 24302 42712 24308 42764
rect 24360 42752 24366 42764
rect 25317 42755 25375 42761
rect 25317 42752 25329 42755
rect 24360 42724 25329 42752
rect 24360 42712 24366 42724
rect 25317 42721 25329 42724
rect 25363 42721 25375 42755
rect 25317 42715 25375 42721
rect 22830 42684 22836 42696
rect 21744 42656 22836 42684
rect 22830 42644 22836 42656
rect 22888 42644 22894 42696
rect 23201 42687 23259 42693
rect 23201 42653 23213 42687
rect 23247 42653 23259 42687
rect 23201 42647 23259 42653
rect 23477 42687 23535 42693
rect 23477 42653 23489 42687
rect 23523 42684 23535 42687
rect 23658 42684 23664 42696
rect 23523 42656 23664 42684
rect 23523 42653 23535 42656
rect 23477 42647 23535 42653
rect 1857 42619 1915 42625
rect 1857 42585 1869 42619
rect 1903 42616 1915 42619
rect 3970 42616 3976 42628
rect 1903 42588 3976 42616
rect 1903 42585 1915 42588
rect 1857 42579 1915 42585
rect 3970 42576 3976 42588
rect 4028 42576 4034 42628
rect 4798 42576 4804 42628
rect 4856 42616 4862 42628
rect 5261 42619 5319 42625
rect 5261 42616 5273 42619
rect 4856 42588 5273 42616
rect 4856 42576 4862 42588
rect 5261 42585 5273 42588
rect 5307 42585 5319 42619
rect 5261 42579 5319 42585
rect 7558 42576 7564 42628
rect 7616 42616 7622 42628
rect 9674 42616 9680 42628
rect 7616 42588 9680 42616
rect 7616 42576 7622 42588
rect 9674 42576 9680 42588
rect 9732 42576 9738 42628
rect 11057 42619 11115 42625
rect 11057 42616 11069 42619
rect 10888 42588 11069 42616
rect 10888 42560 10916 42588
rect 11057 42585 11069 42588
rect 11103 42585 11115 42619
rect 15105 42619 15163 42625
rect 15105 42616 15117 42619
rect 11057 42579 11115 42585
rect 12544 42588 15117 42616
rect 8297 42551 8355 42557
rect 8297 42517 8309 42551
rect 8343 42548 8355 42551
rect 8386 42548 8392 42560
rect 8343 42520 8392 42548
rect 8343 42517 8355 42520
rect 8297 42511 8355 42517
rect 8386 42508 8392 42520
rect 8444 42508 8450 42560
rect 8846 42508 8852 42560
rect 8904 42548 8910 42560
rect 9493 42551 9551 42557
rect 9493 42548 9505 42551
rect 8904 42520 9505 42548
rect 8904 42508 8910 42520
rect 9493 42517 9505 42520
rect 9539 42517 9551 42551
rect 9493 42511 9551 42517
rect 10318 42508 10324 42560
rect 10376 42508 10382 42560
rect 10870 42508 10876 42560
rect 10928 42508 10934 42560
rect 12434 42508 12440 42560
rect 12492 42548 12498 42560
rect 12544 42557 12572 42588
rect 15105 42585 15117 42588
rect 15151 42585 15163 42619
rect 15105 42579 15163 42585
rect 15562 42576 15568 42628
rect 15620 42576 15626 42628
rect 16390 42576 16396 42628
rect 16448 42616 16454 42628
rect 16448 42588 17172 42616
rect 16448 42576 16454 42588
rect 12529 42551 12587 42557
rect 12529 42548 12541 42551
rect 12492 42520 12541 42548
rect 12492 42508 12498 42520
rect 12529 42517 12541 42520
rect 12575 42517 12587 42551
rect 12529 42511 12587 42517
rect 16577 42551 16635 42557
rect 16577 42517 16589 42551
rect 16623 42548 16635 42551
rect 16666 42548 16672 42560
rect 16623 42520 16672 42548
rect 16623 42517 16635 42520
rect 16577 42511 16635 42517
rect 16666 42508 16672 42520
rect 16724 42508 16730 42560
rect 17144 42557 17172 42588
rect 21174 42576 21180 42628
rect 21232 42616 21238 42628
rect 22189 42619 22247 42625
rect 22189 42616 22201 42619
rect 21232 42588 22201 42616
rect 21232 42576 21238 42588
rect 22189 42585 22201 42588
rect 22235 42585 22247 42619
rect 23216 42616 23244 42647
rect 23658 42644 23664 42656
rect 23716 42644 23722 42696
rect 23750 42644 23756 42696
rect 23808 42684 23814 42696
rect 24854 42684 24860 42696
rect 23808 42656 24860 42684
rect 23808 42644 23814 42656
rect 24854 42644 24860 42656
rect 24912 42644 24918 42696
rect 23216 42588 24532 42616
rect 22189 42579 22247 42585
rect 17129 42551 17187 42557
rect 17129 42517 17141 42551
rect 17175 42517 17187 42551
rect 17129 42511 17187 42517
rect 17497 42551 17555 42557
rect 17497 42517 17509 42551
rect 17543 42548 17555 42551
rect 19334 42548 19340 42560
rect 17543 42520 19340 42548
rect 17543 42517 17555 42520
rect 17497 42511 17555 42517
rect 19334 42508 19340 42520
rect 19392 42508 19398 42560
rect 20530 42508 20536 42560
rect 20588 42548 20594 42560
rect 21269 42551 21327 42557
rect 21269 42548 21281 42551
rect 20588 42520 21281 42548
rect 20588 42508 20594 42520
rect 21269 42517 21281 42520
rect 21315 42517 21327 42551
rect 21269 42511 21327 42517
rect 21821 42551 21879 42557
rect 21821 42517 21833 42551
rect 21867 42548 21879 42551
rect 22094 42548 22100 42560
rect 21867 42520 22100 42548
rect 21867 42517 21879 42520
rect 21821 42511 21879 42517
rect 22094 42508 22100 42520
rect 22152 42508 22158 42560
rect 24504 42557 24532 42588
rect 24489 42551 24547 42557
rect 24489 42517 24501 42551
rect 24535 42548 24547 42551
rect 24854 42548 24860 42560
rect 24535 42520 24860 42548
rect 24535 42517 24547 42520
rect 24489 42511 24547 42517
rect 24854 42508 24860 42520
rect 24912 42508 24918 42560
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 4154 42304 4160 42356
rect 4212 42344 4218 42356
rect 4341 42347 4399 42353
rect 4341 42344 4353 42347
rect 4212 42316 4353 42344
rect 4212 42304 4218 42316
rect 4341 42313 4353 42316
rect 4387 42313 4399 42347
rect 4341 42307 4399 42313
rect 5074 42304 5080 42356
rect 5132 42304 5138 42356
rect 5442 42304 5448 42356
rect 5500 42344 5506 42356
rect 6733 42347 6791 42353
rect 6733 42344 6745 42347
rect 5500 42316 6745 42344
rect 5500 42304 5506 42316
rect 6733 42313 6745 42316
rect 6779 42313 6791 42347
rect 8110 42344 8116 42356
rect 6733 42307 6791 42313
rect 7576 42316 8116 42344
rect 7576 42276 7604 42316
rect 8110 42304 8116 42316
rect 8168 42344 8174 42356
rect 9214 42344 9220 42356
rect 8168 42316 9220 42344
rect 8168 42304 8174 42316
rect 9214 42304 9220 42316
rect 9272 42304 9278 42356
rect 9674 42304 9680 42356
rect 9732 42304 9738 42356
rect 11422 42304 11428 42356
rect 11480 42344 11486 42356
rect 11793 42347 11851 42353
rect 11793 42344 11805 42347
rect 11480 42316 11805 42344
rect 11480 42304 11486 42316
rect 11793 42313 11805 42316
rect 11839 42313 11851 42347
rect 11793 42307 11851 42313
rect 12989 42347 13047 42353
rect 12989 42313 13001 42347
rect 13035 42344 13047 42347
rect 13446 42344 13452 42356
rect 13035 42316 13452 42344
rect 13035 42313 13047 42316
rect 12989 42307 13047 42313
rect 13446 42304 13452 42316
rect 13504 42304 13510 42356
rect 15194 42304 15200 42356
rect 15252 42344 15258 42356
rect 15381 42347 15439 42353
rect 15381 42344 15393 42347
rect 15252 42316 15393 42344
rect 15252 42304 15258 42316
rect 15381 42313 15393 42316
rect 15427 42313 15439 42347
rect 15381 42307 15439 42313
rect 15841 42347 15899 42353
rect 15841 42313 15853 42347
rect 15887 42344 15899 42347
rect 16853 42347 16911 42353
rect 16853 42344 16865 42347
rect 15887 42316 16865 42344
rect 15887 42313 15899 42316
rect 15841 42307 15899 42313
rect 16853 42313 16865 42316
rect 16899 42313 16911 42347
rect 16853 42307 16911 42313
rect 17221 42347 17279 42353
rect 17221 42313 17233 42347
rect 17267 42344 17279 42347
rect 18141 42347 18199 42353
rect 18141 42344 18153 42347
rect 17267 42316 18153 42344
rect 17267 42313 17279 42316
rect 17221 42307 17279 42313
rect 18141 42313 18153 42316
rect 18187 42344 18199 42347
rect 19794 42344 19800 42356
rect 18187 42316 19800 42344
rect 18187 42313 18199 42316
rect 18141 42307 18199 42313
rect 19794 42304 19800 42316
rect 19852 42344 19858 42356
rect 20162 42344 20168 42356
rect 19852 42316 20168 42344
rect 19852 42304 19858 42316
rect 20162 42304 20168 42316
rect 20220 42304 20226 42356
rect 20257 42347 20315 42353
rect 20257 42313 20269 42347
rect 20303 42313 20315 42347
rect 20257 42307 20315 42313
rect 7484 42248 7604 42276
rect 12253 42279 12311 42285
rect 3881 42211 3939 42217
rect 3881 42177 3893 42211
rect 3927 42208 3939 42211
rect 4246 42208 4252 42220
rect 3927 42180 4252 42208
rect 3927 42177 3939 42180
rect 3881 42171 3939 42177
rect 4246 42168 4252 42180
rect 4304 42168 4310 42220
rect 4985 42211 5043 42217
rect 4985 42177 4997 42211
rect 5031 42208 5043 42211
rect 6641 42211 6699 42217
rect 5031 42180 5580 42208
rect 5031 42177 5043 42180
rect 4985 42171 5043 42177
rect 5552 42013 5580 42180
rect 6641 42177 6653 42211
rect 6687 42208 6699 42211
rect 7006 42208 7012 42220
rect 6687 42180 7012 42208
rect 6687 42177 6699 42180
rect 6641 42171 6699 42177
rect 7006 42168 7012 42180
rect 7064 42168 7070 42220
rect 7484 42217 7512 42248
rect 12253 42245 12265 42279
rect 12299 42276 12311 42279
rect 15562 42276 15568 42288
rect 12299 42248 15568 42276
rect 12299 42245 12311 42248
rect 12253 42239 12311 42245
rect 15562 42236 15568 42248
rect 15620 42236 15626 42288
rect 15749 42279 15807 42285
rect 15749 42245 15761 42279
rect 15795 42276 15807 42279
rect 17862 42276 17868 42288
rect 15795 42248 17868 42276
rect 15795 42245 15807 42248
rect 15749 42239 15807 42245
rect 17862 42236 17868 42248
rect 17920 42236 17926 42288
rect 20272 42276 20300 42307
rect 20714 42304 20720 42356
rect 20772 42304 20778 42356
rect 21358 42304 21364 42356
rect 21416 42304 21422 42356
rect 23290 42304 23296 42356
rect 23348 42344 23354 42356
rect 25225 42347 25283 42353
rect 25225 42344 25237 42347
rect 23348 42316 25237 42344
rect 23348 42304 23354 42316
rect 25225 42313 25237 42316
rect 25271 42313 25283 42347
rect 25225 42307 25283 42313
rect 21082 42276 21088 42288
rect 20272 42248 21088 42276
rect 21082 42236 21088 42248
rect 21140 42236 21146 42288
rect 24302 42236 24308 42288
rect 24360 42236 24366 42288
rect 7469 42211 7527 42217
rect 7469 42177 7481 42211
rect 7515 42177 7527 42211
rect 7469 42171 7527 42177
rect 8846 42168 8852 42220
rect 8904 42168 8910 42220
rect 9122 42168 9128 42220
rect 9180 42208 9186 42220
rect 10045 42211 10103 42217
rect 9180 42180 9352 42208
rect 9180 42168 9186 42180
rect 7742 42100 7748 42152
rect 7800 42140 7806 42152
rect 9324 42140 9352 42180
rect 10045 42177 10057 42211
rect 10091 42177 10103 42211
rect 10045 42171 10103 42177
rect 10060 42140 10088 42171
rect 11146 42168 11152 42220
rect 11204 42208 11210 42220
rect 12161 42211 12219 42217
rect 12161 42208 12173 42211
rect 11204 42180 12173 42208
rect 11204 42168 11210 42180
rect 12161 42177 12173 42180
rect 12207 42177 12219 42211
rect 12161 42171 12219 42177
rect 13357 42211 13415 42217
rect 13357 42177 13369 42211
rect 13403 42208 13415 42211
rect 14185 42211 14243 42217
rect 14185 42208 14197 42211
rect 13403 42180 14197 42208
rect 13403 42177 13415 42180
rect 13357 42171 13415 42177
rect 14185 42177 14197 42180
rect 14231 42177 14243 42211
rect 14185 42171 14243 42177
rect 18877 42211 18935 42217
rect 18877 42177 18889 42211
rect 18923 42177 18935 42211
rect 18877 42171 18935 42177
rect 7800 42112 9260 42140
rect 9324 42112 10088 42140
rect 7800 42100 7806 42112
rect 9232 42072 9260 42112
rect 10134 42100 10140 42152
rect 10192 42100 10198 42152
rect 10229 42143 10287 42149
rect 10229 42109 10241 42143
rect 10275 42109 10287 42143
rect 10229 42103 10287 42109
rect 10244 42072 10272 42103
rect 12434 42100 12440 42152
rect 12492 42100 12498 42152
rect 13449 42143 13507 42149
rect 13449 42109 13461 42143
rect 13495 42109 13507 42143
rect 13449 42103 13507 42109
rect 13633 42143 13691 42149
rect 13633 42109 13645 42143
rect 13679 42140 13691 42143
rect 14274 42140 14280 42152
rect 13679 42112 14280 42140
rect 13679 42109 13691 42112
rect 13633 42103 13691 42109
rect 9232 42044 10272 42072
rect 13354 42032 13360 42084
rect 13412 42072 13418 42084
rect 13464 42072 13492 42103
rect 14274 42100 14280 42112
rect 14332 42140 14338 42152
rect 15933 42143 15991 42149
rect 15933 42140 15945 42143
rect 14332 42112 15945 42140
rect 14332 42100 14338 42112
rect 15933 42109 15945 42112
rect 15979 42109 15991 42143
rect 17313 42143 17371 42149
rect 17313 42140 17325 42143
rect 15933 42103 15991 42109
rect 16408 42112 17325 42140
rect 13412 42044 13492 42072
rect 13412 42032 13418 42044
rect 5537 42007 5595 42013
rect 5537 41973 5549 42007
rect 5583 42004 5595 42007
rect 6086 42004 6092 42016
rect 5583 41976 6092 42004
rect 5583 41973 5595 41976
rect 5537 41967 5595 41973
rect 6086 41964 6092 41976
rect 6144 41964 6150 42016
rect 7006 41964 7012 42016
rect 7064 42004 7070 42016
rect 7101 42007 7159 42013
rect 7101 42004 7113 42007
rect 7064 41976 7113 42004
rect 7064 41964 7070 41976
rect 7101 41973 7113 41976
rect 7147 41973 7159 42007
rect 7101 41967 7159 41973
rect 9217 42007 9275 42013
rect 9217 41973 9229 42007
rect 9263 42004 9275 42007
rect 9582 42004 9588 42016
rect 9263 41976 9588 42004
rect 9263 41973 9275 41976
rect 9217 41967 9275 41973
rect 9582 41964 9588 41976
rect 9640 41964 9646 42016
rect 10502 41964 10508 42016
rect 10560 42004 10566 42016
rect 10689 42007 10747 42013
rect 10689 42004 10701 42007
rect 10560 41976 10701 42004
rect 10560 41964 10566 41976
rect 10689 41973 10701 41976
rect 10735 41973 10747 42007
rect 10689 41967 10747 41973
rect 15102 41964 15108 42016
rect 15160 42004 15166 42016
rect 16408 42013 16436 42112
rect 17313 42109 17325 42112
rect 17359 42109 17371 42143
rect 17313 42103 17371 42109
rect 17497 42143 17555 42149
rect 17497 42109 17509 42143
rect 17543 42140 17555 42143
rect 17865 42143 17923 42149
rect 17865 42140 17877 42143
rect 17543 42112 17877 42140
rect 17543 42109 17555 42112
rect 17497 42103 17555 42109
rect 17865 42109 17877 42112
rect 17911 42109 17923 42143
rect 17865 42103 17923 42109
rect 16482 42032 16488 42084
rect 16540 42072 16546 42084
rect 17512 42072 17540 42103
rect 16540 42044 17540 42072
rect 18601 42075 18659 42081
rect 16540 42032 16546 42044
rect 18601 42041 18613 42075
rect 18647 42072 18659 42075
rect 18892 42072 18920 42171
rect 19518 42168 19524 42220
rect 19576 42208 19582 42220
rect 20625 42211 20683 42217
rect 20625 42208 20637 42211
rect 19576 42180 20637 42208
rect 19576 42168 19582 42180
rect 20625 42177 20637 42180
rect 20671 42177 20683 42211
rect 22005 42211 22063 42217
rect 22005 42208 22017 42211
rect 20625 42171 20683 42177
rect 21560 42180 22017 42208
rect 19242 42100 19248 42152
rect 19300 42140 19306 42152
rect 19613 42143 19671 42149
rect 19613 42140 19625 42143
rect 19300 42112 19625 42140
rect 19300 42100 19306 42112
rect 19613 42109 19625 42112
rect 19659 42109 19671 42143
rect 19613 42103 19671 42109
rect 19702 42100 19708 42152
rect 19760 42140 19766 42152
rect 20530 42140 20536 42152
rect 19760 42112 20536 42140
rect 19760 42100 19766 42112
rect 20530 42100 20536 42112
rect 20588 42140 20594 42152
rect 20809 42143 20867 42149
rect 20809 42140 20821 42143
rect 20588 42112 20821 42140
rect 20588 42100 20594 42112
rect 20809 42109 20821 42112
rect 20855 42109 20867 42143
rect 20809 42103 20867 42109
rect 21560 42081 21588 42180
rect 22005 42177 22017 42180
rect 22051 42177 22063 42211
rect 22005 42171 22063 42177
rect 22830 42100 22836 42152
rect 22888 42140 22894 42152
rect 23474 42140 23480 42152
rect 22888 42112 23480 42140
rect 22888 42100 22894 42112
rect 23474 42100 23480 42112
rect 23532 42100 23538 42152
rect 23753 42143 23811 42149
rect 23753 42109 23765 42143
rect 23799 42140 23811 42143
rect 25222 42140 25228 42152
rect 23799 42112 25228 42140
rect 23799 42109 23811 42112
rect 23753 42103 23811 42109
rect 25222 42100 25228 42112
rect 25280 42100 25286 42152
rect 21545 42075 21603 42081
rect 21545 42072 21557 42075
rect 18647 42044 21557 42072
rect 18647 42041 18659 42044
rect 18601 42035 18659 42041
rect 20732 42016 20760 42044
rect 21545 42041 21557 42044
rect 21591 42041 21603 42075
rect 21545 42035 21603 42041
rect 16393 42007 16451 42013
rect 16393 42004 16405 42007
rect 15160 41976 16405 42004
rect 15160 41964 15166 41976
rect 16393 41973 16405 41976
rect 16439 41973 16451 42007
rect 16393 41967 16451 41973
rect 20714 41964 20720 42016
rect 20772 41964 20778 42016
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 5166 41760 5172 41812
rect 5224 41760 5230 41812
rect 7653 41803 7711 41809
rect 7653 41769 7665 41803
rect 7699 41800 7711 41803
rect 7742 41800 7748 41812
rect 7699 41772 7748 41800
rect 7699 41769 7711 41772
rect 7653 41763 7711 41769
rect 7742 41760 7748 41772
rect 7800 41760 7806 41812
rect 7834 41760 7840 41812
rect 7892 41800 7898 41812
rect 8110 41800 8116 41812
rect 7892 41772 8116 41800
rect 7892 41760 7898 41772
rect 8110 41760 8116 41772
rect 8168 41760 8174 41812
rect 10689 41803 10747 41809
rect 10689 41769 10701 41803
rect 10735 41800 10747 41803
rect 11054 41800 11060 41812
rect 10735 41772 11060 41800
rect 10735 41769 10747 41772
rect 10689 41763 10747 41769
rect 11054 41760 11060 41772
rect 11112 41760 11118 41812
rect 20806 41760 20812 41812
rect 20864 41800 20870 41812
rect 21177 41803 21235 41809
rect 21177 41800 21189 41803
rect 20864 41772 21189 41800
rect 20864 41760 20870 41772
rect 21177 41769 21189 41772
rect 21223 41800 21235 41803
rect 21266 41800 21272 41812
rect 21223 41772 21272 41800
rect 21223 41769 21235 41772
rect 21177 41763 21235 41769
rect 21266 41760 21272 41772
rect 21324 41760 21330 41812
rect 21726 41760 21732 41812
rect 21784 41800 21790 41812
rect 25866 41800 25872 41812
rect 21784 41772 25872 41800
rect 21784 41760 21790 41772
rect 25866 41760 25872 41772
rect 25924 41760 25930 41812
rect 8021 41735 8079 41741
rect 8021 41701 8033 41735
rect 8067 41732 8079 41735
rect 8294 41732 8300 41744
rect 8067 41704 8300 41732
rect 8067 41701 8079 41704
rect 8021 41695 8079 41701
rect 5905 41667 5963 41673
rect 5905 41633 5917 41667
rect 5951 41664 5963 41667
rect 6178 41664 6184 41676
rect 5951 41636 6184 41664
rect 5951 41633 5963 41636
rect 5905 41627 5963 41633
rect 6178 41624 6184 41636
rect 6236 41624 6242 41676
rect 8036 41596 8064 41695
rect 8294 41692 8300 41704
rect 8352 41732 8358 41744
rect 8754 41732 8760 41744
rect 8352 41704 8760 41732
rect 8352 41692 8358 41704
rect 8754 41692 8760 41704
rect 8812 41692 8818 41744
rect 9674 41692 9680 41744
rect 9732 41732 9738 41744
rect 10870 41732 10876 41744
rect 9732 41704 10876 41732
rect 9732 41692 9738 41704
rect 10870 41692 10876 41704
rect 10928 41692 10934 41744
rect 17313 41735 17371 41741
rect 17313 41701 17325 41735
rect 17359 41732 17371 41735
rect 22833 41735 22891 41741
rect 17359 41704 19564 41732
rect 17359 41701 17371 41704
rect 17313 41695 17371 41701
rect 9214 41624 9220 41676
rect 9272 41664 9278 41676
rect 10045 41667 10103 41673
rect 10045 41664 10057 41667
rect 9272 41636 10057 41664
rect 9272 41624 9278 41636
rect 10045 41633 10057 41636
rect 10091 41664 10103 41667
rect 10594 41664 10600 41676
rect 10091 41636 10600 41664
rect 10091 41633 10103 41636
rect 10045 41627 10103 41633
rect 10594 41624 10600 41636
rect 10652 41624 10658 41676
rect 10778 41624 10784 41676
rect 10836 41664 10842 41676
rect 11241 41667 11299 41673
rect 11241 41664 11253 41667
rect 10836 41636 11253 41664
rect 10836 41624 10842 41636
rect 11241 41633 11253 41636
rect 11287 41633 11299 41667
rect 11241 41627 11299 41633
rect 12342 41624 12348 41676
rect 12400 41664 12406 41676
rect 12713 41667 12771 41673
rect 12713 41664 12725 41667
rect 12400 41636 12725 41664
rect 12400 41624 12406 41636
rect 12713 41633 12725 41636
rect 12759 41664 12771 41667
rect 12802 41664 12808 41676
rect 12759 41636 12808 41664
rect 12759 41633 12771 41636
rect 12713 41627 12771 41633
rect 12802 41624 12808 41636
rect 12860 41664 12866 41676
rect 13630 41664 13636 41676
rect 12860 41636 13636 41664
rect 12860 41624 12866 41636
rect 13630 41624 13636 41636
rect 13688 41624 13694 41676
rect 13906 41624 13912 41676
rect 13964 41664 13970 41676
rect 16114 41664 16120 41676
rect 13964 41636 16120 41664
rect 13964 41624 13970 41636
rect 16114 41624 16120 41636
rect 16172 41664 16178 41676
rect 16761 41667 16819 41673
rect 16761 41664 16773 41667
rect 16172 41636 16773 41664
rect 16172 41624 16178 41636
rect 16761 41633 16773 41636
rect 16807 41633 16819 41667
rect 16761 41627 16819 41633
rect 7314 41568 8064 41596
rect 9309 41599 9367 41605
rect 9309 41565 9321 41599
rect 9355 41596 9367 41599
rect 10502 41596 10508 41608
rect 9355 41568 10508 41596
rect 9355 41565 9367 41568
rect 9309 41559 9367 41565
rect 10502 41556 10508 41568
rect 10560 41596 10566 41608
rect 11977 41599 12035 41605
rect 11977 41596 11989 41599
rect 10560 41568 11989 41596
rect 10560 41556 10566 41568
rect 11977 41565 11989 41568
rect 12023 41596 12035 41599
rect 12023 41568 12434 41596
rect 12023 41565 12035 41568
rect 11977 41559 12035 41565
rect 5077 41531 5135 41537
rect 5077 41497 5089 41531
rect 5123 41497 5135 41531
rect 5077 41491 5135 41497
rect 6181 41531 6239 41537
rect 6181 41497 6193 41531
rect 6227 41497 6239 41531
rect 6181 41491 6239 41497
rect 1394 41420 1400 41472
rect 1452 41420 1458 41472
rect 5092 41460 5120 41491
rect 5629 41463 5687 41469
rect 5629 41460 5641 41463
rect 5092 41432 5641 41460
rect 5629 41429 5641 41432
rect 5675 41460 5687 41463
rect 5718 41460 5724 41472
rect 5675 41432 5724 41460
rect 5675 41429 5687 41432
rect 5629 41423 5687 41429
rect 5718 41420 5724 41432
rect 5776 41420 5782 41472
rect 6196 41460 6224 41491
rect 7742 41488 7748 41540
rect 7800 41528 7806 41540
rect 9122 41528 9128 41540
rect 7800 41500 9128 41528
rect 7800 41488 7806 41500
rect 9122 41488 9128 41500
rect 9180 41488 9186 41540
rect 12406 41528 12434 41568
rect 16574 41556 16580 41608
rect 16632 41596 16638 41608
rect 16669 41599 16727 41605
rect 16669 41596 16681 41599
rect 16632 41568 16681 41596
rect 16632 41556 16638 41568
rect 16669 41565 16681 41568
rect 16715 41565 16727 41599
rect 16669 41559 16727 41565
rect 13173 41531 13231 41537
rect 13173 41528 13185 41531
rect 12406 41500 13185 41528
rect 13173 41497 13185 41500
rect 13219 41497 13231 41531
rect 13173 41491 13231 41497
rect 7558 41460 7564 41472
rect 6196 41432 7564 41460
rect 7558 41420 7564 41432
rect 7616 41420 7622 41472
rect 8570 41420 8576 41472
rect 8628 41460 8634 41472
rect 9306 41460 9312 41472
rect 8628 41432 9312 41460
rect 8628 41420 8634 41432
rect 9306 41420 9312 41432
rect 9364 41420 9370 41472
rect 10778 41420 10784 41472
rect 10836 41460 10842 41472
rect 10962 41460 10968 41472
rect 10836 41432 10968 41460
rect 10836 41420 10842 41432
rect 10962 41420 10968 41432
rect 11020 41420 11026 41472
rect 11054 41420 11060 41472
rect 11112 41420 11118 41472
rect 11149 41463 11207 41469
rect 11149 41429 11161 41463
rect 11195 41460 11207 41463
rect 12342 41460 12348 41472
rect 11195 41432 12348 41460
rect 11195 41429 11207 41432
rect 11149 41423 11207 41429
rect 12342 41420 12348 41432
rect 12400 41420 12406 41472
rect 16206 41420 16212 41472
rect 16264 41420 16270 41472
rect 16577 41463 16635 41469
rect 16577 41429 16589 41463
rect 16623 41460 16635 41463
rect 17328 41460 17356 41695
rect 18506 41624 18512 41676
rect 18564 41664 18570 41676
rect 18601 41667 18659 41673
rect 18601 41664 18613 41667
rect 18564 41636 18613 41664
rect 18564 41624 18570 41636
rect 18601 41633 18613 41636
rect 18647 41633 18659 41667
rect 18601 41627 18659 41633
rect 18785 41667 18843 41673
rect 18785 41633 18797 41667
rect 18831 41664 18843 41667
rect 18966 41664 18972 41676
rect 18831 41636 18972 41664
rect 18831 41633 18843 41636
rect 18785 41627 18843 41633
rect 18966 41624 18972 41636
rect 19024 41624 19030 41676
rect 19242 41624 19248 41676
rect 19300 41664 19306 41676
rect 19429 41667 19487 41673
rect 19429 41664 19441 41667
rect 19300 41636 19441 41664
rect 19300 41624 19306 41636
rect 19429 41633 19441 41636
rect 19475 41633 19487 41667
rect 19536 41664 19564 41704
rect 22833 41701 22845 41735
rect 22879 41732 22891 41735
rect 25038 41732 25044 41744
rect 22879 41704 25044 41732
rect 22879 41701 22891 41704
rect 22833 41695 22891 41701
rect 25038 41692 25044 41704
rect 25096 41692 25102 41744
rect 22281 41667 22339 41673
rect 19536 41636 21128 41664
rect 19429 41627 19487 41633
rect 21100 41596 21128 41636
rect 22281 41633 22293 41667
rect 22327 41664 22339 41667
rect 22554 41664 22560 41676
rect 22327 41636 22560 41664
rect 22327 41633 22339 41636
rect 22281 41627 22339 41633
rect 22554 41624 22560 41636
rect 22612 41624 22618 41676
rect 22738 41624 22744 41676
rect 22796 41664 22802 41676
rect 23293 41667 23351 41673
rect 23293 41664 23305 41667
rect 22796 41636 23305 41664
rect 22796 41624 22802 41636
rect 23293 41633 23305 41636
rect 23339 41633 23351 41667
rect 23293 41627 23351 41633
rect 23385 41667 23443 41673
rect 23385 41633 23397 41667
rect 23431 41664 23443 41667
rect 23474 41664 23480 41676
rect 23431 41636 23480 41664
rect 23431 41633 23443 41636
rect 23385 41627 23443 41633
rect 23474 41624 23480 41636
rect 23532 41664 23538 41676
rect 23842 41664 23848 41676
rect 23532 41636 23848 41664
rect 23532 41624 23538 41636
rect 23842 41624 23848 41636
rect 23900 41624 23906 41676
rect 23750 41596 23756 41608
rect 21100 41568 23756 41596
rect 23750 41556 23756 41568
rect 23808 41556 23814 41608
rect 24489 41599 24547 41605
rect 24489 41565 24501 41599
rect 24535 41596 24547 41599
rect 25314 41596 25320 41608
rect 24535 41568 25320 41596
rect 24535 41565 24547 41568
rect 24489 41559 24547 41565
rect 25314 41556 25320 41568
rect 25372 41556 25378 41608
rect 19702 41488 19708 41540
rect 19760 41488 19766 41540
rect 21358 41528 21364 41540
rect 20930 41500 21364 41528
rect 21358 41488 21364 41500
rect 21416 41488 21422 41540
rect 21542 41488 21548 41540
rect 21600 41528 21606 41540
rect 22097 41531 22155 41537
rect 22097 41528 22109 41531
rect 21600 41500 22109 41528
rect 21600 41488 21606 41500
rect 22097 41497 22109 41500
rect 22143 41497 22155 41531
rect 22097 41491 22155 41497
rect 22278 41488 22284 41540
rect 22336 41528 22342 41540
rect 23201 41531 23259 41537
rect 23201 41528 23213 41531
rect 22336 41500 23213 41528
rect 22336 41488 22342 41500
rect 23201 41497 23213 41500
rect 23247 41497 23259 41531
rect 23201 41491 23259 41497
rect 24213 41531 24271 41537
rect 24213 41497 24225 41531
rect 24259 41528 24271 41531
rect 24259 41500 25360 41528
rect 24259 41497 24271 41500
rect 24213 41491 24271 41497
rect 25332 41472 25360 41500
rect 16623 41432 17356 41460
rect 18141 41463 18199 41469
rect 16623 41429 16635 41432
rect 16577 41423 16635 41429
rect 18141 41429 18153 41463
rect 18187 41460 18199 41463
rect 18414 41460 18420 41472
rect 18187 41432 18420 41460
rect 18187 41429 18199 41432
rect 18141 41423 18199 41429
rect 18414 41420 18420 41432
rect 18472 41420 18478 41472
rect 18509 41463 18567 41469
rect 18509 41429 18521 41463
rect 18555 41460 18567 41463
rect 19150 41460 19156 41472
rect 18555 41432 19156 41460
rect 18555 41429 18567 41432
rect 18509 41423 18567 41429
rect 19150 41420 19156 41432
rect 19208 41420 19214 41472
rect 21634 41420 21640 41472
rect 21692 41420 21698 41472
rect 22002 41420 22008 41472
rect 22060 41420 22066 41472
rect 23842 41420 23848 41472
rect 23900 41460 23906 41472
rect 24302 41460 24308 41472
rect 23900 41432 24308 41460
rect 23900 41420 23906 41432
rect 24302 41420 24308 41432
rect 24360 41460 24366 41472
rect 24581 41463 24639 41469
rect 24581 41460 24593 41463
rect 24360 41432 24593 41460
rect 24360 41420 24366 41432
rect 24581 41429 24593 41432
rect 24627 41429 24639 41463
rect 24581 41423 24639 41429
rect 24854 41420 24860 41472
rect 24912 41420 24918 41472
rect 25130 41420 25136 41472
rect 25188 41420 25194 41472
rect 25314 41420 25320 41472
rect 25372 41420 25378 41472
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 1946 41216 1952 41268
rect 2004 41256 2010 41268
rect 3329 41259 3387 41265
rect 3329 41256 3341 41259
rect 2004 41228 3341 41256
rect 2004 41216 2010 41228
rect 3329 41225 3341 41228
rect 3375 41225 3387 41259
rect 3329 41219 3387 41225
rect 6178 41216 6184 41268
rect 6236 41256 6242 41268
rect 7834 41256 7840 41268
rect 6236 41228 7840 41256
rect 6236 41216 6242 41228
rect 7834 41216 7840 41228
rect 7892 41256 7898 41268
rect 8021 41259 8079 41265
rect 8021 41256 8033 41259
rect 7892 41228 8033 41256
rect 7892 41216 7898 41228
rect 8021 41225 8033 41228
rect 8067 41225 8079 41259
rect 9398 41256 9404 41268
rect 8021 41219 8079 41225
rect 8956 41228 9404 41256
rect 1302 41080 1308 41132
rect 1360 41120 1366 41132
rect 1581 41123 1639 41129
rect 1581 41120 1593 41123
rect 1360 41092 1593 41120
rect 1360 41080 1366 41092
rect 1581 41089 1593 41092
rect 1627 41089 1639 41123
rect 1581 41083 1639 41089
rect 3237 41123 3295 41129
rect 3237 41089 3249 41123
rect 3283 41120 3295 41123
rect 3697 41123 3755 41129
rect 3697 41120 3709 41123
rect 3283 41092 3709 41120
rect 3283 41089 3295 41092
rect 3237 41083 3295 41089
rect 3697 41089 3709 41092
rect 3743 41120 3755 41123
rect 4614 41120 4620 41132
rect 3743 41092 4620 41120
rect 3743 41089 3755 41092
rect 3697 41083 3755 41089
rect 4614 41080 4620 41092
rect 4672 41080 4678 41132
rect 8956 41129 8984 41228
rect 9398 41216 9404 41228
rect 9456 41216 9462 41268
rect 10042 41256 10048 41268
rect 9600 41228 10048 41256
rect 9122 41148 9128 41200
rect 9180 41188 9186 41200
rect 9600 41188 9628 41228
rect 10042 41216 10048 41228
rect 10100 41256 10106 41268
rect 10965 41259 11023 41265
rect 10965 41256 10977 41259
rect 10100 41228 10977 41256
rect 10100 41216 10106 41228
rect 10965 41225 10977 41228
rect 11011 41256 11023 41259
rect 11514 41256 11520 41268
rect 11011 41228 11520 41256
rect 11011 41225 11023 41228
rect 10965 41219 11023 41225
rect 11514 41216 11520 41228
rect 11572 41216 11578 41268
rect 11698 41216 11704 41268
rect 11756 41216 11762 41268
rect 12161 41259 12219 41265
rect 12161 41225 12173 41259
rect 12207 41256 12219 41259
rect 14918 41256 14924 41268
rect 12207 41228 14924 41256
rect 12207 41225 12219 41228
rect 12161 41219 12219 41225
rect 14918 41216 14924 41228
rect 14976 41216 14982 41268
rect 15749 41259 15807 41265
rect 15749 41256 15761 41259
rect 15028 41228 15761 41256
rect 9180 41160 9706 41188
rect 9180 41148 9186 41160
rect 15028 41132 15056 41228
rect 15749 41225 15761 41228
rect 15795 41256 15807 41259
rect 15838 41256 15844 41268
rect 15795 41228 15844 41256
rect 15795 41225 15807 41228
rect 15749 41219 15807 41225
rect 15838 41216 15844 41228
rect 15896 41216 15902 41268
rect 19242 41256 19248 41268
rect 16868 41228 19248 41256
rect 8941 41123 8999 41129
rect 8941 41089 8953 41123
rect 8987 41089 8999 41123
rect 8941 41083 8999 41089
rect 10502 41080 10508 41132
rect 10560 41120 10566 41132
rect 12069 41123 12127 41129
rect 12069 41120 12081 41123
rect 10560 41092 12081 41120
rect 10560 41080 10566 41092
rect 12069 41089 12081 41092
rect 12115 41089 12127 41123
rect 12069 41083 12127 41089
rect 13630 41080 13636 41132
rect 13688 41080 13694 41132
rect 15010 41080 15016 41132
rect 15068 41080 15074 41132
rect 16868 41129 16896 41228
rect 19242 41216 19248 41228
rect 19300 41216 19306 41268
rect 19886 41216 19892 41268
rect 19944 41216 19950 41268
rect 22002 41216 22008 41268
rect 22060 41216 22066 41268
rect 23474 41216 23480 41268
rect 23532 41256 23538 41268
rect 24673 41259 24731 41265
rect 24673 41256 24685 41259
rect 23532 41228 24685 41256
rect 23532 41216 23538 41228
rect 24673 41225 24685 41228
rect 24719 41225 24731 41259
rect 24673 41219 24731 41225
rect 18874 41188 18880 41200
rect 18354 41160 18880 41188
rect 18874 41148 18880 41160
rect 18932 41148 18938 41200
rect 24486 41188 24492 41200
rect 24426 41160 24492 41188
rect 24486 41148 24492 41160
rect 24544 41148 24550 41200
rect 16853 41123 16911 41129
rect 16853 41089 16865 41123
rect 16899 41089 16911 41123
rect 16853 41083 16911 41089
rect 19797 41123 19855 41129
rect 19797 41089 19809 41123
rect 19843 41120 19855 41123
rect 20438 41120 20444 41132
rect 19843 41092 20444 41120
rect 19843 41089 19855 41092
rect 19797 41083 19855 41089
rect 20438 41080 20444 41092
rect 20496 41080 20502 41132
rect 20898 41080 20904 41132
rect 20956 41120 20962 41132
rect 21085 41123 21143 41129
rect 21085 41120 21097 41123
rect 20956 41092 21097 41120
rect 20956 41080 20962 41092
rect 21085 41089 21097 41092
rect 21131 41089 21143 41123
rect 21085 41083 21143 41089
rect 25314 41080 25320 41132
rect 25372 41080 25378 41132
rect 9217 41055 9275 41061
rect 9217 41021 9229 41055
rect 9263 41052 9275 41055
rect 10226 41052 10232 41064
rect 9263 41024 10232 41052
rect 9263 41021 9275 41024
rect 9217 41015 9275 41021
rect 10226 41012 10232 41024
rect 10284 41012 10290 41064
rect 12250 41012 12256 41064
rect 12308 41012 12314 41064
rect 13906 41012 13912 41064
rect 13964 41012 13970 41064
rect 16666 41012 16672 41064
rect 16724 41052 16730 41064
rect 17129 41055 17187 41061
rect 17129 41052 17141 41055
rect 16724 41024 17141 41052
rect 16724 41012 16730 41024
rect 17129 41021 17141 41024
rect 17175 41052 17187 41055
rect 17175 41024 18368 41052
rect 17175 41021 17187 41024
rect 17129 41015 17187 41021
rect 15378 40944 15384 40996
rect 15436 40984 15442 40996
rect 16390 40984 16396 40996
rect 15436 40956 16396 40984
rect 15436 40944 15442 40956
rect 16390 40944 16396 40956
rect 16448 40944 16454 40996
rect 18340 40984 18368 41024
rect 19978 41012 19984 41064
rect 20036 41012 20042 41064
rect 20990 41012 20996 41064
rect 21048 41052 21054 41064
rect 21177 41055 21235 41061
rect 21177 41052 21189 41055
rect 21048 41024 21189 41052
rect 21048 41012 21054 41024
rect 21177 41021 21189 41024
rect 21223 41021 21235 41055
rect 21177 41015 21235 41021
rect 21269 41055 21327 41061
rect 21269 41021 21281 41055
rect 21315 41021 21327 41055
rect 21269 41015 21327 41021
rect 21284 40984 21312 41015
rect 22462 41012 22468 41064
rect 22520 41052 22526 41064
rect 22646 41052 22652 41064
rect 22520 41024 22652 41052
rect 22520 41012 22526 41024
rect 22646 41012 22652 41024
rect 22704 41012 22710 41064
rect 22830 41012 22836 41064
rect 22888 41052 22894 41064
rect 22925 41055 22983 41061
rect 22925 41052 22937 41055
rect 22888 41024 22937 41052
rect 22888 41012 22894 41024
rect 22925 41021 22937 41024
rect 22971 41021 22983 41055
rect 23201 41055 23259 41061
rect 23201 41052 23213 41055
rect 22925 41015 22983 41021
rect 23032 41024 23213 41052
rect 18340 40956 21312 40984
rect 22186 40944 22192 40996
rect 22244 40984 22250 40996
rect 23032 40984 23060 41024
rect 23201 41021 23213 41024
rect 23247 41052 23259 41055
rect 24854 41052 24860 41064
rect 23247 41024 24860 41052
rect 23247 41021 23259 41024
rect 23201 41015 23259 41021
rect 24854 41012 24860 41024
rect 24912 41012 24918 41064
rect 25133 40987 25191 40993
rect 25133 40984 25145 40987
rect 22244 40956 23060 40984
rect 24228 40956 25145 40984
rect 22244 40944 22250 40956
rect 1762 40876 1768 40928
rect 1820 40916 1826 40928
rect 2225 40919 2283 40925
rect 2225 40916 2237 40919
rect 1820 40888 2237 40916
rect 1820 40876 1826 40888
rect 2225 40885 2237 40888
rect 2271 40885 2283 40919
rect 2225 40879 2283 40885
rect 8478 40876 8484 40928
rect 8536 40916 8542 40928
rect 9030 40916 9036 40928
rect 8536 40888 9036 40916
rect 8536 40876 8542 40888
rect 9030 40876 9036 40888
rect 9088 40876 9094 40928
rect 10318 40876 10324 40928
rect 10376 40916 10382 40928
rect 10686 40916 10692 40928
rect 10376 40888 10692 40916
rect 10376 40876 10382 40888
rect 10686 40876 10692 40888
rect 10744 40876 10750 40928
rect 18322 40876 18328 40928
rect 18380 40916 18386 40928
rect 18601 40919 18659 40925
rect 18601 40916 18613 40919
rect 18380 40888 18613 40916
rect 18380 40876 18386 40888
rect 18601 40885 18613 40888
rect 18647 40885 18659 40919
rect 18601 40879 18659 40885
rect 19150 40876 19156 40928
rect 19208 40876 19214 40928
rect 19426 40876 19432 40928
rect 19484 40876 19490 40928
rect 20717 40919 20775 40925
rect 20717 40885 20729 40919
rect 20763 40916 20775 40919
rect 20806 40916 20812 40928
rect 20763 40888 20812 40916
rect 20763 40885 20775 40888
rect 20717 40879 20775 40885
rect 20806 40876 20812 40888
rect 20864 40876 20870 40928
rect 20898 40876 20904 40928
rect 20956 40916 20962 40928
rect 24228 40916 24256 40956
rect 25133 40953 25145 40956
rect 25179 40953 25191 40987
rect 25133 40947 25191 40953
rect 20956 40888 24256 40916
rect 20956 40876 20962 40888
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 7558 40672 7564 40724
rect 7616 40712 7622 40724
rect 7929 40715 7987 40721
rect 7929 40712 7941 40715
rect 7616 40684 7941 40712
rect 7616 40672 7622 40684
rect 7929 40681 7941 40684
rect 7975 40681 7987 40715
rect 7929 40675 7987 40681
rect 8478 40672 8484 40724
rect 8536 40712 8542 40724
rect 9582 40712 9588 40724
rect 8536 40684 9588 40712
rect 8536 40672 8542 40684
rect 9582 40672 9588 40684
rect 9640 40672 9646 40724
rect 10594 40672 10600 40724
rect 10652 40672 10658 40724
rect 17678 40672 17684 40724
rect 17736 40712 17742 40724
rect 19978 40712 19984 40724
rect 17736 40684 19984 40712
rect 17736 40672 17742 40684
rect 19978 40672 19984 40684
rect 20036 40672 20042 40724
rect 20901 40715 20959 40721
rect 20901 40681 20913 40715
rect 20947 40712 20959 40715
rect 21174 40712 21180 40724
rect 20947 40684 21180 40712
rect 20947 40681 20959 40684
rect 20901 40675 20959 40681
rect 21174 40672 21180 40684
rect 21232 40672 21238 40724
rect 22189 40715 22247 40721
rect 22189 40712 22201 40715
rect 21468 40684 22201 40712
rect 7760 40616 11560 40644
rect 6457 40579 6515 40585
rect 6457 40545 6469 40579
rect 6503 40576 6515 40579
rect 6546 40576 6552 40588
rect 6503 40548 6552 40576
rect 6503 40545 6515 40548
rect 6457 40539 6515 40545
rect 6546 40536 6552 40548
rect 6604 40576 6610 40588
rect 7760 40576 7788 40616
rect 6604 40548 7788 40576
rect 6604 40536 6610 40548
rect 9398 40536 9404 40588
rect 9456 40576 9462 40588
rect 11532 40585 11560 40616
rect 14642 40604 14648 40656
rect 14700 40644 14706 40656
rect 18690 40644 18696 40656
rect 14700 40616 18696 40644
rect 14700 40604 14706 40616
rect 18690 40604 18696 40616
rect 18748 40644 18754 40656
rect 18748 40616 20116 40644
rect 18748 40604 18754 40616
rect 9769 40579 9827 40585
rect 9769 40576 9781 40579
rect 9456 40548 9781 40576
rect 9456 40536 9462 40548
rect 9769 40545 9781 40548
rect 9815 40576 9827 40579
rect 10229 40579 10287 40585
rect 10229 40576 10241 40579
rect 9815 40548 10241 40576
rect 9815 40545 9827 40548
rect 9769 40539 9827 40545
rect 10229 40545 10241 40548
rect 10275 40545 10287 40579
rect 10229 40539 10287 40545
rect 11517 40579 11575 40585
rect 11517 40545 11529 40579
rect 11563 40545 11575 40579
rect 11517 40539 11575 40545
rect 13265 40579 13323 40585
rect 13265 40545 13277 40579
rect 13311 40576 13323 40579
rect 13630 40576 13636 40588
rect 13311 40548 13636 40576
rect 13311 40545 13323 40548
rect 13265 40539 13323 40545
rect 13630 40536 13636 40548
rect 13688 40536 13694 40588
rect 13814 40536 13820 40588
rect 13872 40576 13878 40588
rect 13998 40576 14004 40588
rect 13872 40548 14004 40576
rect 13872 40536 13878 40548
rect 13998 40536 14004 40548
rect 14056 40576 14062 40588
rect 14737 40579 14795 40585
rect 14737 40576 14749 40579
rect 14056 40548 14749 40576
rect 14056 40536 14062 40548
rect 14737 40545 14749 40548
rect 14783 40576 14795 40579
rect 15841 40579 15899 40585
rect 15841 40576 15853 40579
rect 14783 40548 15853 40576
rect 14783 40545 14795 40548
rect 14737 40539 14795 40545
rect 15841 40545 15853 40548
rect 15887 40576 15899 40579
rect 16942 40576 16948 40588
rect 15887 40548 16948 40576
rect 15887 40545 15899 40548
rect 15841 40539 15899 40545
rect 16942 40536 16948 40548
rect 17000 40536 17006 40588
rect 17034 40536 17040 40588
rect 17092 40576 17098 40588
rect 17129 40579 17187 40585
rect 17129 40576 17141 40579
rect 17092 40548 17141 40576
rect 17092 40536 17098 40548
rect 17129 40545 17141 40548
rect 17175 40545 17187 40579
rect 17129 40539 17187 40545
rect 17218 40536 17224 40588
rect 17276 40536 17282 40588
rect 1762 40468 1768 40520
rect 1820 40468 1826 40520
rect 6178 40468 6184 40520
rect 6236 40468 6242 40520
rect 8757 40511 8815 40517
rect 1581 40375 1639 40381
rect 1581 40341 1593 40375
rect 1627 40372 1639 40375
rect 1854 40372 1860 40384
rect 1627 40344 1860 40372
rect 1627 40341 1639 40344
rect 1581 40335 1639 40341
rect 1854 40332 1860 40344
rect 1912 40332 1918 40384
rect 7282 40332 7288 40384
rect 7340 40372 7346 40384
rect 7576 40372 7604 40494
rect 8757 40477 8769 40511
rect 8803 40508 8815 40511
rect 9214 40508 9220 40520
rect 8803 40480 9220 40508
rect 8803 40477 8815 40480
rect 8757 40471 8815 40477
rect 9214 40468 9220 40480
rect 9272 40508 9278 40520
rect 9677 40511 9735 40517
rect 9677 40508 9689 40511
rect 9272 40480 9689 40508
rect 9272 40468 9278 40480
rect 9677 40477 9689 40480
rect 9723 40508 9735 40511
rect 11882 40508 11888 40520
rect 9723 40480 11888 40508
rect 9723 40477 9735 40480
rect 9677 40471 9735 40477
rect 11882 40468 11888 40480
rect 11940 40468 11946 40520
rect 11974 40468 11980 40520
rect 12032 40508 12038 40520
rect 12032 40480 12434 40508
rect 12032 40468 12038 40480
rect 9490 40400 9496 40452
rect 9548 40440 9554 40452
rect 11057 40443 11115 40449
rect 11057 40440 11069 40443
rect 9548 40412 11069 40440
rect 9548 40400 9554 40412
rect 11057 40409 11069 40412
rect 11103 40409 11115 40443
rect 11057 40403 11115 40409
rect 11333 40443 11391 40449
rect 11333 40409 11345 40443
rect 11379 40440 11391 40443
rect 11793 40443 11851 40449
rect 11793 40440 11805 40443
rect 11379 40412 11805 40440
rect 11379 40409 11391 40412
rect 11333 40403 11391 40409
rect 11793 40409 11805 40412
rect 11839 40440 11851 40443
rect 12250 40440 12256 40452
rect 11839 40412 12256 40440
rect 11839 40409 11851 40412
rect 11793 40403 11851 40409
rect 8294 40372 8300 40384
rect 7340 40344 8300 40372
rect 7340 40332 7346 40344
rect 8294 40332 8300 40344
rect 8352 40372 8358 40384
rect 9122 40372 9128 40384
rect 8352 40344 9128 40372
rect 8352 40332 8358 40344
rect 9122 40332 9128 40344
rect 9180 40332 9186 40384
rect 9214 40332 9220 40384
rect 9272 40332 9278 40384
rect 9582 40332 9588 40384
rect 9640 40332 9646 40384
rect 11072 40372 11100 40403
rect 12250 40400 12256 40412
rect 12308 40400 12314 40452
rect 12406 40440 12434 40480
rect 12710 40468 12716 40520
rect 12768 40508 12774 40520
rect 12989 40511 13047 40517
rect 12989 40508 13001 40511
rect 12768 40480 13001 40508
rect 12768 40468 12774 40480
rect 12989 40477 13001 40480
rect 13035 40477 13047 40511
rect 12989 40471 13047 40477
rect 13081 40511 13139 40517
rect 13081 40477 13093 40511
rect 13127 40508 13139 40511
rect 13725 40511 13783 40517
rect 13725 40508 13737 40511
rect 13127 40480 13737 40508
rect 13127 40477 13139 40480
rect 13081 40471 13139 40477
rect 13725 40477 13737 40480
rect 13771 40508 13783 40511
rect 16850 40508 16856 40520
rect 13771 40480 16856 40508
rect 13771 40477 13783 40480
rect 13725 40471 13783 40477
rect 16850 40468 16856 40480
rect 16908 40468 16914 40520
rect 19334 40468 19340 40520
rect 19392 40508 19398 40520
rect 19978 40508 19984 40520
rect 19392 40480 19984 40508
rect 19392 40468 19398 40480
rect 19978 40468 19984 40480
rect 20036 40468 20042 40520
rect 20088 40508 20116 40616
rect 21174 40508 21180 40520
rect 20088 40480 21180 40508
rect 21174 40468 21180 40480
rect 21232 40468 21238 40520
rect 21269 40511 21327 40517
rect 21269 40477 21281 40511
rect 21315 40508 21327 40511
rect 21468 40508 21496 40684
rect 22189 40681 22201 40684
rect 22235 40712 22247 40715
rect 22738 40712 22744 40724
rect 22235 40684 22744 40712
rect 22235 40681 22247 40684
rect 22189 40675 22247 40681
rect 22738 40672 22744 40684
rect 22796 40712 22802 40724
rect 25774 40712 25780 40724
rect 22796 40684 25780 40712
rect 22796 40672 22802 40684
rect 25774 40672 25780 40684
rect 25832 40672 25838 40724
rect 21542 40536 21548 40588
rect 21600 40536 21606 40588
rect 21726 40536 21732 40588
rect 21784 40576 21790 40588
rect 21913 40579 21971 40585
rect 21913 40576 21925 40579
rect 21784 40548 21925 40576
rect 21784 40536 21790 40548
rect 21913 40545 21925 40548
rect 21959 40545 21971 40579
rect 21913 40539 21971 40545
rect 22094 40536 22100 40588
rect 22152 40576 22158 40588
rect 22925 40579 22983 40585
rect 22925 40576 22937 40579
rect 22152 40548 22937 40576
rect 22152 40536 22158 40548
rect 22925 40545 22937 40548
rect 22971 40545 22983 40579
rect 22925 40539 22983 40545
rect 23109 40579 23167 40585
rect 23109 40545 23121 40579
rect 23155 40576 23167 40579
rect 23382 40576 23388 40588
rect 23155 40548 23388 40576
rect 23155 40545 23167 40548
rect 23109 40539 23167 40545
rect 23382 40536 23388 40548
rect 23440 40536 23446 40588
rect 21315 40480 21496 40508
rect 21315 40477 21327 40480
rect 21269 40471 21327 40477
rect 21634 40468 21640 40520
rect 21692 40508 21698 40520
rect 22833 40511 22891 40517
rect 22833 40508 22845 40511
rect 21692 40480 22845 40508
rect 21692 40468 21698 40480
rect 22833 40477 22845 40480
rect 22879 40477 22891 40511
rect 22833 40471 22891 40477
rect 23014 40468 23020 40520
rect 23072 40508 23078 40520
rect 24394 40508 24400 40520
rect 23072 40480 24400 40508
rect 23072 40468 23078 40480
rect 24394 40468 24400 40480
rect 24452 40468 24458 40520
rect 24673 40511 24731 40517
rect 24673 40477 24685 40511
rect 24719 40508 24731 40511
rect 24762 40508 24768 40520
rect 24719 40480 24768 40508
rect 24719 40477 24731 40480
rect 24673 40471 24731 40477
rect 24762 40468 24768 40480
rect 24820 40508 24826 40520
rect 25317 40511 25375 40517
rect 25317 40508 25329 40511
rect 24820 40480 25329 40508
rect 24820 40468 24826 40480
rect 25317 40477 25329 40480
rect 25363 40477 25375 40511
rect 25317 40471 25375 40477
rect 14829 40443 14887 40449
rect 14829 40440 14841 40443
rect 12406 40412 14841 40440
rect 14829 40409 14841 40412
rect 14875 40440 14887 40443
rect 15657 40443 15715 40449
rect 15657 40440 15669 40443
rect 14875 40412 15669 40440
rect 14875 40409 14887 40412
rect 14829 40403 14887 40409
rect 15657 40409 15669 40412
rect 15703 40409 15715 40443
rect 15657 40403 15715 40409
rect 15838 40400 15844 40452
rect 15896 40440 15902 40452
rect 17037 40443 17095 40449
rect 17037 40440 17049 40443
rect 15896 40412 17049 40440
rect 15896 40400 15902 40412
rect 17037 40409 17049 40412
rect 17083 40409 17095 40443
rect 17037 40403 17095 40409
rect 19150 40400 19156 40452
rect 19208 40440 19214 40452
rect 19208 40412 21404 40440
rect 19208 40400 19214 40412
rect 11701 40375 11759 40381
rect 11701 40372 11713 40375
rect 11072 40344 11713 40372
rect 11701 40341 11713 40344
rect 11747 40341 11759 40375
rect 11701 40335 11759 40341
rect 12158 40332 12164 40384
rect 12216 40332 12222 40384
rect 12618 40332 12624 40384
rect 12676 40332 12682 40384
rect 15194 40332 15200 40384
rect 15252 40332 15258 40384
rect 15565 40375 15623 40381
rect 15565 40341 15577 40375
rect 15611 40372 15623 40375
rect 16298 40372 16304 40384
rect 15611 40344 16304 40372
rect 15611 40341 15623 40344
rect 15565 40335 15623 40341
rect 16298 40332 16304 40344
rect 16356 40332 16362 40384
rect 16669 40375 16727 40381
rect 16669 40341 16681 40375
rect 16715 40372 16727 40375
rect 17494 40372 17500 40384
rect 16715 40344 17500 40372
rect 16715 40341 16727 40344
rect 16669 40335 16727 40341
rect 17494 40332 17500 40344
rect 17552 40332 17558 40384
rect 20349 40375 20407 40381
rect 20349 40341 20361 40375
rect 20395 40372 20407 40375
rect 20438 40372 20444 40384
rect 20395 40344 20444 40372
rect 20395 40341 20407 40344
rect 20349 40335 20407 40341
rect 20438 40332 20444 40344
rect 20496 40332 20502 40384
rect 21376 40381 21404 40412
rect 21542 40400 21548 40452
rect 21600 40440 21606 40452
rect 22370 40440 22376 40452
rect 21600 40412 22376 40440
rect 21600 40400 21606 40412
rect 22370 40400 22376 40412
rect 22428 40440 22434 40452
rect 23750 40440 23756 40452
rect 22428 40412 23756 40440
rect 22428 40400 22434 40412
rect 23750 40400 23756 40412
rect 23808 40400 23814 40452
rect 24029 40443 24087 40449
rect 24029 40409 24041 40443
rect 24075 40440 24087 40443
rect 24857 40443 24915 40449
rect 24075 40412 24532 40440
rect 24075 40409 24087 40412
rect 24029 40403 24087 40409
rect 24504 40384 24532 40412
rect 24857 40409 24869 40443
rect 24903 40440 24915 40443
rect 24903 40412 25360 40440
rect 24903 40409 24915 40412
rect 24857 40403 24915 40409
rect 25332 40384 25360 40412
rect 21361 40375 21419 40381
rect 21361 40341 21373 40375
rect 21407 40372 21419 40375
rect 21726 40372 21732 40384
rect 21407 40344 21732 40372
rect 21407 40341 21419 40344
rect 21361 40335 21419 40341
rect 21726 40332 21732 40344
rect 21784 40332 21790 40384
rect 22465 40375 22523 40381
rect 22465 40341 22477 40375
rect 22511 40372 22523 40375
rect 23382 40372 23388 40384
rect 22511 40344 23388 40372
rect 22511 40341 22523 40344
rect 22465 40335 22523 40341
rect 23382 40332 23388 40344
rect 23440 40332 23446 40384
rect 24210 40332 24216 40384
rect 24268 40332 24274 40384
rect 24486 40332 24492 40384
rect 24544 40332 24550 40384
rect 24578 40332 24584 40384
rect 24636 40372 24642 40384
rect 25133 40375 25191 40381
rect 25133 40372 25145 40375
rect 24636 40344 25145 40372
rect 24636 40332 24642 40344
rect 25133 40341 25145 40344
rect 25179 40341 25191 40375
rect 25133 40335 25191 40341
rect 25314 40332 25320 40384
rect 25372 40332 25378 40384
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 7190 40128 7196 40180
rect 7248 40168 7254 40180
rect 7285 40171 7343 40177
rect 7285 40168 7297 40171
rect 7248 40140 7297 40168
rect 7248 40128 7254 40140
rect 7285 40137 7297 40140
rect 7331 40137 7343 40171
rect 7285 40131 7343 40137
rect 9122 40128 9128 40180
rect 9180 40128 9186 40180
rect 9398 40128 9404 40180
rect 9456 40168 9462 40180
rect 9456 40140 10548 40168
rect 9456 40128 9462 40140
rect 7653 40103 7711 40109
rect 7653 40069 7665 40103
rect 7699 40100 7711 40103
rect 8754 40100 8760 40112
rect 7699 40072 8760 40100
rect 7699 40069 7711 40072
rect 7653 40063 7711 40069
rect 8754 40060 8760 40072
rect 8812 40060 8818 40112
rect 9140 40100 9168 40128
rect 10520 40109 10548 40140
rect 11514 40128 11520 40180
rect 11572 40128 11578 40180
rect 12250 40128 12256 40180
rect 12308 40168 12314 40180
rect 14642 40168 14648 40180
rect 12308 40140 14648 40168
rect 12308 40128 12314 40140
rect 14642 40128 14648 40140
rect 14700 40128 14706 40180
rect 15010 40128 15016 40180
rect 15068 40128 15074 40180
rect 15562 40128 15568 40180
rect 15620 40128 15626 40180
rect 16298 40128 16304 40180
rect 16356 40168 16362 40180
rect 22094 40168 22100 40180
rect 16356 40140 22100 40168
rect 16356 40128 16362 40140
rect 22094 40128 22100 40140
rect 22152 40168 22158 40180
rect 22646 40168 22652 40180
rect 22152 40140 22652 40168
rect 22152 40128 22158 40140
rect 22646 40128 22652 40140
rect 22704 40128 22710 40180
rect 23658 40168 23664 40180
rect 22756 40140 23664 40168
rect 10505 40103 10563 40109
rect 9140 40072 9246 40100
rect 10505 40069 10517 40103
rect 10551 40069 10563 40103
rect 14550 40100 14556 40112
rect 14398 40072 14556 40100
rect 10505 40063 10563 40069
rect 14550 40060 14556 40072
rect 14608 40100 14614 40112
rect 15028 40100 15056 40128
rect 14608 40072 15056 40100
rect 15933 40103 15991 40109
rect 14608 40060 14614 40072
rect 15933 40069 15945 40103
rect 15979 40069 15991 40103
rect 15933 40063 15991 40069
rect 7926 39992 7932 40044
rect 7984 40032 7990 40044
rect 8481 40035 8539 40041
rect 8481 40032 8493 40035
rect 7984 40004 8493 40032
rect 7984 39992 7990 40004
rect 8481 40001 8493 40004
rect 8527 40001 8539 40035
rect 8481 39995 8539 40001
rect 12434 39992 12440 40044
rect 12492 40032 12498 40044
rect 12802 40032 12808 40044
rect 12492 40004 12808 40032
rect 12492 39992 12498 40004
rect 12802 39992 12808 40004
rect 12860 40032 12866 40044
rect 12897 40035 12955 40041
rect 12897 40032 12909 40035
rect 12860 40004 12909 40032
rect 12860 39992 12866 40004
rect 12897 40001 12909 40004
rect 12943 40001 12955 40035
rect 15948 40032 15976 40063
rect 18598 40060 18604 40112
rect 18656 40060 18662 40112
rect 20165 40103 20223 40109
rect 20165 40100 20177 40103
rect 19306 40072 20177 40100
rect 16298 40032 16304 40044
rect 15948 40004 16304 40032
rect 12897 39995 12955 40001
rect 16298 39992 16304 40004
rect 16356 39992 16362 40044
rect 7745 39967 7803 39973
rect 7745 39933 7757 39967
rect 7791 39933 7803 39967
rect 7745 39927 7803 39933
rect 7760 39896 7788 39927
rect 7834 39924 7840 39976
rect 7892 39924 7898 39976
rect 8757 39967 8815 39973
rect 8757 39933 8769 39967
rect 8803 39964 8815 39967
rect 10318 39964 10324 39976
rect 8803 39936 10324 39964
rect 8803 39933 8815 39936
rect 8757 39927 8815 39933
rect 10318 39924 10324 39936
rect 10376 39924 10382 39976
rect 10962 39924 10968 39976
rect 11020 39924 11026 39976
rect 13173 39967 13231 39973
rect 13173 39933 13185 39967
rect 13219 39964 13231 39967
rect 15378 39964 15384 39976
rect 13219 39936 15384 39964
rect 13219 39933 13231 39936
rect 13173 39927 13231 39933
rect 15378 39924 15384 39936
rect 15436 39924 15442 39976
rect 16022 39924 16028 39976
rect 16080 39924 16086 39976
rect 16117 39967 16175 39973
rect 16117 39933 16129 39967
rect 16163 39933 16175 39967
rect 16117 39927 16175 39933
rect 8478 39896 8484 39908
rect 7760 39868 8484 39896
rect 8478 39856 8484 39868
rect 8536 39856 8542 39908
rect 16132 39896 16160 39927
rect 18414 39924 18420 39976
rect 18472 39964 18478 39976
rect 18693 39967 18751 39973
rect 18693 39964 18705 39967
rect 18472 39936 18705 39964
rect 18472 39924 18478 39936
rect 18693 39933 18705 39936
rect 18739 39933 18751 39967
rect 18693 39927 18751 39933
rect 18782 39924 18788 39976
rect 18840 39924 18846 39976
rect 19306 39964 19334 40072
rect 20165 40069 20177 40072
rect 20211 40100 20223 40103
rect 20211 40072 21128 40100
rect 20211 40069 20223 40072
rect 20165 40063 20223 40069
rect 20254 39992 20260 40044
rect 20312 39992 20318 40044
rect 21100 40041 21128 40072
rect 21174 40060 21180 40112
rect 21232 40100 21238 40112
rect 22756 40100 22784 40140
rect 23658 40128 23664 40140
rect 23716 40128 23722 40180
rect 23750 40128 23756 40180
rect 23808 40168 23814 40180
rect 25225 40171 25283 40177
rect 25225 40168 25237 40171
rect 23808 40140 25237 40168
rect 23808 40128 23814 40140
rect 25225 40137 25237 40140
rect 25271 40137 25283 40171
rect 25225 40131 25283 40137
rect 21232 40072 22784 40100
rect 21232 40060 21238 40072
rect 22830 40060 22836 40112
rect 22888 40100 22894 40112
rect 22888 40072 23428 40100
rect 22888 40060 22894 40072
rect 21085 40035 21143 40041
rect 21085 40001 21097 40035
rect 21131 40032 21143 40035
rect 21358 40032 21364 40044
rect 21131 40004 21364 40032
rect 21131 40001 21143 40004
rect 21085 39995 21143 40001
rect 21358 39992 21364 40004
rect 21416 39992 21422 40044
rect 21726 39992 21732 40044
rect 21784 40032 21790 40044
rect 22281 40035 22339 40041
rect 22281 40032 22293 40035
rect 21784 40004 22293 40032
rect 21784 39992 21790 40004
rect 22281 40001 22293 40004
rect 22327 40001 22339 40035
rect 22281 39995 22339 40001
rect 22557 40035 22615 40041
rect 22557 40001 22569 40035
rect 22603 40032 22615 40035
rect 22738 40032 22744 40044
rect 22603 40004 22744 40032
rect 22603 40001 22615 40004
rect 22557 39995 22615 40001
rect 22738 39992 22744 40004
rect 22796 39992 22802 40044
rect 23400 40032 23428 40072
rect 24486 40060 24492 40112
rect 24544 40060 24550 40112
rect 23477 40035 23535 40041
rect 23477 40032 23489 40035
rect 23400 40004 23489 40032
rect 23477 40001 23489 40004
rect 23523 40001 23535 40035
rect 23477 39995 23535 40001
rect 18984 39936 19334 39964
rect 14200 39868 16160 39896
rect 13722 39788 13728 39840
rect 13780 39828 13786 39840
rect 14200 39828 14228 39868
rect 18230 39856 18236 39908
rect 18288 39856 18294 39908
rect 13780 39800 14228 39828
rect 13780 39788 13786 39800
rect 14642 39788 14648 39840
rect 14700 39828 14706 39840
rect 14826 39828 14832 39840
rect 14700 39800 14832 39828
rect 14700 39788 14706 39800
rect 14826 39788 14832 39800
rect 14884 39788 14890 39840
rect 16298 39788 16304 39840
rect 16356 39828 16362 39840
rect 16669 39831 16727 39837
rect 16669 39828 16681 39831
rect 16356 39800 16681 39828
rect 16356 39788 16362 39800
rect 16669 39797 16681 39800
rect 16715 39797 16727 39831
rect 16669 39791 16727 39797
rect 17126 39788 17132 39840
rect 17184 39828 17190 39840
rect 18984 39828 19012 39936
rect 20438 39924 20444 39976
rect 20496 39924 20502 39976
rect 20530 39924 20536 39976
rect 20588 39964 20594 39976
rect 21542 39964 21548 39976
rect 20588 39936 21548 39964
rect 20588 39924 20594 39936
rect 21542 39924 21548 39936
rect 21600 39924 21606 39976
rect 22646 39924 22652 39976
rect 22704 39964 22710 39976
rect 23014 39964 23020 39976
rect 22704 39936 23020 39964
rect 22704 39924 22710 39936
rect 23014 39924 23020 39936
rect 23072 39924 23078 39976
rect 23753 39967 23811 39973
rect 23753 39933 23765 39967
rect 23799 39964 23811 39967
rect 24486 39964 24492 39976
rect 23799 39936 24492 39964
rect 23799 39933 23811 39936
rect 23753 39927 23811 39933
rect 24486 39924 24492 39936
rect 24544 39924 24550 39976
rect 19518 39856 19524 39908
rect 19576 39896 19582 39908
rect 19797 39899 19855 39905
rect 19797 39896 19809 39899
rect 19576 39868 19809 39896
rect 19576 39856 19582 39868
rect 19797 39865 19809 39868
rect 19843 39865 19855 39899
rect 21818 39896 21824 39908
rect 19797 39859 19855 39865
rect 20180 39868 21824 39896
rect 17184 39800 19012 39828
rect 17184 39788 17190 39800
rect 19058 39788 19064 39840
rect 19116 39828 19122 39840
rect 20180 39828 20208 39868
rect 21818 39856 21824 39868
rect 21876 39856 21882 39908
rect 19116 39800 20208 39828
rect 19116 39788 19122 39800
rect 20254 39788 20260 39840
rect 20312 39828 20318 39840
rect 20901 39831 20959 39837
rect 20901 39828 20913 39831
rect 20312 39800 20913 39828
rect 20312 39788 20318 39800
rect 20901 39797 20913 39800
rect 20947 39828 20959 39831
rect 23750 39828 23756 39840
rect 20947 39800 23756 39828
rect 20947 39797 20959 39800
rect 20901 39791 20959 39797
rect 23750 39788 23756 39800
rect 23808 39788 23814 39840
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 6546 39584 6552 39636
rect 6604 39624 6610 39636
rect 6641 39627 6699 39633
rect 6641 39624 6653 39627
rect 6604 39596 6653 39624
rect 6604 39584 6610 39596
rect 6641 39593 6653 39596
rect 6687 39593 6699 39627
rect 6641 39587 6699 39593
rect 8478 39584 8484 39636
rect 8536 39624 8542 39636
rect 9769 39627 9827 39633
rect 9769 39624 9781 39627
rect 8536 39596 9781 39624
rect 8536 39584 8542 39596
rect 9769 39593 9781 39596
rect 9815 39593 9827 39627
rect 9769 39587 9827 39593
rect 11228 39627 11286 39633
rect 11228 39593 11240 39627
rect 11274 39624 11286 39627
rect 12250 39624 12256 39636
rect 11274 39596 12256 39624
rect 11274 39593 11286 39596
rect 11228 39587 11286 39593
rect 12250 39584 12256 39596
rect 12308 39624 12314 39636
rect 12308 39596 12940 39624
rect 12308 39584 12314 39596
rect 12713 39559 12771 39565
rect 12713 39525 12725 39559
rect 12759 39556 12771 39559
rect 12912 39556 12940 39596
rect 13078 39584 13084 39636
rect 13136 39624 13142 39636
rect 14274 39624 14280 39636
rect 13136 39596 14280 39624
rect 13136 39584 13142 39596
rect 14274 39584 14280 39596
rect 14332 39624 14338 39636
rect 14550 39624 14556 39636
rect 14332 39596 14556 39624
rect 14332 39584 14338 39596
rect 14550 39584 14556 39596
rect 14608 39584 14614 39636
rect 14734 39584 14740 39636
rect 14792 39624 14798 39636
rect 15565 39627 15623 39633
rect 15565 39624 15577 39627
rect 14792 39596 15577 39624
rect 14792 39584 14798 39596
rect 15565 39593 15577 39596
rect 15611 39593 15623 39627
rect 15565 39587 15623 39593
rect 18506 39584 18512 39636
rect 18564 39624 18570 39636
rect 18785 39627 18843 39633
rect 18785 39624 18797 39627
rect 18564 39596 18797 39624
rect 18564 39584 18570 39596
rect 18785 39593 18797 39596
rect 18831 39593 18843 39627
rect 18785 39587 18843 39593
rect 19058 39584 19064 39636
rect 19116 39584 19122 39636
rect 19610 39584 19616 39636
rect 19668 39624 19674 39636
rect 20438 39624 20444 39636
rect 19668 39596 20444 39624
rect 19668 39584 19674 39596
rect 20438 39584 20444 39596
rect 20496 39584 20502 39636
rect 21269 39627 21327 39633
rect 21269 39593 21281 39627
rect 21315 39624 21327 39627
rect 22278 39624 22284 39636
rect 21315 39596 22284 39624
rect 21315 39593 21327 39596
rect 21269 39587 21327 39593
rect 22278 39584 22284 39596
rect 22336 39584 22342 39636
rect 13265 39559 13323 39565
rect 13265 39556 13277 39559
rect 12759 39528 12848 39556
rect 12912 39528 13277 39556
rect 12759 39525 12771 39528
rect 12713 39519 12771 39525
rect 4893 39491 4951 39497
rect 4893 39457 4905 39491
rect 4939 39488 4951 39491
rect 6178 39488 6184 39500
rect 4939 39460 6184 39488
rect 4939 39457 4951 39460
rect 4893 39451 4951 39457
rect 6178 39448 6184 39460
rect 6236 39488 6242 39500
rect 7101 39491 7159 39497
rect 7101 39488 7113 39491
rect 6236 39460 7113 39488
rect 6236 39448 6242 39460
rect 7101 39457 7113 39460
rect 7147 39457 7159 39491
rect 7101 39451 7159 39457
rect 9214 39448 9220 39500
rect 9272 39488 9278 39500
rect 10229 39491 10287 39497
rect 10229 39488 10241 39491
rect 9272 39460 10241 39488
rect 9272 39448 9278 39460
rect 10229 39457 10241 39460
rect 10275 39457 10287 39491
rect 10229 39451 10287 39457
rect 10318 39448 10324 39500
rect 10376 39448 10382 39500
rect 10965 39491 11023 39497
rect 10965 39457 10977 39491
rect 11011 39488 11023 39491
rect 12434 39488 12440 39500
rect 11011 39460 12440 39488
rect 11011 39457 11023 39460
rect 10965 39451 11023 39457
rect 12434 39448 12440 39460
rect 12492 39448 12498 39500
rect 12820 39488 12848 39528
rect 13265 39525 13277 39528
rect 13311 39556 13323 39559
rect 13814 39556 13820 39568
rect 13311 39528 13820 39556
rect 13311 39525 13323 39528
rect 13265 39519 13323 39525
rect 13814 39516 13820 39528
rect 13872 39516 13878 39568
rect 14369 39559 14427 39565
rect 14369 39525 14381 39559
rect 14415 39556 14427 39559
rect 15838 39556 15844 39568
rect 14415 39528 15844 39556
rect 14415 39525 14427 39528
rect 14369 39519 14427 39525
rect 15838 39516 15844 39528
rect 15896 39516 15902 39568
rect 16022 39516 16028 39568
rect 16080 39556 16086 39568
rect 25130 39556 25136 39568
rect 16080 39528 25136 39556
rect 16080 39516 16086 39528
rect 25130 39516 25136 39528
rect 25188 39516 25194 39568
rect 13446 39488 13452 39500
rect 12820 39460 13452 39488
rect 13446 39448 13452 39460
rect 13504 39448 13510 39500
rect 15013 39491 15071 39497
rect 15013 39457 15025 39491
rect 15059 39488 15071 39491
rect 15654 39488 15660 39500
rect 15059 39460 15660 39488
rect 15059 39457 15071 39460
rect 15013 39451 15071 39457
rect 15654 39448 15660 39460
rect 15712 39448 15718 39500
rect 16209 39491 16267 39497
rect 16209 39457 16221 39491
rect 16255 39488 16267 39491
rect 17770 39488 17776 39500
rect 16255 39460 17776 39488
rect 16255 39457 16267 39460
rect 16209 39451 16267 39457
rect 17770 39448 17776 39460
rect 17828 39448 17834 39500
rect 19426 39448 19432 39500
rect 19484 39488 19490 39500
rect 19889 39491 19947 39497
rect 19889 39488 19901 39491
rect 19484 39460 19901 39488
rect 19484 39448 19490 39460
rect 19889 39457 19901 39460
rect 19935 39457 19947 39491
rect 19889 39451 19947 39457
rect 20070 39448 20076 39500
rect 20128 39448 20134 39500
rect 21542 39448 21548 39500
rect 21600 39488 21606 39500
rect 21913 39491 21971 39497
rect 21913 39488 21925 39491
rect 21600 39460 21925 39488
rect 21600 39448 21606 39460
rect 21913 39457 21925 39460
rect 21959 39488 21971 39491
rect 22186 39488 22192 39500
rect 21959 39460 22192 39488
rect 21959 39457 21971 39460
rect 21913 39451 21971 39457
rect 22186 39448 22192 39460
rect 22244 39488 22250 39500
rect 22281 39491 22339 39497
rect 22281 39488 22293 39491
rect 22244 39460 22293 39488
rect 22244 39448 22250 39460
rect 22281 39457 22293 39460
rect 22327 39457 22339 39491
rect 22281 39451 22339 39457
rect 23293 39491 23351 39497
rect 23293 39457 23305 39491
rect 23339 39488 23351 39491
rect 23474 39488 23480 39500
rect 23339 39460 23480 39488
rect 23339 39457 23351 39460
rect 23293 39451 23351 39457
rect 23474 39448 23480 39460
rect 23532 39448 23538 39500
rect 25038 39448 25044 39500
rect 25096 39448 25102 39500
rect 25222 39448 25228 39500
rect 25280 39448 25286 39500
rect 15838 39420 15844 39432
rect 13740 39392 15844 39420
rect 5169 39355 5227 39361
rect 5169 39321 5181 39355
rect 5215 39321 5227 39355
rect 6917 39355 6975 39361
rect 6917 39352 6929 39355
rect 6394 39324 6929 39352
rect 5169 39315 5227 39321
rect 6917 39321 6929 39324
rect 6963 39352 6975 39355
rect 7282 39352 7288 39364
rect 6963 39324 7288 39352
rect 6963 39321 6975 39324
rect 6917 39315 6975 39321
rect 5184 39284 5212 39315
rect 7282 39312 7288 39324
rect 7340 39312 7346 39364
rect 10137 39355 10195 39361
rect 10137 39321 10149 39355
rect 10183 39352 10195 39355
rect 10183 39324 11192 39352
rect 10183 39321 10195 39324
rect 10137 39315 10195 39321
rect 5810 39284 5816 39296
rect 5184 39256 5816 39284
rect 5810 39244 5816 39256
rect 5868 39244 5874 39296
rect 8294 39244 8300 39296
rect 8352 39284 8358 39296
rect 9125 39287 9183 39293
rect 9125 39284 9137 39287
rect 8352 39256 9137 39284
rect 8352 39244 8358 39256
rect 9125 39253 9137 39256
rect 9171 39253 9183 39287
rect 11164 39284 11192 39324
rect 11514 39312 11520 39364
rect 11572 39352 11578 39364
rect 11572 39324 11730 39352
rect 11572 39312 11578 39324
rect 13740 39284 13768 39392
rect 15838 39380 15844 39392
rect 15896 39380 15902 39432
rect 16960 39392 20208 39420
rect 14829 39355 14887 39361
rect 14829 39352 14841 39355
rect 13832 39324 14841 39352
rect 13832 39296 13860 39324
rect 14829 39321 14841 39324
rect 14875 39321 14887 39355
rect 14829 39315 14887 39321
rect 15010 39312 15016 39364
rect 15068 39352 15074 39364
rect 16960 39352 16988 39392
rect 15068 39324 16988 39352
rect 15068 39312 15074 39324
rect 17034 39312 17040 39364
rect 17092 39352 17098 39364
rect 19797 39355 19855 39361
rect 19797 39352 19809 39355
rect 17092 39324 19809 39352
rect 17092 39312 17098 39324
rect 19797 39321 19809 39324
rect 19843 39321 19855 39355
rect 20180 39352 20208 39392
rect 20254 39380 20260 39432
rect 20312 39420 20318 39432
rect 23109 39423 23167 39429
rect 23109 39420 23121 39423
rect 20312 39392 23121 39420
rect 20312 39380 20318 39392
rect 23109 39389 23121 39392
rect 23155 39389 23167 39423
rect 23109 39383 23167 39389
rect 20180 39324 21680 39352
rect 19797 39315 19855 39321
rect 11164 39256 13768 39284
rect 9125 39247 9183 39253
rect 13814 39244 13820 39296
rect 13872 39244 13878 39296
rect 14734 39244 14740 39296
rect 14792 39244 14798 39296
rect 15378 39244 15384 39296
rect 15436 39284 15442 39296
rect 15933 39287 15991 39293
rect 15933 39284 15945 39287
rect 15436 39256 15945 39284
rect 15436 39244 15442 39256
rect 15933 39253 15945 39256
rect 15979 39253 15991 39287
rect 15933 39247 15991 39253
rect 16022 39244 16028 39296
rect 16080 39244 16086 39296
rect 18414 39244 18420 39296
rect 18472 39284 18478 39296
rect 18601 39287 18659 39293
rect 18601 39284 18613 39287
rect 18472 39256 18613 39284
rect 18472 39244 18478 39256
rect 18601 39253 18613 39256
rect 18647 39253 18659 39287
rect 18601 39247 18659 39253
rect 19429 39287 19487 39293
rect 19429 39253 19441 39287
rect 19475 39284 19487 39287
rect 19886 39284 19892 39296
rect 19475 39256 19892 39284
rect 19475 39253 19487 39256
rect 19429 39247 19487 39253
rect 19886 39244 19892 39256
rect 19944 39244 19950 39296
rect 21652 39293 21680 39324
rect 21726 39312 21732 39364
rect 21784 39312 21790 39364
rect 22738 39352 22744 39364
rect 22112 39324 22744 39352
rect 21637 39287 21695 39293
rect 21637 39253 21649 39287
rect 21683 39284 21695 39287
rect 22112 39284 22140 39324
rect 22738 39312 22744 39324
rect 22796 39312 22802 39364
rect 23017 39355 23075 39361
rect 23017 39321 23029 39355
rect 23063 39352 23075 39355
rect 23845 39355 23903 39361
rect 23845 39352 23857 39355
rect 23063 39324 23857 39352
rect 23063 39321 23075 39324
rect 23017 39315 23075 39321
rect 23845 39321 23857 39324
rect 23891 39321 23903 39355
rect 24949 39355 25007 39361
rect 24949 39352 24961 39355
rect 23845 39315 23903 39321
rect 23952 39324 24961 39352
rect 21683 39256 22140 39284
rect 22649 39287 22707 39293
rect 21683 39253 21695 39256
rect 21637 39247 21695 39253
rect 22649 39253 22661 39287
rect 22695 39284 22707 39287
rect 23952 39284 23980 39324
rect 24949 39321 24961 39324
rect 24995 39321 25007 39355
rect 24949 39315 25007 39321
rect 22695 39256 23980 39284
rect 24581 39287 24639 39293
rect 22695 39253 22707 39256
rect 22649 39247 22707 39253
rect 24581 39253 24593 39287
rect 24627 39284 24639 39287
rect 24762 39284 24768 39296
rect 24627 39256 24768 39284
rect 24627 39253 24639 39256
rect 24581 39247 24639 39253
rect 24762 39244 24768 39256
rect 24820 39244 24826 39296
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 7282 39040 7288 39092
rect 7340 39040 7346 39092
rect 8205 39083 8263 39089
rect 8205 39049 8217 39083
rect 8251 39080 8263 39083
rect 9490 39080 9496 39092
rect 8251 39052 9496 39080
rect 8251 39049 8263 39052
rect 8205 39043 8263 39049
rect 9490 39040 9496 39052
rect 9548 39040 9554 39092
rect 10781 39083 10839 39089
rect 10781 39049 10793 39083
rect 10827 39080 10839 39083
rect 10962 39080 10968 39092
rect 10827 39052 10968 39080
rect 10827 39049 10839 39052
rect 10781 39043 10839 39049
rect 10962 39040 10968 39052
rect 11020 39040 11026 39092
rect 13722 39080 13728 39092
rect 11624 39052 13728 39080
rect 7300 39012 7328 39040
rect 8665 39015 8723 39021
rect 8665 39012 8677 39015
rect 7300 38984 8677 39012
rect 8665 38981 8677 38984
rect 8711 38981 8723 39015
rect 8665 38975 8723 38981
rect 10873 39015 10931 39021
rect 10873 38981 10885 39015
rect 10919 39012 10931 39015
rect 11514 39012 11520 39024
rect 10919 38984 11520 39012
rect 10919 38981 10931 38984
rect 10873 38975 10931 38981
rect 11514 38972 11520 38984
rect 11572 38972 11578 39024
rect 4062 38904 4068 38956
rect 4120 38944 4126 38956
rect 8297 38947 8355 38953
rect 8297 38944 8309 38947
rect 4120 38916 8309 38944
rect 4120 38904 4126 38916
rect 8297 38913 8309 38916
rect 8343 38944 8355 38947
rect 9585 38947 9643 38953
rect 9585 38944 9597 38947
rect 8343 38916 9597 38944
rect 8343 38913 8355 38916
rect 8297 38907 8355 38913
rect 9585 38913 9597 38916
rect 9631 38913 9643 38947
rect 9585 38907 9643 38913
rect 8573 38811 8631 38817
rect 8573 38777 8585 38811
rect 8619 38808 8631 38811
rect 9490 38808 9496 38820
rect 8619 38780 9496 38808
rect 8619 38777 8631 38780
rect 8573 38771 8631 38777
rect 9490 38768 9496 38780
rect 9548 38768 9554 38820
rect 1394 38700 1400 38752
rect 1452 38700 1458 38752
rect 9122 38700 9128 38752
rect 9180 38700 9186 38752
rect 9600 38740 9628 38907
rect 9674 38836 9680 38888
rect 9732 38836 9738 38888
rect 10962 38836 10968 38888
rect 11020 38876 11026 38888
rect 11057 38879 11115 38885
rect 11057 38876 11069 38879
rect 11020 38848 11069 38876
rect 11020 38836 11026 38848
rect 11057 38845 11069 38848
rect 11103 38876 11115 38879
rect 11624 38876 11652 39052
rect 13722 39040 13728 39052
rect 13780 39040 13786 39092
rect 14277 39083 14335 39089
rect 14277 39049 14289 39083
rect 14323 39080 14335 39083
rect 14734 39080 14740 39092
rect 14323 39052 14740 39080
rect 14323 39049 14335 39052
rect 14277 39043 14335 39049
rect 14734 39040 14740 39052
rect 14792 39040 14798 39092
rect 14826 39040 14832 39092
rect 14884 39080 14890 39092
rect 15010 39080 15016 39092
rect 14884 39052 15016 39080
rect 14884 39040 14890 39052
rect 15010 39040 15016 39052
rect 15068 39040 15074 39092
rect 15289 39083 15347 39089
rect 15289 39049 15301 39083
rect 15335 39080 15347 39083
rect 15930 39080 15936 39092
rect 15335 39052 15936 39080
rect 15335 39049 15347 39052
rect 15289 39043 15347 39049
rect 15930 39040 15936 39052
rect 15988 39040 15994 39092
rect 16022 39040 16028 39092
rect 16080 39080 16086 39092
rect 19153 39083 19211 39089
rect 19153 39080 19165 39083
rect 16080 39052 19165 39080
rect 16080 39040 16086 39052
rect 19153 39049 19165 39052
rect 19199 39049 19211 39083
rect 19153 39043 19211 39049
rect 20717 39083 20775 39089
rect 20717 39049 20729 39083
rect 20763 39080 20775 39083
rect 20990 39080 20996 39092
rect 20763 39052 20996 39080
rect 20763 39049 20775 39052
rect 20717 39043 20775 39049
rect 20990 39040 20996 39052
rect 21048 39040 21054 39092
rect 22094 39040 22100 39092
rect 22152 39080 22158 39092
rect 24489 39083 24547 39089
rect 24489 39080 24501 39083
rect 22152 39052 24501 39080
rect 22152 39040 22158 39052
rect 24489 39049 24501 39052
rect 24535 39049 24547 39083
rect 24489 39043 24547 39049
rect 12434 39012 12440 39024
rect 12084 38984 12440 39012
rect 12084 38953 12112 38984
rect 12434 38972 12440 38984
rect 12492 38972 12498 39024
rect 13078 38972 13084 39024
rect 13136 38972 13142 39024
rect 18325 39015 18383 39021
rect 18325 38981 18337 39015
rect 18371 39012 18383 39015
rect 18506 39012 18512 39024
rect 18371 38984 18512 39012
rect 18371 38981 18383 38984
rect 18325 38975 18383 38981
rect 18506 38972 18512 38984
rect 18564 38972 18570 39024
rect 19613 39015 19671 39021
rect 19613 38981 19625 39015
rect 19659 39012 19671 39015
rect 20806 39012 20812 39024
rect 19659 38984 20812 39012
rect 19659 38981 19671 38984
rect 19613 38975 19671 38981
rect 20806 38972 20812 38984
rect 20864 38972 20870 39024
rect 23658 38972 23664 39024
rect 23716 39012 23722 39024
rect 24121 39015 24179 39021
rect 24121 39012 24133 39015
rect 23716 38984 24133 39012
rect 23716 38972 23722 38984
rect 24121 38981 24133 38984
rect 24167 39012 24179 39015
rect 25406 39012 25412 39024
rect 24167 38984 25412 39012
rect 24167 38981 24179 38984
rect 24121 38975 24179 38981
rect 25406 38972 25412 38984
rect 25464 38972 25470 39024
rect 12069 38947 12127 38953
rect 12069 38913 12081 38947
rect 12115 38913 12127 38947
rect 12069 38907 12127 38913
rect 19521 38947 19579 38953
rect 19521 38913 19533 38947
rect 19567 38944 19579 38947
rect 21358 38944 21364 38956
rect 19567 38916 21364 38944
rect 19567 38913 19579 38916
rect 19521 38907 19579 38913
rect 21358 38904 21364 38916
rect 21416 38904 21422 38956
rect 23506 38916 24164 38944
rect 11103 38848 11652 38876
rect 12345 38879 12403 38885
rect 11103 38845 11115 38848
rect 11057 38839 11115 38845
rect 12345 38845 12357 38879
rect 12391 38876 12403 38879
rect 14642 38876 14648 38888
rect 12391 38848 14648 38876
rect 12391 38845 12403 38848
rect 12345 38839 12403 38845
rect 14642 38836 14648 38848
rect 14700 38836 14706 38888
rect 15381 38879 15439 38885
rect 15381 38845 15393 38879
rect 15427 38845 15439 38879
rect 15381 38839 15439 38845
rect 10413 38811 10471 38817
rect 10413 38777 10425 38811
rect 10459 38808 10471 38811
rect 11146 38808 11152 38820
rect 10459 38780 11152 38808
rect 10459 38777 10471 38780
rect 10413 38771 10471 38777
rect 11146 38768 11152 38780
rect 11204 38768 11210 38820
rect 11974 38808 11980 38820
rect 11243 38780 11980 38808
rect 11243 38740 11271 38780
rect 11974 38768 11980 38780
rect 12032 38768 12038 38820
rect 14921 38811 14979 38817
rect 14921 38808 14933 38811
rect 13648 38780 14933 38808
rect 9600 38712 11271 38740
rect 11514 38700 11520 38752
rect 11572 38700 11578 38752
rect 11698 38700 11704 38752
rect 11756 38740 11762 38752
rect 13648 38740 13676 38780
rect 14921 38777 14933 38780
rect 14967 38777 14979 38811
rect 15396 38808 15424 38839
rect 15562 38836 15568 38888
rect 15620 38836 15626 38888
rect 16850 38836 16856 38888
rect 16908 38836 16914 38888
rect 18414 38836 18420 38888
rect 18472 38836 18478 38888
rect 18601 38879 18659 38885
rect 18601 38845 18613 38879
rect 18647 38876 18659 38879
rect 19150 38876 19156 38888
rect 18647 38848 19156 38876
rect 18647 38845 18659 38848
rect 18601 38839 18659 38845
rect 19150 38836 19156 38848
rect 19208 38836 19214 38888
rect 19705 38879 19763 38885
rect 19705 38845 19717 38879
rect 19751 38845 19763 38879
rect 19705 38839 19763 38845
rect 15396 38780 16068 38808
rect 14921 38771 14979 38777
rect 16040 38752 16068 38780
rect 18322 38768 18328 38820
rect 18380 38808 18386 38820
rect 19720 38808 19748 38839
rect 20438 38836 20444 38888
rect 20496 38876 20502 38888
rect 20809 38879 20867 38885
rect 20809 38876 20821 38879
rect 20496 38848 20821 38876
rect 20496 38836 20502 38848
rect 20809 38845 20821 38848
rect 20855 38845 20867 38879
rect 20809 38839 20867 38845
rect 20990 38836 20996 38888
rect 21048 38836 21054 38888
rect 22104 38879 22162 38885
rect 22104 38845 22116 38879
rect 22150 38876 22162 38879
rect 22373 38879 22431 38885
rect 22150 38848 22232 38876
rect 22150 38845 22162 38848
rect 22104 38839 22162 38845
rect 18380 38780 19748 38808
rect 18380 38768 18386 38780
rect 11756 38712 13676 38740
rect 13817 38743 13875 38749
rect 11756 38700 11762 38712
rect 13817 38709 13829 38743
rect 13863 38740 13875 38743
rect 13998 38740 14004 38752
rect 13863 38712 14004 38740
rect 13863 38709 13875 38712
rect 13817 38703 13875 38709
rect 13998 38700 14004 38712
rect 14056 38700 14062 38752
rect 16022 38700 16028 38752
rect 16080 38700 16086 38752
rect 16574 38700 16580 38752
rect 16632 38740 16638 38752
rect 17957 38743 18015 38749
rect 17957 38740 17969 38743
rect 16632 38712 17969 38740
rect 16632 38700 16638 38712
rect 17957 38709 17969 38712
rect 18003 38709 18015 38743
rect 17957 38703 18015 38709
rect 18506 38700 18512 38752
rect 18564 38740 18570 38752
rect 18690 38740 18696 38752
rect 18564 38712 18696 38740
rect 18564 38700 18570 38712
rect 18690 38700 18696 38712
rect 18748 38700 18754 38752
rect 20346 38700 20352 38752
rect 20404 38700 20410 38752
rect 20438 38700 20444 38752
rect 20496 38740 20502 38752
rect 22094 38740 22100 38752
rect 20496 38712 22100 38740
rect 20496 38700 20502 38712
rect 22094 38700 22100 38712
rect 22152 38700 22158 38752
rect 22204 38740 22232 38848
rect 22373 38845 22385 38879
rect 22419 38876 22431 38879
rect 23106 38876 23112 38888
rect 22419 38848 23112 38876
rect 22419 38845 22431 38848
rect 22373 38839 22431 38845
rect 23106 38836 23112 38848
rect 23164 38876 23170 38888
rect 23750 38876 23756 38888
rect 23164 38848 23756 38876
rect 23164 38836 23170 38848
rect 23750 38836 23756 38848
rect 23808 38836 23814 38888
rect 24136 38876 24164 38916
rect 24210 38904 24216 38956
rect 24268 38944 24274 38956
rect 24673 38947 24731 38953
rect 24673 38944 24685 38947
rect 24268 38916 24685 38944
rect 24268 38904 24274 38916
rect 24673 38913 24685 38916
rect 24719 38944 24731 38947
rect 24854 38944 24860 38956
rect 24719 38916 24860 38944
rect 24719 38913 24731 38916
rect 24673 38907 24731 38913
rect 24854 38904 24860 38916
rect 24912 38904 24918 38956
rect 25314 38904 25320 38956
rect 25372 38904 25378 38956
rect 24578 38876 24584 38888
rect 24136 38848 24584 38876
rect 24578 38836 24584 38848
rect 24636 38836 24642 38888
rect 22830 38740 22836 38752
rect 22204 38712 22836 38740
rect 22830 38700 22836 38712
rect 22888 38700 22894 38752
rect 23658 38700 23664 38752
rect 23716 38740 23722 38752
rect 23845 38743 23903 38749
rect 23845 38740 23857 38743
rect 23716 38712 23857 38740
rect 23716 38700 23722 38712
rect 23845 38709 23857 38712
rect 23891 38709 23903 38743
rect 23845 38703 23903 38709
rect 25130 38700 25136 38752
rect 25188 38700 25194 38752
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 6914 38496 6920 38548
rect 6972 38536 6978 38548
rect 7190 38536 7196 38548
rect 6972 38508 7196 38536
rect 6972 38496 6978 38508
rect 7190 38496 7196 38508
rect 7248 38496 7254 38548
rect 7742 38496 7748 38548
rect 7800 38536 7806 38548
rect 7837 38539 7895 38545
rect 7837 38536 7849 38539
rect 7800 38508 7849 38536
rect 7800 38496 7806 38508
rect 7837 38505 7849 38508
rect 7883 38505 7895 38539
rect 9858 38536 9864 38548
rect 7837 38499 7895 38505
rect 8588 38508 9864 38536
rect 8588 38480 8616 38508
rect 9858 38496 9864 38508
rect 9916 38536 9922 38548
rect 10318 38536 10324 38548
rect 9916 38508 10324 38536
rect 9916 38496 9922 38508
rect 10318 38496 10324 38508
rect 10376 38496 10382 38548
rect 10413 38539 10471 38545
rect 10413 38505 10425 38539
rect 10459 38536 10471 38539
rect 11054 38536 11060 38548
rect 10459 38508 11060 38536
rect 10459 38505 10471 38508
rect 10413 38499 10471 38505
rect 11054 38496 11060 38508
rect 11112 38496 11118 38548
rect 12342 38496 12348 38548
rect 12400 38536 12406 38548
rect 14277 38539 14335 38545
rect 14277 38536 14289 38539
rect 12400 38508 14289 38536
rect 12400 38496 12406 38508
rect 14277 38505 14289 38508
rect 14323 38505 14335 38539
rect 14277 38499 14335 38505
rect 15838 38496 15844 38548
rect 15896 38536 15902 38548
rect 15896 38508 17264 38536
rect 15896 38496 15902 38508
rect 8570 38468 8576 38480
rect 6840 38440 8576 38468
rect 5721 38403 5779 38409
rect 5721 38369 5733 38403
rect 5767 38400 5779 38403
rect 6840 38400 6868 38440
rect 8570 38428 8576 38440
rect 8628 38428 8634 38480
rect 10134 38428 10140 38480
rect 10192 38468 10198 38480
rect 11885 38471 11943 38477
rect 11885 38468 11897 38471
rect 10192 38440 11897 38468
rect 10192 38428 10198 38440
rect 11885 38437 11897 38440
rect 11931 38437 11943 38471
rect 13446 38468 13452 38480
rect 11885 38431 11943 38437
rect 11992 38440 13452 38468
rect 5767 38372 6868 38400
rect 5767 38369 5779 38372
rect 5721 38363 5779 38369
rect 6914 38360 6920 38412
rect 6972 38400 6978 38412
rect 7193 38403 7251 38409
rect 7193 38400 7205 38403
rect 6972 38372 7205 38400
rect 6972 38360 6978 38372
rect 7193 38369 7205 38372
rect 7239 38400 7251 38403
rect 7834 38400 7840 38412
rect 7239 38372 7840 38400
rect 7239 38369 7251 38372
rect 7193 38363 7251 38369
rect 7834 38360 7840 38372
rect 7892 38360 7898 38412
rect 8481 38403 8539 38409
rect 8481 38369 8493 38403
rect 8527 38369 8539 38403
rect 8481 38363 8539 38369
rect 1302 38292 1308 38344
rect 1360 38332 1366 38344
rect 1581 38335 1639 38341
rect 1581 38332 1593 38335
rect 1360 38304 1593 38332
rect 1360 38292 1366 38304
rect 1581 38301 1593 38304
rect 1627 38301 1639 38335
rect 1581 38295 1639 38301
rect 5445 38335 5503 38341
rect 5445 38301 5457 38335
rect 5491 38301 5503 38335
rect 5445 38295 5503 38301
rect 8205 38335 8263 38341
rect 8205 38301 8217 38335
rect 8251 38332 8263 38335
rect 8294 38332 8300 38344
rect 8251 38304 8300 38332
rect 8251 38301 8263 38304
rect 8205 38295 8263 38301
rect 1762 38156 1768 38208
rect 1820 38196 1826 38208
rect 2225 38199 2283 38205
rect 2225 38196 2237 38199
rect 1820 38168 2237 38196
rect 1820 38156 1826 38168
rect 2225 38165 2237 38168
rect 2271 38165 2283 38199
rect 5460 38196 5488 38295
rect 8294 38292 8300 38304
rect 8352 38292 8358 38344
rect 7374 38264 7380 38276
rect 6946 38236 7380 38264
rect 7374 38224 7380 38236
rect 7432 38224 7438 38276
rect 7558 38224 7564 38276
rect 7616 38264 7622 38276
rect 8496 38264 8524 38363
rect 9122 38360 9128 38412
rect 9180 38400 9186 38412
rect 9677 38403 9735 38409
rect 9677 38400 9689 38403
rect 9180 38372 9689 38400
rect 9180 38360 9186 38372
rect 9677 38369 9689 38372
rect 9723 38369 9735 38403
rect 9677 38363 9735 38369
rect 9769 38403 9827 38409
rect 9769 38369 9781 38403
rect 9815 38369 9827 38403
rect 9769 38363 9827 38369
rect 9214 38292 9220 38344
rect 9272 38332 9278 38344
rect 9784 38332 9812 38363
rect 10226 38360 10232 38412
rect 10284 38400 10290 38412
rect 10965 38403 11023 38409
rect 10965 38400 10977 38403
rect 10284 38372 10977 38400
rect 10284 38360 10290 38372
rect 10965 38369 10977 38372
rect 11011 38400 11023 38403
rect 11992 38400 12020 38440
rect 13446 38428 13452 38440
rect 13504 38468 13510 38480
rect 17236 38468 17264 38508
rect 17862 38496 17868 38548
rect 17920 38536 17926 38548
rect 19429 38539 19487 38545
rect 19429 38536 19441 38539
rect 17920 38508 19441 38536
rect 17920 38496 17926 38508
rect 19429 38505 19441 38508
rect 19475 38505 19487 38539
rect 25958 38536 25964 38548
rect 19429 38499 19487 38505
rect 21652 38508 25964 38536
rect 18141 38471 18199 38477
rect 18141 38468 18153 38471
rect 13504 38440 14872 38468
rect 17236 38440 18153 38468
rect 13504 38428 13510 38440
rect 11011 38372 12020 38400
rect 11011 38369 11023 38372
rect 10965 38363 11023 38369
rect 12158 38360 12164 38412
rect 12216 38400 12222 38412
rect 12345 38403 12403 38409
rect 12345 38400 12357 38403
rect 12216 38372 12357 38400
rect 12216 38360 12222 38372
rect 12345 38369 12357 38372
rect 12391 38369 12403 38403
rect 12345 38363 12403 38369
rect 12437 38403 12495 38409
rect 12437 38369 12449 38403
rect 12483 38369 12495 38403
rect 12437 38363 12495 38369
rect 12452 38332 12480 38363
rect 13262 38360 13268 38412
rect 13320 38360 13326 38412
rect 13909 38403 13967 38409
rect 13909 38369 13921 38403
rect 13955 38400 13967 38403
rect 14274 38400 14280 38412
rect 13955 38372 14280 38400
rect 13955 38369 13967 38372
rect 13909 38363 13967 38369
rect 14274 38360 14280 38372
rect 14332 38360 14338 38412
rect 14844 38409 14872 38440
rect 18141 38437 18153 38440
rect 18187 38437 18199 38471
rect 20806 38468 20812 38480
rect 18141 38431 18199 38437
rect 18524 38440 20812 38468
rect 14829 38403 14887 38409
rect 14829 38369 14841 38403
rect 14875 38369 14887 38403
rect 18322 38400 18328 38412
rect 14829 38363 14887 38369
rect 15856 38372 18328 38400
rect 9272 38304 9812 38332
rect 9876 38304 12480 38332
rect 9272 38292 9278 38304
rect 9876 38264 9904 38304
rect 12710 38292 12716 38344
rect 12768 38332 12774 38344
rect 13280 38332 13308 38360
rect 12768 38304 13308 38332
rect 14737 38335 14795 38341
rect 12768 38292 12774 38304
rect 14737 38301 14749 38335
rect 14783 38332 14795 38335
rect 15194 38332 15200 38344
rect 14783 38304 15200 38332
rect 14783 38301 14795 38304
rect 14737 38295 14795 38301
rect 15194 38292 15200 38304
rect 15252 38292 15258 38344
rect 7616 38236 9904 38264
rect 7616 38224 7622 38236
rect 11974 38224 11980 38276
rect 12032 38264 12038 38276
rect 15102 38264 15108 38276
rect 12032 38236 15108 38264
rect 12032 38224 12038 38236
rect 15102 38224 15108 38236
rect 15160 38224 15166 38276
rect 15654 38224 15660 38276
rect 15712 38264 15718 38276
rect 15856 38264 15884 38372
rect 18322 38360 18328 38372
rect 18380 38360 18386 38412
rect 15930 38292 15936 38344
rect 15988 38292 15994 38344
rect 17310 38292 17316 38344
rect 17368 38292 17374 38344
rect 18524 38341 18552 38440
rect 20806 38428 20812 38440
rect 20864 38428 20870 38480
rect 18690 38360 18696 38412
rect 18748 38360 18754 38412
rect 18874 38360 18880 38412
rect 18932 38400 18938 38412
rect 19981 38403 20039 38409
rect 19981 38400 19993 38403
rect 18932 38372 19993 38400
rect 18932 38360 18938 38372
rect 19981 38369 19993 38372
rect 20027 38369 20039 38403
rect 19981 38363 20039 38369
rect 21082 38360 21088 38412
rect 21140 38360 21146 38412
rect 21266 38360 21272 38412
rect 21324 38360 21330 38412
rect 18509 38335 18567 38341
rect 18509 38301 18521 38335
rect 18555 38301 18567 38335
rect 18509 38295 18567 38301
rect 18601 38335 18659 38341
rect 18601 38301 18613 38335
rect 18647 38332 18659 38335
rect 19058 38332 19064 38344
rect 18647 38304 19064 38332
rect 18647 38301 18659 38304
rect 18601 38295 18659 38301
rect 19058 38292 19064 38304
rect 19116 38292 19122 38344
rect 19889 38335 19947 38341
rect 19889 38301 19901 38335
rect 19935 38332 19947 38335
rect 20438 38332 20444 38344
rect 19935 38304 20444 38332
rect 19935 38301 19947 38304
rect 19889 38295 19947 38301
rect 20438 38292 20444 38304
rect 20496 38292 20502 38344
rect 20622 38292 20628 38344
rect 20680 38332 20686 38344
rect 21652 38341 21680 38508
rect 25958 38496 25964 38508
rect 26016 38496 26022 38548
rect 22278 38428 22284 38480
rect 22336 38468 22342 38480
rect 24670 38468 24676 38480
rect 22336 38440 24676 38468
rect 22336 38428 22342 38440
rect 24670 38428 24676 38440
rect 24728 38428 24734 38480
rect 21910 38360 21916 38412
rect 21968 38400 21974 38412
rect 22465 38403 22523 38409
rect 22465 38400 22477 38403
rect 21968 38372 22477 38400
rect 21968 38360 21974 38372
rect 22465 38369 22477 38372
rect 22511 38369 22523 38403
rect 22465 38363 22523 38369
rect 22646 38360 22652 38412
rect 22704 38400 22710 38412
rect 23658 38400 23664 38412
rect 22704 38372 23664 38400
rect 22704 38360 22710 38372
rect 23658 38360 23664 38372
rect 23716 38360 23722 38412
rect 23750 38360 23756 38412
rect 23808 38360 23814 38412
rect 24946 38360 24952 38412
rect 25004 38400 25010 38412
rect 25041 38403 25099 38409
rect 25041 38400 25053 38403
rect 25004 38372 25053 38400
rect 25004 38360 25010 38372
rect 25041 38369 25053 38372
rect 25087 38369 25099 38403
rect 25041 38363 25099 38369
rect 25133 38403 25191 38409
rect 25133 38369 25145 38403
rect 25179 38369 25191 38403
rect 25133 38363 25191 38369
rect 21637 38335 21695 38341
rect 21637 38332 21649 38335
rect 20680 38304 21649 38332
rect 20680 38292 20686 38304
rect 21637 38301 21649 38304
rect 21683 38301 21695 38335
rect 21637 38295 21695 38301
rect 23842 38292 23848 38344
rect 23900 38332 23906 38344
rect 25148 38332 25176 38363
rect 23900 38304 25176 38332
rect 23900 38292 23906 38304
rect 16209 38267 16267 38273
rect 16209 38264 16221 38267
rect 15712 38236 16221 38264
rect 15712 38224 15718 38236
rect 16209 38233 16221 38236
rect 16255 38233 16267 38267
rect 19242 38264 19248 38276
rect 16209 38227 16267 38233
rect 17604 38236 19248 38264
rect 6546 38196 6552 38208
rect 5460 38168 6552 38196
rect 2225 38159 2283 38165
rect 6546 38156 6552 38168
rect 6604 38156 6610 38208
rect 7190 38156 7196 38208
rect 7248 38196 7254 38208
rect 7469 38199 7527 38205
rect 7469 38196 7481 38199
rect 7248 38168 7481 38196
rect 7248 38156 7254 38168
rect 7469 38165 7481 38168
rect 7515 38196 7527 38199
rect 8202 38196 8208 38208
rect 7515 38168 8208 38196
rect 7515 38165 7527 38168
rect 7469 38159 7527 38165
rect 8202 38156 8208 38168
rect 8260 38196 8266 38208
rect 8297 38199 8355 38205
rect 8297 38196 8309 38199
rect 8260 38168 8309 38196
rect 8260 38156 8266 38168
rect 8297 38165 8309 38168
rect 8343 38165 8355 38199
rect 8297 38159 8355 38165
rect 8478 38156 8484 38208
rect 8536 38196 8542 38208
rect 9217 38199 9275 38205
rect 9217 38196 9229 38199
rect 8536 38168 9229 38196
rect 8536 38156 8542 38168
rect 9217 38165 9229 38168
rect 9263 38165 9275 38199
rect 9217 38159 9275 38165
rect 9585 38199 9643 38205
rect 9585 38165 9597 38199
rect 9631 38196 9643 38199
rect 10686 38196 10692 38208
rect 9631 38168 10692 38196
rect 9631 38165 9643 38168
rect 9585 38159 9643 38165
rect 10686 38156 10692 38168
rect 10744 38156 10750 38208
rect 10778 38156 10784 38208
rect 10836 38156 10842 38208
rect 10873 38199 10931 38205
rect 10873 38165 10885 38199
rect 10919 38196 10931 38199
rect 11054 38196 11060 38208
rect 10919 38168 11060 38196
rect 10919 38165 10931 38168
rect 10873 38159 10931 38165
rect 11054 38156 11060 38168
rect 11112 38156 11118 38208
rect 12253 38199 12311 38205
rect 12253 38165 12265 38199
rect 12299 38196 12311 38199
rect 12897 38199 12955 38205
rect 12897 38196 12909 38199
rect 12299 38168 12909 38196
rect 12299 38165 12311 38168
rect 12253 38159 12311 38165
rect 12897 38165 12909 38168
rect 12943 38196 12955 38199
rect 14550 38196 14556 38208
rect 12943 38168 14556 38196
rect 12943 38165 12955 38168
rect 12897 38159 12955 38165
rect 14550 38156 14556 38168
rect 14608 38156 14614 38208
rect 14645 38199 14703 38205
rect 14645 38165 14657 38199
rect 14691 38196 14703 38199
rect 17604 38196 17632 38236
rect 19242 38224 19248 38236
rect 19300 38224 19306 38276
rect 19334 38224 19340 38276
rect 19392 38264 19398 38276
rect 19797 38267 19855 38273
rect 19797 38264 19809 38267
rect 19392 38236 19809 38264
rect 19392 38224 19398 38236
rect 19797 38233 19809 38236
rect 19843 38233 19855 38267
rect 20993 38267 21051 38273
rect 20993 38264 21005 38267
rect 19797 38227 19855 38233
rect 19904 38236 21005 38264
rect 14691 38168 17632 38196
rect 17681 38199 17739 38205
rect 14691 38165 14703 38168
rect 14645 38159 14703 38165
rect 17681 38165 17693 38199
rect 17727 38196 17739 38199
rect 17770 38196 17776 38208
rect 17727 38168 17776 38196
rect 17727 38165 17739 38168
rect 17681 38159 17739 38165
rect 17770 38156 17776 38168
rect 17828 38156 17834 38208
rect 18782 38156 18788 38208
rect 18840 38196 18846 38208
rect 19904 38196 19932 38236
rect 20993 38233 21005 38236
rect 21039 38233 21051 38267
rect 20993 38227 21051 38233
rect 22373 38267 22431 38273
rect 22373 38233 22385 38267
rect 22419 38264 22431 38267
rect 23934 38264 23940 38276
rect 22419 38236 23244 38264
rect 22419 38233 22431 38236
rect 22373 38227 22431 38233
rect 18840 38168 19932 38196
rect 20625 38199 20683 38205
rect 18840 38156 18846 38168
rect 20625 38165 20637 38199
rect 20671 38196 20683 38199
rect 21082 38196 21088 38208
rect 20671 38168 21088 38196
rect 20671 38165 20683 38168
rect 20625 38159 20683 38165
rect 21082 38156 21088 38168
rect 21140 38156 21146 38208
rect 21910 38156 21916 38208
rect 21968 38196 21974 38208
rect 23216 38205 23244 38236
rect 23584 38236 23940 38264
rect 23584 38208 23612 38236
rect 23934 38224 23940 38236
rect 23992 38224 23998 38276
rect 22005 38199 22063 38205
rect 22005 38196 22017 38199
rect 21968 38168 22017 38196
rect 21968 38156 21974 38168
rect 22005 38165 22017 38168
rect 22051 38165 22063 38199
rect 22005 38159 22063 38165
rect 23201 38199 23259 38205
rect 23201 38165 23213 38199
rect 23247 38165 23259 38199
rect 23201 38159 23259 38165
rect 23566 38156 23572 38208
rect 23624 38156 23630 38208
rect 23658 38156 23664 38208
rect 23716 38156 23722 38208
rect 23750 38156 23756 38208
rect 23808 38196 23814 38208
rect 24581 38199 24639 38205
rect 24581 38196 24593 38199
rect 23808 38168 24593 38196
rect 23808 38156 23814 38168
rect 24581 38165 24593 38168
rect 24627 38165 24639 38199
rect 24581 38159 24639 38165
rect 24670 38156 24676 38208
rect 24728 38196 24734 38208
rect 24949 38199 25007 38205
rect 24949 38196 24961 38199
rect 24728 38168 24961 38196
rect 24728 38156 24734 38168
rect 24949 38165 24961 38168
rect 24995 38165 25007 38199
rect 24949 38159 25007 38165
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 5258 37952 5264 38004
rect 5316 37952 5322 38004
rect 5721 37995 5779 38001
rect 5721 37961 5733 37995
rect 5767 37992 5779 37995
rect 9122 37992 9128 38004
rect 5767 37964 9128 37992
rect 5767 37961 5779 37964
rect 5721 37955 5779 37961
rect 9122 37952 9128 37964
rect 9180 37952 9186 38004
rect 10045 37995 10103 38001
rect 10045 37961 10057 37995
rect 10091 37992 10103 37995
rect 10502 37992 10508 38004
rect 10091 37964 10508 37992
rect 10091 37961 10103 37964
rect 10045 37955 10103 37961
rect 10502 37952 10508 37964
rect 10560 37952 10566 38004
rect 10778 37952 10784 38004
rect 10836 37992 10842 38004
rect 11701 37995 11759 38001
rect 11701 37992 11713 37995
rect 10836 37964 11713 37992
rect 10836 37952 10842 37964
rect 11701 37961 11713 37964
rect 11747 37961 11759 37995
rect 11701 37955 11759 37961
rect 12434 37952 12440 38004
rect 12492 37992 12498 38004
rect 12492 37964 12940 37992
rect 12492 37952 12498 37964
rect 6825 37927 6883 37933
rect 6825 37893 6837 37927
rect 6871 37924 6883 37927
rect 6914 37924 6920 37936
rect 6871 37896 6920 37924
rect 6871 37893 6883 37896
rect 6825 37887 6883 37893
rect 6914 37884 6920 37896
rect 6972 37884 6978 37936
rect 7558 37884 7564 37936
rect 7616 37884 7622 37936
rect 8573 37927 8631 37933
rect 8573 37893 8585 37927
rect 8619 37924 8631 37927
rect 9582 37924 9588 37936
rect 8619 37896 9588 37924
rect 8619 37893 8631 37896
rect 8573 37887 8631 37893
rect 1762 37816 1768 37868
rect 1820 37816 1826 37868
rect 4982 37816 4988 37868
rect 5040 37856 5046 37868
rect 5629 37859 5687 37865
rect 5629 37856 5641 37859
rect 5040 37828 5641 37856
rect 5040 37816 5046 37828
rect 5629 37825 5641 37828
rect 5675 37825 5687 37859
rect 5629 37819 5687 37825
rect 5810 37748 5816 37800
rect 5868 37748 5874 37800
rect 6546 37748 6552 37800
rect 6604 37748 6610 37800
rect 7374 37748 7380 37800
rect 7432 37788 7438 37800
rect 7558 37788 7564 37800
rect 7432 37760 7564 37788
rect 7432 37748 7438 37760
rect 7558 37748 7564 37760
rect 7616 37748 7622 37800
rect 7834 37748 7840 37800
rect 7892 37788 7898 37800
rect 8588 37788 8616 37887
rect 9582 37884 9588 37896
rect 9640 37924 9646 37936
rect 9640 37896 11192 37924
rect 9640 37884 9646 37896
rect 9125 37859 9183 37865
rect 9125 37825 9137 37859
rect 9171 37856 9183 37859
rect 9306 37856 9312 37868
rect 9171 37828 9312 37856
rect 9171 37825 9183 37828
rect 9125 37819 9183 37825
rect 9306 37816 9312 37828
rect 9364 37816 9370 37868
rect 9401 37859 9459 37865
rect 9401 37825 9413 37859
rect 9447 37856 9459 37859
rect 10413 37859 10471 37865
rect 10413 37856 10425 37859
rect 9447 37828 10425 37856
rect 9447 37825 9459 37828
rect 9401 37819 9459 37825
rect 10413 37825 10425 37828
rect 10459 37825 10471 37859
rect 10413 37819 10471 37825
rect 10502 37816 10508 37868
rect 10560 37816 10566 37868
rect 7892 37760 8616 37788
rect 7892 37748 7898 37760
rect 9324 37720 9352 37816
rect 10689 37791 10747 37797
rect 10689 37757 10701 37791
rect 10735 37757 10747 37791
rect 10689 37751 10747 37757
rect 9324 37692 10548 37720
rect 1581 37655 1639 37661
rect 1581 37621 1593 37655
rect 1627 37652 1639 37655
rect 2682 37652 2688 37664
rect 1627 37624 2688 37652
rect 1627 37621 1639 37624
rect 1581 37615 1639 37621
rect 2682 37612 2688 37624
rect 2740 37612 2746 37664
rect 6638 37612 6644 37664
rect 6696 37652 6702 37664
rect 8849 37655 8907 37661
rect 8849 37652 8861 37655
rect 6696 37624 8861 37652
rect 6696 37612 6702 37624
rect 8849 37621 8861 37624
rect 8895 37652 8907 37655
rect 10042 37652 10048 37664
rect 8895 37624 10048 37652
rect 8895 37621 8907 37624
rect 8849 37615 8907 37621
rect 10042 37612 10048 37624
rect 10100 37652 10106 37664
rect 10226 37652 10232 37664
rect 10100 37624 10232 37652
rect 10100 37612 10106 37624
rect 10226 37612 10232 37624
rect 10284 37612 10290 37664
rect 10520 37652 10548 37692
rect 10704 37652 10732 37751
rect 11164 37720 11192 37896
rect 11238 37884 11244 37936
rect 11296 37924 11302 37936
rect 12805 37927 12863 37933
rect 12805 37924 12817 37927
rect 11296 37896 12817 37924
rect 11296 37884 11302 37896
rect 12805 37893 12817 37896
rect 12851 37893 12863 37927
rect 12912 37924 12940 37964
rect 13538 37952 13544 38004
rect 13596 37992 13602 38004
rect 13722 37992 13728 38004
rect 13596 37964 13728 37992
rect 13596 37952 13602 37964
rect 13722 37952 13728 37964
rect 13780 37952 13786 38004
rect 14093 37995 14151 38001
rect 14093 37961 14105 37995
rect 14139 37992 14151 37995
rect 14366 37992 14372 38004
rect 14139 37964 14372 37992
rect 14139 37961 14151 37964
rect 14093 37955 14151 37961
rect 14366 37952 14372 37964
rect 14424 37992 14430 38004
rect 15470 37992 15476 38004
rect 14424 37964 15476 37992
rect 14424 37952 14430 37964
rect 15470 37952 15476 37964
rect 15528 37952 15534 38004
rect 16114 37952 16120 38004
rect 16172 37992 16178 38004
rect 16393 37995 16451 38001
rect 16393 37992 16405 37995
rect 16172 37964 16405 37992
rect 16172 37952 16178 37964
rect 16393 37961 16405 37964
rect 16439 37992 16451 37995
rect 16666 37992 16672 38004
rect 16439 37964 16672 37992
rect 16439 37961 16451 37964
rect 16393 37955 16451 37961
rect 16666 37952 16672 37964
rect 16724 37952 16730 38004
rect 16850 37952 16856 38004
rect 16908 37992 16914 38004
rect 17221 37995 17279 38001
rect 17221 37992 17233 37995
rect 16908 37964 17233 37992
rect 16908 37952 16914 37964
rect 17221 37961 17233 37964
rect 17267 37961 17279 37995
rect 17221 37955 17279 37961
rect 17310 37952 17316 38004
rect 17368 37992 17374 38004
rect 18049 37995 18107 38001
rect 18049 37992 18061 37995
rect 17368 37964 18061 37992
rect 17368 37952 17374 37964
rect 18049 37961 18061 37964
rect 18095 37992 18107 37995
rect 18230 37992 18236 38004
rect 18095 37964 18236 37992
rect 18095 37961 18107 37964
rect 18049 37955 18107 37961
rect 18230 37952 18236 37964
rect 18288 37952 18294 38004
rect 18325 37995 18383 38001
rect 18325 37961 18337 37995
rect 18371 37992 18383 37995
rect 18690 37992 18696 38004
rect 18371 37964 18696 37992
rect 18371 37961 18383 37964
rect 18325 37955 18383 37961
rect 18340 37924 18368 37955
rect 18690 37952 18696 37964
rect 18748 37952 18754 38004
rect 18969 37995 19027 38001
rect 18969 37961 18981 37995
rect 19015 37961 19027 37995
rect 18969 37955 19027 37961
rect 19429 37995 19487 38001
rect 19429 37961 19441 37995
rect 19475 37992 19487 37995
rect 20622 37992 20628 38004
rect 19475 37964 20628 37992
rect 19475 37961 19487 37964
rect 19429 37955 19487 37961
rect 18874 37924 18880 37936
rect 12912 37896 18368 37924
rect 18432 37896 18880 37924
rect 12805 37887 12863 37893
rect 12710 37816 12716 37868
rect 12768 37816 12774 37868
rect 14369 37859 14427 37865
rect 14369 37825 14381 37859
rect 14415 37856 14427 37859
rect 15381 37859 15439 37865
rect 15381 37856 15393 37859
rect 14415 37828 15393 37856
rect 14415 37825 14427 37828
rect 14369 37819 14427 37825
rect 15381 37825 15393 37828
rect 15427 37825 15439 37859
rect 15381 37819 15439 37825
rect 15473 37859 15531 37865
rect 15473 37825 15485 37859
rect 15519 37856 15531 37859
rect 16298 37856 16304 37868
rect 15519 37828 16304 37856
rect 15519 37825 15531 37828
rect 15473 37819 15531 37825
rect 16298 37816 16304 37828
rect 16356 37816 16362 37868
rect 16482 37816 16488 37868
rect 16540 37856 16546 37868
rect 17402 37856 17408 37868
rect 16540 37828 17408 37856
rect 16540 37816 16546 37828
rect 17402 37816 17408 37828
rect 17460 37856 17466 37868
rect 18432 37865 18460 37896
rect 18874 37884 18880 37896
rect 18932 37884 18938 37936
rect 18984 37924 19012 37955
rect 20622 37952 20628 37964
rect 20680 37992 20686 38004
rect 20717 37995 20775 38001
rect 20717 37992 20729 37995
rect 20680 37964 20729 37992
rect 20680 37952 20686 37964
rect 20717 37961 20729 37964
rect 20763 37961 20775 37995
rect 20717 37955 20775 37961
rect 21542 37952 21548 38004
rect 21600 37952 21606 38004
rect 22005 37995 22063 38001
rect 22005 37961 22017 37995
rect 22051 37992 22063 37995
rect 24670 37992 24676 38004
rect 22051 37964 24676 37992
rect 22051 37961 22063 37964
rect 22005 37955 22063 37961
rect 24670 37952 24676 37964
rect 24728 37952 24734 38004
rect 21450 37924 21456 37936
rect 18984 37896 21456 37924
rect 21450 37884 21456 37896
rect 21508 37884 21514 37936
rect 22462 37924 22468 37936
rect 22296 37896 22468 37924
rect 18417 37859 18475 37865
rect 18417 37856 18429 37859
rect 17460 37828 18429 37856
rect 17460 37816 17466 37828
rect 18417 37825 18429 37828
rect 18463 37825 18475 37859
rect 18417 37819 18475 37825
rect 18690 37816 18696 37868
rect 18748 37856 18754 37868
rect 19337 37859 19395 37865
rect 19337 37856 19349 37859
rect 18748 37828 19349 37856
rect 18748 37816 18754 37828
rect 19337 37825 19349 37828
rect 19383 37825 19395 37859
rect 19337 37819 19395 37825
rect 20254 37816 20260 37868
rect 20312 37856 20318 37868
rect 20625 37859 20683 37865
rect 20625 37856 20637 37859
rect 20312 37828 20637 37856
rect 20312 37816 20318 37828
rect 20625 37825 20637 37828
rect 20671 37856 20683 37859
rect 21269 37859 21327 37865
rect 21269 37856 21281 37859
rect 20671 37828 21281 37856
rect 20671 37825 20683 37828
rect 20625 37819 20683 37825
rect 21269 37825 21281 37828
rect 21315 37825 21327 37859
rect 21269 37819 21327 37825
rect 12989 37791 13047 37797
rect 12989 37757 13001 37791
rect 13035 37788 13047 37791
rect 13446 37788 13452 37800
rect 13035 37760 13452 37788
rect 13035 37757 13047 37760
rect 12989 37751 13047 37757
rect 13446 37748 13452 37760
rect 13504 37748 13510 37800
rect 13538 37748 13544 37800
rect 13596 37748 13602 37800
rect 15562 37748 15568 37800
rect 15620 37788 15626 37800
rect 15657 37791 15715 37797
rect 15657 37788 15669 37791
rect 15620 37760 15669 37788
rect 15620 37748 15626 37760
rect 15657 37757 15669 37760
rect 15703 37788 15715 37791
rect 16114 37788 16120 37800
rect 15703 37760 16120 37788
rect 15703 37757 15715 37760
rect 15657 37751 15715 37757
rect 16114 37748 16120 37760
rect 16172 37748 16178 37800
rect 16666 37748 16672 37800
rect 16724 37788 16730 37800
rect 17313 37791 17371 37797
rect 17313 37788 17325 37791
rect 16724 37760 17325 37788
rect 16724 37748 16730 37760
rect 17313 37757 17325 37760
rect 17359 37757 17371 37791
rect 17313 37751 17371 37757
rect 17497 37791 17555 37797
rect 17497 37757 17509 37791
rect 17543 37788 17555 37791
rect 18966 37788 18972 37800
rect 17543 37760 18972 37788
rect 17543 37757 17555 37760
rect 17497 37751 17555 37757
rect 18966 37748 18972 37760
rect 19024 37748 19030 37800
rect 19613 37791 19671 37797
rect 19613 37757 19625 37791
rect 19659 37788 19671 37791
rect 20530 37788 20536 37800
rect 19659 37760 20536 37788
rect 19659 37757 19671 37760
rect 19613 37751 19671 37757
rect 20530 37748 20536 37760
rect 20588 37748 20594 37800
rect 20901 37791 20959 37797
rect 20901 37757 20913 37791
rect 20947 37788 20959 37791
rect 21542 37788 21548 37800
rect 20947 37760 21548 37788
rect 20947 37757 20959 37760
rect 20901 37751 20959 37757
rect 21542 37748 21548 37760
rect 21600 37748 21606 37800
rect 17862 37720 17868 37732
rect 11164 37692 17868 37720
rect 17862 37680 17868 37692
rect 17920 37680 17926 37732
rect 18598 37720 18604 37732
rect 17972 37692 18604 37720
rect 12066 37652 12072 37664
rect 10520 37624 12072 37652
rect 12066 37612 12072 37624
rect 12124 37612 12130 37664
rect 12342 37612 12348 37664
rect 12400 37612 12406 37664
rect 15010 37612 15016 37664
rect 15068 37612 15074 37664
rect 16117 37655 16175 37661
rect 16117 37621 16129 37655
rect 16163 37652 16175 37655
rect 16298 37652 16304 37664
rect 16163 37624 16304 37652
rect 16163 37621 16175 37624
rect 16117 37615 16175 37621
rect 16298 37612 16304 37624
rect 16356 37612 16362 37664
rect 16853 37655 16911 37661
rect 16853 37621 16865 37655
rect 16899 37652 16911 37655
rect 17972 37652 18000 37692
rect 18598 37680 18604 37692
rect 18656 37680 18662 37732
rect 19058 37680 19064 37732
rect 19116 37720 19122 37732
rect 21634 37720 21640 37732
rect 19116 37692 21640 37720
rect 19116 37680 19122 37692
rect 21634 37680 21640 37692
rect 21692 37680 21698 37732
rect 16899 37624 18000 37652
rect 16899 37621 16911 37624
rect 16853 37615 16911 37621
rect 18690 37612 18696 37664
rect 18748 37612 18754 37664
rect 18966 37612 18972 37664
rect 19024 37652 19030 37664
rect 19426 37652 19432 37664
rect 19024 37624 19432 37652
rect 19024 37612 19030 37624
rect 19426 37612 19432 37624
rect 19484 37612 19490 37664
rect 20162 37612 20168 37664
rect 20220 37652 20226 37664
rect 20257 37655 20315 37661
rect 20257 37652 20269 37655
rect 20220 37624 20269 37652
rect 20220 37612 20226 37624
rect 20257 37621 20269 37624
rect 20303 37621 20315 37655
rect 20257 37615 20315 37621
rect 22002 37612 22008 37664
rect 22060 37652 22066 37664
rect 22296 37652 22324 37896
rect 22462 37884 22468 37896
rect 22520 37884 22526 37936
rect 24578 37884 24584 37936
rect 24636 37884 24642 37936
rect 22373 37859 22431 37865
rect 22373 37825 22385 37859
rect 22419 37856 22431 37859
rect 22738 37856 22744 37868
rect 22419 37828 22744 37856
rect 22419 37825 22431 37828
rect 22373 37819 22431 37825
rect 22738 37816 22744 37828
rect 22796 37856 22802 37868
rect 23201 37859 23259 37865
rect 23201 37856 23213 37859
rect 22796 37828 23213 37856
rect 22796 37816 22802 37828
rect 23201 37825 23213 37828
rect 23247 37856 23259 37859
rect 23290 37856 23296 37868
rect 23247 37828 23296 37856
rect 23247 37825 23259 37828
rect 23201 37819 23259 37825
rect 23290 37816 23296 37828
rect 23348 37816 23354 37868
rect 22462 37748 22468 37800
rect 22520 37788 22526 37800
rect 22557 37791 22615 37797
rect 22557 37788 22569 37791
rect 22520 37760 22569 37788
rect 22520 37748 22526 37760
rect 22557 37757 22569 37760
rect 22603 37757 22615 37791
rect 22557 37751 22615 37757
rect 22830 37748 22836 37800
rect 22888 37788 22894 37800
rect 23569 37791 23627 37797
rect 23569 37788 23581 37791
rect 22888 37760 23581 37788
rect 22888 37748 22894 37760
rect 23569 37757 23581 37760
rect 23615 37757 23627 37791
rect 23569 37751 23627 37757
rect 23842 37748 23848 37800
rect 23900 37748 23906 37800
rect 24486 37748 24492 37800
rect 24544 37788 24550 37800
rect 25317 37791 25375 37797
rect 25317 37788 25329 37791
rect 24544 37760 25329 37788
rect 24544 37748 24550 37760
rect 25317 37757 25329 37760
rect 25363 37757 25375 37791
rect 25317 37751 25375 37757
rect 23017 37655 23075 37661
rect 23017 37652 23029 37655
rect 22060 37624 23029 37652
rect 22060 37612 22066 37624
rect 23017 37621 23029 37624
rect 23063 37621 23075 37655
rect 23017 37615 23075 37621
rect 23474 37612 23480 37664
rect 23532 37652 23538 37664
rect 23658 37652 23664 37664
rect 23532 37624 23664 37652
rect 23532 37612 23538 37624
rect 23658 37612 23664 37624
rect 23716 37612 23722 37664
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 8570 37408 8576 37460
rect 8628 37408 8634 37460
rect 8662 37408 8668 37460
rect 8720 37448 8726 37460
rect 8720 37420 8892 37448
rect 8720 37408 8726 37420
rect 8864 37392 8892 37420
rect 10410 37408 10416 37460
rect 10468 37408 10474 37460
rect 10870 37408 10876 37460
rect 10928 37408 10934 37460
rect 14645 37451 14703 37457
rect 14645 37417 14657 37451
rect 14691 37448 14703 37451
rect 15102 37448 15108 37460
rect 14691 37420 15108 37448
rect 14691 37417 14703 37420
rect 14645 37411 14703 37417
rect 15102 37408 15108 37420
rect 15160 37408 15166 37460
rect 16298 37408 16304 37460
rect 16356 37448 16362 37460
rect 23474 37448 23480 37460
rect 16356 37420 23480 37448
rect 16356 37408 16362 37420
rect 23474 37408 23480 37420
rect 23532 37408 23538 37460
rect 23566 37408 23572 37460
rect 23624 37448 23630 37460
rect 23937 37451 23995 37457
rect 23937 37448 23949 37451
rect 23624 37420 23949 37448
rect 23624 37408 23630 37420
rect 23937 37417 23949 37420
rect 23983 37417 23995 37451
rect 23937 37411 23995 37417
rect 24670 37408 24676 37460
rect 24728 37408 24734 37460
rect 8846 37340 8852 37392
rect 8904 37380 8910 37392
rect 11514 37380 11520 37392
rect 8904 37352 11520 37380
rect 8904 37340 8910 37352
rect 11514 37340 11520 37352
rect 11572 37380 11578 37392
rect 11572 37352 11928 37380
rect 11572 37340 11578 37352
rect 7101 37315 7159 37321
rect 7101 37281 7113 37315
rect 7147 37312 7159 37315
rect 8662 37312 8668 37324
rect 7147 37284 8668 37312
rect 7147 37281 7159 37284
rect 7101 37275 7159 37281
rect 8662 37272 8668 37284
rect 8720 37312 8726 37324
rect 9398 37312 9404 37324
rect 8720 37284 9404 37312
rect 8720 37272 8726 37284
rect 9398 37272 9404 37284
rect 9456 37272 9462 37324
rect 10870 37272 10876 37324
rect 10928 37312 10934 37324
rect 11793 37315 11851 37321
rect 11793 37312 11805 37315
rect 10928 37284 11805 37312
rect 10928 37272 10934 37284
rect 11793 37281 11805 37284
rect 11839 37281 11851 37315
rect 11900 37312 11928 37352
rect 13814 37340 13820 37392
rect 13872 37380 13878 37392
rect 14185 37383 14243 37389
rect 14185 37380 14197 37383
rect 13872 37352 14197 37380
rect 13872 37340 13878 37352
rect 14185 37349 14197 37352
rect 14231 37380 14243 37383
rect 14826 37380 14832 37392
rect 14231 37352 14832 37380
rect 14231 37349 14243 37352
rect 14185 37343 14243 37349
rect 14826 37340 14832 37352
rect 14884 37340 14890 37392
rect 16390 37340 16396 37392
rect 16448 37380 16454 37392
rect 16448 37352 16712 37380
rect 16448 37340 16454 37352
rect 12437 37315 12495 37321
rect 12437 37312 12449 37315
rect 11900 37284 12449 37312
rect 11793 37275 11851 37281
rect 12437 37281 12449 37284
rect 12483 37312 12495 37315
rect 13357 37315 13415 37321
rect 13357 37312 13369 37315
rect 12483 37284 13369 37312
rect 12483 37281 12495 37284
rect 12437 37275 12495 37281
rect 13357 37281 13369 37284
rect 13403 37281 13415 37315
rect 13357 37275 13415 37281
rect 13449 37315 13507 37321
rect 13449 37281 13461 37315
rect 13495 37312 13507 37315
rect 13906 37312 13912 37324
rect 13495 37284 13912 37312
rect 13495 37281 13507 37284
rect 13449 37275 13507 37281
rect 13906 37272 13912 37284
rect 13964 37272 13970 37324
rect 15010 37312 15016 37324
rect 14016 37284 15016 37312
rect 6546 37204 6552 37256
rect 6604 37244 6610 37256
rect 6825 37247 6883 37253
rect 6825 37244 6837 37247
rect 6604 37216 6837 37244
rect 6604 37204 6610 37216
rect 6825 37213 6837 37216
rect 6871 37213 6883 37247
rect 9861 37247 9919 37253
rect 9861 37244 9873 37247
rect 6825 37207 6883 37213
rect 8404 37216 9873 37244
rect 6840 37108 6868 37207
rect 7558 37136 7564 37188
rect 7616 37136 7622 37188
rect 8404 37108 8432 37216
rect 9861 37213 9873 37216
rect 9907 37213 9919 37247
rect 9861 37207 9919 37213
rect 11609 37247 11667 37253
rect 11609 37213 11621 37247
rect 11655 37244 11667 37247
rect 13265 37247 13323 37253
rect 11655 37216 13216 37244
rect 11655 37213 11667 37216
rect 11609 37207 11667 37213
rect 9125 37179 9183 37185
rect 9125 37145 9137 37179
rect 9171 37176 9183 37179
rect 10410 37176 10416 37188
rect 9171 37148 10416 37176
rect 9171 37145 9183 37148
rect 9125 37139 9183 37145
rect 10410 37136 10416 37148
rect 10468 37136 10474 37188
rect 10686 37136 10692 37188
rect 10744 37176 10750 37188
rect 10744 37148 11652 37176
rect 10744 37136 10750 37148
rect 6840 37080 8432 37108
rect 10597 37111 10655 37117
rect 10597 37077 10609 37111
rect 10643 37108 10655 37111
rect 10778 37108 10784 37120
rect 10643 37080 10784 37108
rect 10643 37077 10655 37080
rect 10597 37071 10655 37077
rect 10778 37068 10784 37080
rect 10836 37068 10842 37120
rect 11238 37068 11244 37120
rect 11296 37068 11302 37120
rect 11624 37108 11652 37148
rect 11698 37136 11704 37188
rect 11756 37136 11762 37188
rect 13078 37176 13084 37188
rect 12406 37148 13084 37176
rect 12406 37108 12434 37148
rect 13078 37136 13084 37148
rect 13136 37136 13142 37188
rect 13188 37176 13216 37216
rect 13265 37213 13277 37247
rect 13311 37244 13323 37247
rect 13538 37244 13544 37256
rect 13311 37216 13544 37244
rect 13311 37213 13323 37216
rect 13265 37207 13323 37213
rect 13538 37204 13544 37216
rect 13596 37204 13602 37256
rect 14016 37176 14044 37284
rect 15010 37272 15016 37284
rect 15068 37272 15074 37324
rect 15194 37272 15200 37324
rect 15252 37312 15258 37324
rect 15473 37315 15531 37321
rect 15473 37312 15485 37315
rect 15252 37284 15485 37312
rect 15252 37272 15258 37284
rect 15473 37281 15485 37284
rect 15519 37281 15531 37315
rect 15473 37275 15531 37281
rect 16206 37272 16212 37324
rect 16264 37312 16270 37324
rect 16684 37321 16712 37352
rect 20530 37340 20536 37392
rect 20588 37380 20594 37392
rect 20625 37383 20683 37389
rect 20625 37380 20637 37383
rect 20588 37352 20637 37380
rect 20588 37340 20594 37352
rect 20625 37349 20637 37352
rect 20671 37349 20683 37383
rect 20625 37343 20683 37349
rect 21542 37340 21548 37392
rect 21600 37380 21606 37392
rect 25038 37380 25044 37392
rect 21600 37352 25044 37380
rect 21600 37340 21606 37352
rect 25038 37340 25044 37352
rect 25096 37340 25102 37392
rect 16577 37315 16635 37321
rect 16577 37312 16589 37315
rect 16264 37284 16589 37312
rect 16264 37272 16270 37284
rect 16577 37281 16589 37284
rect 16623 37281 16635 37315
rect 16577 37275 16635 37281
rect 16669 37315 16727 37321
rect 16669 37281 16681 37315
rect 16715 37281 16727 37315
rect 16669 37275 16727 37281
rect 17862 37272 17868 37324
rect 17920 37272 17926 37324
rect 19061 37315 19119 37321
rect 19061 37281 19073 37315
rect 19107 37312 19119 37315
rect 20254 37312 20260 37324
rect 19107 37284 20260 37312
rect 19107 37281 19119 37284
rect 19061 37275 19119 37281
rect 16485 37247 16543 37253
rect 16485 37244 16497 37247
rect 13188 37148 14044 37176
rect 14108 37216 16497 37244
rect 11624 37080 12434 37108
rect 12621 37111 12679 37117
rect 12621 37077 12633 37111
rect 12667 37108 12679 37111
rect 12710 37108 12716 37120
rect 12667 37080 12716 37108
rect 12667 37077 12679 37080
rect 12621 37071 12679 37077
rect 12710 37068 12716 37080
rect 12768 37068 12774 37120
rect 12897 37111 12955 37117
rect 12897 37077 12909 37111
rect 12943 37108 12955 37111
rect 14108 37108 14136 37216
rect 16485 37213 16497 37216
rect 16531 37213 16543 37247
rect 16485 37207 16543 37213
rect 17773 37247 17831 37253
rect 17773 37213 17785 37247
rect 17819 37244 17831 37247
rect 19076 37244 19104 37275
rect 20254 37272 20260 37284
rect 20312 37312 20318 37324
rect 24026 37312 24032 37324
rect 20312 37284 24032 37312
rect 20312 37272 20318 37284
rect 24026 37272 24032 37284
rect 24084 37272 24090 37324
rect 24581 37315 24639 37321
rect 24581 37281 24593 37315
rect 24627 37312 24639 37315
rect 24627 37284 25360 37312
rect 24627 37281 24639 37284
rect 24581 37275 24639 37281
rect 25332 37256 25360 37284
rect 20714 37244 20720 37256
rect 17819 37216 19104 37244
rect 19444 37216 20720 37244
rect 17819 37213 17831 37216
rect 17773 37207 17831 37213
rect 19444 37188 19472 37216
rect 20714 37204 20720 37216
rect 20772 37244 20778 37256
rect 21085 37247 21143 37253
rect 21085 37244 21097 37247
rect 20772 37216 21097 37244
rect 20772 37204 20778 37216
rect 21085 37213 21097 37216
rect 21131 37244 21143 37247
rect 21453 37247 21511 37253
rect 21453 37244 21465 37247
rect 21131 37216 21465 37244
rect 21131 37213 21143 37216
rect 21085 37207 21143 37213
rect 21453 37213 21465 37216
rect 21499 37213 21511 37247
rect 21453 37207 21511 37213
rect 22066 37216 24072 37244
rect 15381 37179 15439 37185
rect 15381 37145 15393 37179
rect 15427 37176 15439 37179
rect 17586 37176 17592 37188
rect 15427 37148 17592 37176
rect 15427 37145 15439 37148
rect 15381 37139 15439 37145
rect 17586 37136 17592 37148
rect 17644 37136 17650 37188
rect 17681 37179 17739 37185
rect 17681 37145 17693 37179
rect 17727 37176 17739 37179
rect 17727 37148 19380 37176
rect 17727 37145 17739 37148
rect 17681 37139 17739 37145
rect 12943 37080 14136 37108
rect 14461 37111 14519 37117
rect 12943 37077 12955 37080
rect 12897 37071 12955 37077
rect 14461 37077 14473 37111
rect 14507 37108 14519 37111
rect 14550 37108 14556 37120
rect 14507 37080 14556 37108
rect 14507 37077 14519 37080
rect 14461 37071 14519 37077
rect 14550 37068 14556 37080
rect 14608 37068 14614 37120
rect 14918 37068 14924 37120
rect 14976 37068 14982 37120
rect 15289 37111 15347 37117
rect 15289 37077 15301 37111
rect 15335 37108 15347 37111
rect 15470 37108 15476 37120
rect 15335 37080 15476 37108
rect 15335 37077 15347 37080
rect 15289 37071 15347 37077
rect 15470 37068 15476 37080
rect 15528 37068 15534 37120
rect 16117 37111 16175 37117
rect 16117 37077 16129 37111
rect 16163 37108 16175 37111
rect 16390 37108 16396 37120
rect 16163 37080 16396 37108
rect 16163 37077 16175 37080
rect 16117 37071 16175 37077
rect 16390 37068 16396 37080
rect 16448 37068 16454 37120
rect 17310 37068 17316 37120
rect 17368 37068 17374 37120
rect 18506 37068 18512 37120
rect 18564 37068 18570 37120
rect 19352 37108 19380 37148
rect 19426 37136 19432 37188
rect 19484 37136 19490 37188
rect 20162 37136 20168 37188
rect 20220 37136 20226 37188
rect 20806 37136 20812 37188
rect 20864 37176 20870 37188
rect 21174 37176 21180 37188
rect 20864 37148 21180 37176
rect 20864 37136 20870 37148
rect 21174 37136 21180 37148
rect 21232 37176 21238 37188
rect 22066 37176 22094 37216
rect 21232 37148 22094 37176
rect 22281 37179 22339 37185
rect 21232 37136 21238 37148
rect 22281 37145 22293 37179
rect 22327 37176 22339 37179
rect 22830 37176 22836 37188
rect 22327 37148 22836 37176
rect 22327 37145 22339 37148
rect 22281 37139 22339 37145
rect 22830 37136 22836 37148
rect 22888 37136 22894 37188
rect 20070 37108 20076 37120
rect 19352 37080 20076 37108
rect 20070 37068 20076 37080
rect 20128 37068 20134 37120
rect 23845 37111 23903 37117
rect 23845 37077 23857 37111
rect 23891 37108 23903 37111
rect 23934 37108 23940 37120
rect 23891 37080 23940 37108
rect 23891 37077 23903 37080
rect 23845 37071 23903 37077
rect 23934 37068 23940 37080
rect 23992 37068 23998 37120
rect 24044 37108 24072 37216
rect 25314 37204 25320 37256
rect 25372 37204 25378 37256
rect 24213 37179 24271 37185
rect 24213 37145 24225 37179
rect 24259 37176 24271 37179
rect 24259 37148 25360 37176
rect 24259 37145 24271 37148
rect 24213 37139 24271 37145
rect 25332 37120 25360 37148
rect 25133 37111 25191 37117
rect 25133 37108 25145 37111
rect 24044 37080 25145 37108
rect 25133 37077 25145 37080
rect 25179 37077 25191 37111
rect 25133 37071 25191 37077
rect 25314 37068 25320 37120
rect 25372 37068 25378 37120
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 5534 36904 5540 36916
rect 3988 36876 5540 36904
rect 3988 36777 4016 36876
rect 5534 36864 5540 36876
rect 5592 36904 5598 36916
rect 6546 36904 6552 36916
rect 5592 36876 6552 36904
rect 5592 36864 5598 36876
rect 6546 36864 6552 36876
rect 6604 36864 6610 36916
rect 7466 36864 7472 36916
rect 7524 36864 7530 36916
rect 7929 36907 7987 36913
rect 7929 36873 7941 36907
rect 7975 36904 7987 36907
rect 8478 36904 8484 36916
rect 7975 36876 8484 36904
rect 7975 36873 7987 36876
rect 7929 36867 7987 36873
rect 8478 36864 8484 36876
rect 8536 36864 8542 36916
rect 9030 36864 9036 36916
rect 9088 36864 9094 36916
rect 12069 36907 12127 36913
rect 12069 36873 12081 36907
rect 12115 36904 12127 36907
rect 12529 36907 12587 36913
rect 12529 36904 12541 36907
rect 12115 36876 12541 36904
rect 12115 36873 12127 36876
rect 12069 36867 12127 36873
rect 12529 36873 12541 36876
rect 12575 36904 12587 36907
rect 12710 36904 12716 36916
rect 12575 36876 12716 36904
rect 12575 36873 12587 36876
rect 12529 36867 12587 36873
rect 12710 36864 12716 36876
rect 12768 36904 12774 36916
rect 13538 36904 13544 36916
rect 12768 36876 13544 36904
rect 12768 36864 12774 36876
rect 13538 36864 13544 36876
rect 13596 36864 13602 36916
rect 13817 36907 13875 36913
rect 13817 36873 13829 36907
rect 13863 36904 13875 36907
rect 14182 36904 14188 36916
rect 13863 36876 14188 36904
rect 13863 36873 13875 36876
rect 13817 36867 13875 36873
rect 14182 36864 14188 36876
rect 14240 36864 14246 36916
rect 15013 36907 15071 36913
rect 15013 36873 15025 36907
rect 15059 36904 15071 36907
rect 15102 36904 15108 36916
rect 15059 36876 15108 36904
rect 15059 36873 15071 36876
rect 15013 36867 15071 36873
rect 15102 36864 15108 36876
rect 15160 36864 15166 36916
rect 15194 36864 15200 36916
rect 15252 36904 15258 36916
rect 15565 36907 15623 36913
rect 15565 36904 15577 36907
rect 15252 36876 15577 36904
rect 15252 36864 15258 36876
rect 15565 36873 15577 36876
rect 15611 36873 15623 36907
rect 15565 36867 15623 36873
rect 17034 36864 17040 36916
rect 17092 36864 17098 36916
rect 17405 36907 17463 36913
rect 17405 36873 17417 36907
rect 17451 36904 17463 36907
rect 18506 36904 18512 36916
rect 17451 36876 18512 36904
rect 17451 36873 17463 36876
rect 17405 36867 17463 36873
rect 18506 36864 18512 36876
rect 18564 36864 18570 36916
rect 20349 36907 20407 36913
rect 20349 36873 20361 36907
rect 20395 36904 20407 36907
rect 20438 36904 20444 36916
rect 20395 36876 20444 36904
rect 20395 36873 20407 36876
rect 20349 36867 20407 36873
rect 20438 36864 20444 36876
rect 20496 36864 20502 36916
rect 23934 36864 23940 36916
rect 23992 36904 23998 36916
rect 23992 36876 24440 36904
rect 23992 36864 23998 36876
rect 5626 36836 5632 36848
rect 5474 36808 5632 36836
rect 5626 36796 5632 36808
rect 5684 36836 5690 36848
rect 5997 36839 6055 36845
rect 5997 36836 6009 36839
rect 5684 36808 6009 36836
rect 5684 36796 5690 36808
rect 5997 36805 6009 36808
rect 6043 36836 6055 36839
rect 7558 36836 7564 36848
rect 6043 36808 7564 36836
rect 6043 36805 6055 36808
rect 5997 36799 6055 36805
rect 7558 36796 7564 36808
rect 7616 36796 7622 36848
rect 10229 36839 10287 36845
rect 10229 36805 10241 36839
rect 10275 36836 10287 36839
rect 10410 36836 10416 36848
rect 10275 36808 10416 36836
rect 10275 36805 10287 36808
rect 10229 36799 10287 36805
rect 10410 36796 10416 36808
rect 10468 36836 10474 36848
rect 11517 36839 11575 36845
rect 11517 36836 11529 36839
rect 10468 36808 11529 36836
rect 10468 36796 10474 36808
rect 11517 36805 11529 36808
rect 11563 36805 11575 36839
rect 11517 36799 11575 36805
rect 3973 36771 4031 36777
rect 3973 36737 3985 36771
rect 4019 36737 4031 36771
rect 3973 36731 4031 36737
rect 7834 36728 7840 36780
rect 7892 36728 7898 36780
rect 9306 36728 9312 36780
rect 9364 36768 9370 36780
rect 9401 36771 9459 36777
rect 9401 36768 9413 36771
rect 9364 36740 9413 36768
rect 9364 36728 9370 36740
rect 9401 36737 9413 36740
rect 9447 36737 9459 36771
rect 9401 36731 9459 36737
rect 4249 36703 4307 36709
rect 4249 36669 4261 36703
rect 4295 36700 4307 36703
rect 5258 36700 5264 36712
rect 4295 36672 5264 36700
rect 4295 36669 4307 36672
rect 4249 36663 4307 36669
rect 5258 36660 5264 36672
rect 5316 36700 5322 36712
rect 5721 36703 5779 36709
rect 5316 36672 5672 36700
rect 5316 36660 5322 36672
rect 5644 36632 5672 36672
rect 5721 36669 5733 36703
rect 5767 36700 5779 36703
rect 5810 36700 5816 36712
rect 5767 36672 5816 36700
rect 5767 36669 5779 36672
rect 5721 36663 5779 36669
rect 5810 36660 5816 36672
rect 5868 36660 5874 36712
rect 5994 36660 6000 36712
rect 6052 36700 6058 36712
rect 8021 36703 8079 36709
rect 8021 36700 8033 36703
rect 6052 36672 8033 36700
rect 6052 36660 6058 36672
rect 8021 36669 8033 36672
rect 8067 36669 8079 36703
rect 8021 36663 8079 36669
rect 9493 36703 9551 36709
rect 9493 36669 9505 36703
rect 9539 36669 9551 36703
rect 9493 36663 9551 36669
rect 7374 36632 7380 36644
rect 5644 36604 7380 36632
rect 7374 36592 7380 36604
rect 7432 36592 7438 36644
rect 9398 36592 9404 36644
rect 9456 36632 9462 36644
rect 9508 36632 9536 36663
rect 9582 36660 9588 36712
rect 9640 36660 9646 36712
rect 10962 36660 10968 36712
rect 11020 36660 11026 36712
rect 9456 36604 9536 36632
rect 11532 36632 11560 36799
rect 13078 36796 13084 36848
rect 13136 36836 13142 36848
rect 17310 36836 17316 36848
rect 13136 36808 17316 36836
rect 13136 36796 13142 36808
rect 17310 36796 17316 36808
rect 17368 36796 17374 36848
rect 24412 36836 24440 36876
rect 24670 36836 24676 36848
rect 24334 36808 24676 36836
rect 24670 36796 24676 36808
rect 24728 36796 24734 36848
rect 12066 36728 12072 36780
rect 12124 36768 12130 36780
rect 13725 36771 13783 36777
rect 12124 36740 13400 36768
rect 12124 36728 12130 36740
rect 11882 36660 11888 36712
rect 11940 36700 11946 36712
rect 12621 36703 12679 36709
rect 12621 36700 12633 36703
rect 11940 36672 12633 36700
rect 11940 36660 11946 36672
rect 12621 36669 12633 36672
rect 12667 36669 12679 36703
rect 12621 36663 12679 36669
rect 12802 36660 12808 36712
rect 12860 36660 12866 36712
rect 13372 36700 13400 36740
rect 13725 36737 13737 36771
rect 13771 36768 13783 36771
rect 13906 36768 13912 36780
rect 13771 36740 13912 36768
rect 13771 36737 13783 36740
rect 13725 36731 13783 36737
rect 13906 36728 13912 36740
rect 13964 36728 13970 36780
rect 14921 36771 14979 36777
rect 14921 36737 14933 36771
rect 14967 36768 14979 36771
rect 14967 36740 15884 36768
rect 14967 36737 14979 36740
rect 14921 36731 14979 36737
rect 15856 36712 15884 36740
rect 16666 36728 16672 36780
rect 16724 36768 16730 36780
rect 17497 36771 17555 36777
rect 17497 36768 17509 36771
rect 16724 36740 17509 36768
rect 16724 36728 16730 36740
rect 17497 36737 17509 36740
rect 17543 36737 17555 36771
rect 17497 36731 17555 36737
rect 19794 36728 19800 36780
rect 19852 36768 19858 36780
rect 20441 36771 20499 36777
rect 20441 36768 20453 36771
rect 19852 36740 20453 36768
rect 19852 36728 19858 36740
rect 20441 36737 20453 36740
rect 20487 36768 20499 36771
rect 20993 36771 21051 36777
rect 20993 36768 21005 36771
rect 20487 36740 21005 36768
rect 20487 36737 20499 36740
rect 20441 36731 20499 36737
rect 20993 36737 21005 36740
rect 21039 36737 21051 36771
rect 20993 36731 21051 36737
rect 25314 36728 25320 36780
rect 25372 36728 25378 36780
rect 13998 36700 14004 36712
rect 13372 36672 14004 36700
rect 13998 36660 14004 36672
rect 14056 36660 14062 36712
rect 14550 36660 14556 36712
rect 14608 36700 14614 36712
rect 15194 36700 15200 36712
rect 14608 36672 15200 36700
rect 14608 36660 14614 36672
rect 15194 36660 15200 36672
rect 15252 36660 15258 36712
rect 15838 36660 15844 36712
rect 15896 36660 15902 36712
rect 17678 36660 17684 36712
rect 17736 36660 17742 36712
rect 18506 36660 18512 36712
rect 18564 36700 18570 36712
rect 20533 36703 20591 36709
rect 20533 36700 20545 36703
rect 18564 36672 20545 36700
rect 18564 36660 18570 36672
rect 20533 36669 20545 36672
rect 20579 36669 20591 36703
rect 20533 36663 20591 36669
rect 22830 36660 22836 36712
rect 22888 36660 22894 36712
rect 23109 36703 23167 36709
rect 23109 36700 23121 36703
rect 22940 36672 23121 36700
rect 16022 36632 16028 36644
rect 11532 36604 16028 36632
rect 9456 36592 9462 36604
rect 16022 36592 16028 36604
rect 16080 36632 16086 36644
rect 19337 36635 19395 36641
rect 19337 36632 19349 36635
rect 16080 36604 19349 36632
rect 16080 36592 16086 36604
rect 19337 36601 19349 36604
rect 19383 36632 19395 36635
rect 19426 36632 19432 36644
rect 19383 36604 19432 36632
rect 19383 36601 19395 36604
rect 19337 36595 19395 36601
rect 19426 36592 19432 36604
rect 19484 36592 19490 36644
rect 20438 36592 20444 36644
rect 20496 36632 20502 36644
rect 22462 36632 22468 36644
rect 20496 36604 22468 36632
rect 20496 36592 20502 36604
rect 22462 36592 22468 36604
rect 22520 36632 22526 36644
rect 22940 36632 22968 36672
rect 23109 36669 23121 36672
rect 23155 36700 23167 36703
rect 23566 36700 23572 36712
rect 23155 36672 23572 36700
rect 23155 36669 23167 36672
rect 23109 36663 23167 36669
rect 23566 36660 23572 36672
rect 23624 36660 23630 36712
rect 23842 36660 23848 36712
rect 23900 36700 23906 36712
rect 24581 36703 24639 36709
rect 24581 36700 24593 36703
rect 23900 36672 24593 36700
rect 23900 36660 23906 36672
rect 24581 36669 24593 36672
rect 24627 36669 24639 36703
rect 24581 36663 24639 36669
rect 25133 36635 25191 36641
rect 25133 36632 25145 36635
rect 22520 36604 22968 36632
rect 24136 36604 25145 36632
rect 22520 36592 22526 36604
rect 1489 36567 1547 36573
rect 1489 36533 1501 36567
rect 1535 36564 1547 36567
rect 1578 36564 1584 36576
rect 1535 36536 1584 36564
rect 1535 36533 1547 36536
rect 1489 36527 1547 36533
rect 1578 36524 1584 36536
rect 1636 36524 1642 36576
rect 8662 36524 8668 36576
rect 8720 36524 8726 36576
rect 10870 36524 10876 36576
rect 10928 36564 10934 36576
rect 12161 36567 12219 36573
rect 12161 36564 12173 36567
rect 10928 36536 12173 36564
rect 10928 36524 10934 36536
rect 12161 36533 12173 36536
rect 12207 36533 12219 36567
rect 12161 36527 12219 36533
rect 13357 36567 13415 36573
rect 13357 36533 13369 36567
rect 13403 36564 13415 36567
rect 14274 36564 14280 36576
rect 13403 36536 14280 36564
rect 13403 36533 13415 36536
rect 13357 36527 13415 36533
rect 14274 36524 14280 36536
rect 14332 36524 14338 36576
rect 14550 36524 14556 36576
rect 14608 36524 14614 36576
rect 17218 36524 17224 36576
rect 17276 36564 17282 36576
rect 19981 36567 20039 36573
rect 19981 36564 19993 36567
rect 17276 36536 19993 36564
rect 17276 36524 17282 36536
rect 19981 36533 19993 36536
rect 20027 36533 20039 36567
rect 19981 36527 20039 36533
rect 20070 36524 20076 36576
rect 20128 36564 20134 36576
rect 24136 36564 24164 36604
rect 25133 36601 25145 36604
rect 25179 36601 25191 36635
rect 25133 36595 25191 36601
rect 20128 36536 24164 36564
rect 20128 36524 20134 36536
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 7650 36320 7656 36372
rect 7708 36320 7714 36372
rect 9122 36320 9128 36372
rect 9180 36320 9186 36372
rect 12437 36363 12495 36369
rect 12437 36329 12449 36363
rect 12483 36360 12495 36363
rect 12526 36360 12532 36372
rect 12483 36332 12532 36360
rect 12483 36329 12495 36332
rect 12437 36323 12495 36329
rect 12526 36320 12532 36332
rect 12584 36320 12590 36372
rect 12713 36363 12771 36369
rect 12713 36329 12725 36363
rect 12759 36360 12771 36363
rect 13354 36360 13360 36372
rect 12759 36332 13360 36360
rect 12759 36329 12771 36332
rect 12713 36323 12771 36329
rect 13354 36320 13360 36332
rect 13412 36320 13418 36372
rect 13538 36320 13544 36372
rect 13596 36360 13602 36372
rect 14277 36363 14335 36369
rect 13596 36332 13676 36360
rect 13596 36320 13602 36332
rect 7098 36252 7104 36304
rect 7156 36292 7162 36304
rect 12161 36295 12219 36301
rect 12161 36292 12173 36295
rect 7156 36264 12173 36292
rect 7156 36252 7162 36264
rect 12161 36261 12173 36264
rect 12207 36292 12219 36295
rect 12544 36292 12572 36320
rect 12207 36264 12434 36292
rect 12544 36264 13216 36292
rect 12207 36261 12219 36264
rect 12161 36255 12219 36261
rect 7558 36184 7564 36236
rect 7616 36224 7622 36236
rect 8205 36227 8263 36233
rect 8205 36224 8217 36227
rect 7616 36196 8217 36224
rect 7616 36184 7622 36196
rect 8205 36193 8217 36196
rect 8251 36193 8263 36227
rect 9677 36227 9735 36233
rect 9677 36224 9689 36227
rect 8205 36187 8263 36193
rect 8312 36196 9689 36224
rect 1578 36116 1584 36168
rect 1636 36116 1642 36168
rect 7374 36116 7380 36168
rect 7432 36156 7438 36168
rect 8312 36156 8340 36196
rect 9677 36193 9689 36196
rect 9723 36193 9735 36227
rect 12406 36224 12434 36264
rect 12710 36224 12716 36236
rect 12406 36196 12716 36224
rect 9677 36187 9735 36193
rect 12710 36184 12716 36196
rect 12768 36184 12774 36236
rect 13188 36233 13216 36264
rect 13173 36227 13231 36233
rect 13173 36193 13185 36227
rect 13219 36193 13231 36227
rect 13173 36187 13231 36193
rect 13357 36227 13415 36233
rect 13357 36193 13369 36227
rect 13403 36224 13415 36227
rect 13538 36224 13544 36236
rect 13403 36196 13544 36224
rect 13403 36193 13415 36196
rect 13357 36187 13415 36193
rect 13538 36184 13544 36196
rect 13596 36184 13602 36236
rect 7432 36128 8340 36156
rect 9585 36159 9643 36165
rect 7432 36116 7438 36128
rect 9585 36125 9597 36159
rect 9631 36156 9643 36159
rect 12342 36156 12348 36168
rect 9631 36128 12348 36156
rect 9631 36125 9643 36128
rect 9585 36119 9643 36125
rect 12342 36116 12348 36128
rect 12400 36116 12406 36168
rect 13648 36156 13676 36332
rect 14277 36329 14289 36363
rect 14323 36360 14335 36363
rect 15378 36360 15384 36372
rect 14323 36332 15384 36360
rect 14323 36329 14335 36332
rect 14277 36323 14335 36329
rect 15378 36320 15384 36332
rect 15436 36320 15442 36372
rect 16117 36363 16175 36369
rect 16117 36329 16129 36363
rect 16163 36360 16175 36363
rect 18782 36360 18788 36372
rect 16163 36332 18788 36360
rect 16163 36329 16175 36332
rect 16117 36323 16175 36329
rect 18782 36320 18788 36332
rect 18840 36320 18846 36372
rect 19242 36320 19248 36372
rect 19300 36360 19306 36372
rect 19429 36363 19487 36369
rect 19429 36360 19441 36363
rect 19300 36332 19441 36360
rect 19300 36320 19306 36332
rect 19429 36329 19441 36332
rect 19475 36329 19487 36363
rect 21726 36360 21732 36372
rect 19429 36323 19487 36329
rect 20088 36332 21732 36360
rect 13814 36252 13820 36304
rect 13872 36292 13878 36304
rect 13872 36264 14780 36292
rect 13872 36252 13878 36264
rect 14752 36233 14780 36264
rect 16942 36252 16948 36304
rect 17000 36292 17006 36304
rect 19061 36295 19119 36301
rect 19061 36292 19073 36295
rect 17000 36264 19073 36292
rect 17000 36252 17006 36264
rect 19061 36261 19073 36264
rect 19107 36292 19119 36295
rect 19107 36264 20024 36292
rect 19107 36261 19119 36264
rect 19061 36255 19119 36261
rect 14737 36227 14795 36233
rect 14737 36193 14749 36227
rect 14783 36193 14795 36227
rect 14737 36187 14795 36193
rect 14921 36227 14979 36233
rect 14921 36193 14933 36227
rect 14967 36224 14979 36227
rect 15654 36224 15660 36236
rect 14967 36196 15660 36224
rect 14967 36193 14979 36196
rect 14921 36187 14979 36193
rect 15654 36184 15660 36196
rect 15712 36184 15718 36236
rect 16761 36227 16819 36233
rect 16761 36193 16773 36227
rect 16807 36224 16819 36227
rect 19702 36224 19708 36236
rect 16807 36196 19708 36224
rect 16807 36193 16819 36196
rect 16761 36187 16819 36193
rect 19702 36184 19708 36196
rect 19760 36184 19766 36236
rect 19996 36233 20024 36264
rect 19981 36227 20039 36233
rect 19981 36193 19993 36227
rect 20027 36193 20039 36227
rect 19981 36187 20039 36193
rect 16577 36159 16635 36165
rect 16577 36156 16589 36159
rect 13648 36128 14780 36156
rect 8113 36091 8171 36097
rect 8113 36057 8125 36091
rect 8159 36088 8171 36091
rect 10410 36088 10416 36100
rect 8159 36060 10416 36088
rect 8159 36057 8171 36060
rect 8113 36051 8171 36057
rect 10410 36048 10416 36060
rect 10468 36048 10474 36100
rect 1762 35980 1768 36032
rect 1820 36020 1826 36032
rect 2225 36023 2283 36029
rect 2225 36020 2237 36023
rect 1820 35992 2237 36020
rect 1820 35980 1826 35992
rect 2225 35989 2237 35992
rect 2271 35989 2283 36023
rect 2225 35983 2283 35989
rect 7466 35980 7472 36032
rect 7524 36020 7530 36032
rect 8021 36023 8079 36029
rect 8021 36020 8033 36023
rect 7524 35992 8033 36020
rect 7524 35980 7530 35992
rect 8021 35989 8033 35992
rect 8067 35989 8079 36023
rect 8021 35983 8079 35989
rect 9493 36023 9551 36029
rect 9493 35989 9505 36023
rect 9539 36020 9551 36023
rect 11330 36020 11336 36032
rect 9539 35992 11336 36020
rect 9539 35989 9551 35992
rect 9493 35983 9551 35989
rect 11330 35980 11336 35992
rect 11388 35980 11394 36032
rect 12710 35980 12716 36032
rect 12768 36020 12774 36032
rect 13081 36023 13139 36029
rect 13081 36020 13093 36023
rect 12768 35992 13093 36020
rect 12768 35980 12774 35992
rect 13081 35989 13093 35992
rect 13127 35989 13139 36023
rect 13081 35983 13139 35989
rect 14642 35980 14648 36032
rect 14700 35980 14706 36032
rect 14752 36020 14780 36128
rect 15764 36128 16589 36156
rect 15654 36048 15660 36100
rect 15712 36088 15718 36100
rect 15764 36097 15792 36128
rect 16577 36125 16589 36128
rect 16623 36125 16635 36159
rect 20088 36156 20116 36332
rect 21726 36320 21732 36332
rect 21784 36360 21790 36372
rect 21784 36332 22094 36360
rect 21784 36320 21790 36332
rect 20346 36184 20352 36236
rect 20404 36224 20410 36236
rect 21269 36227 21327 36233
rect 21269 36224 21281 36227
rect 20404 36196 21281 36224
rect 20404 36184 20410 36196
rect 21269 36193 21281 36196
rect 21315 36193 21327 36227
rect 21269 36187 21327 36193
rect 21358 36184 21364 36236
rect 21416 36184 21422 36236
rect 16577 36119 16635 36125
rect 17420 36128 20116 36156
rect 15749 36091 15807 36097
rect 15749 36088 15761 36091
rect 15712 36060 15761 36088
rect 15712 36048 15718 36060
rect 15749 36057 15761 36060
rect 15795 36057 15807 36091
rect 15749 36051 15807 36057
rect 16485 36091 16543 36097
rect 16485 36057 16497 36091
rect 16531 36088 16543 36091
rect 17313 36091 17371 36097
rect 17313 36088 17325 36091
rect 16531 36060 17325 36088
rect 16531 36057 16543 36060
rect 16485 36051 16543 36057
rect 17313 36057 17325 36060
rect 17359 36057 17371 36091
rect 17313 36051 17371 36057
rect 17420 36020 17448 36128
rect 20898 36116 20904 36168
rect 20956 36156 20962 36168
rect 21177 36159 21235 36165
rect 21177 36156 21189 36159
rect 20956 36128 21189 36156
rect 20956 36116 20962 36128
rect 21177 36125 21189 36128
rect 21223 36125 21235 36159
rect 22066 36156 22094 36332
rect 23198 36320 23204 36372
rect 23256 36360 23262 36372
rect 25130 36360 25136 36372
rect 23256 36332 25136 36360
rect 23256 36320 23262 36332
rect 25130 36320 25136 36332
rect 25188 36320 25194 36372
rect 23293 36295 23351 36301
rect 23293 36261 23305 36295
rect 23339 36292 23351 36295
rect 24394 36292 24400 36304
rect 23339 36264 24400 36292
rect 23339 36261 23351 36264
rect 23293 36255 23351 36261
rect 24394 36252 24400 36264
rect 24452 36252 24458 36304
rect 23750 36184 23756 36236
rect 23808 36184 23814 36236
rect 23937 36227 23995 36233
rect 23937 36193 23949 36227
rect 23983 36224 23995 36227
rect 24486 36224 24492 36236
rect 23983 36196 24492 36224
rect 23983 36193 23995 36196
rect 23937 36187 23995 36193
rect 24486 36184 24492 36196
rect 24544 36184 24550 36236
rect 24118 36156 24124 36168
rect 22066 36128 24124 36156
rect 21177 36119 21235 36125
rect 24118 36116 24124 36128
rect 24176 36116 24182 36168
rect 24857 36159 24915 36165
rect 24857 36125 24869 36159
rect 24903 36156 24915 36159
rect 25314 36156 25320 36168
rect 24903 36128 25320 36156
rect 24903 36125 24915 36128
rect 24857 36119 24915 36125
rect 25314 36116 25320 36128
rect 25372 36116 25378 36168
rect 19889 36091 19947 36097
rect 19889 36057 19901 36091
rect 19935 36088 19947 36091
rect 19935 36060 21404 36088
rect 19935 36057 19947 36060
rect 19889 36051 19947 36057
rect 14752 35992 17448 36020
rect 19610 35980 19616 36032
rect 19668 36020 19674 36032
rect 19797 36023 19855 36029
rect 19797 36020 19809 36023
rect 19668 35992 19809 36020
rect 19668 35980 19674 35992
rect 19797 35989 19809 35992
rect 19843 35989 19855 36023
rect 19797 35983 19855 35989
rect 20809 36023 20867 36029
rect 20809 35989 20821 36023
rect 20855 36020 20867 36023
rect 20898 36020 20904 36032
rect 20855 35992 20904 36020
rect 20855 35989 20867 35992
rect 20809 35983 20867 35989
rect 20898 35980 20904 35992
rect 20956 35980 20962 36032
rect 21376 36020 21404 36060
rect 21818 36048 21824 36100
rect 21876 36088 21882 36100
rect 21876 36060 25176 36088
rect 21876 36048 21882 36060
rect 22278 36020 22284 36032
rect 21376 35992 22284 36020
rect 22278 35980 22284 35992
rect 22336 36020 22342 36032
rect 23198 36020 23204 36032
rect 22336 35992 23204 36020
rect 22336 35980 22342 35992
rect 23198 35980 23204 35992
rect 23256 35980 23262 36032
rect 23658 35980 23664 36032
rect 23716 35980 23722 36032
rect 25148 36029 25176 36060
rect 25133 36023 25191 36029
rect 25133 35989 25145 36023
rect 25179 35989 25191 36023
rect 25133 35983 25191 35989
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 5534 35816 5540 35828
rect 4264 35788 5540 35816
rect 1762 35640 1768 35692
rect 1820 35640 1826 35692
rect 4264 35689 4292 35788
rect 5534 35776 5540 35788
rect 5592 35776 5598 35828
rect 5994 35776 6000 35828
rect 6052 35776 6058 35828
rect 7282 35776 7288 35828
rect 7340 35816 7346 35828
rect 8570 35816 8576 35828
rect 7340 35788 8576 35816
rect 7340 35776 7346 35788
rect 8570 35776 8576 35788
rect 8628 35776 8634 35828
rect 10226 35816 10232 35828
rect 8772 35788 10232 35816
rect 8772 35748 8800 35788
rect 10226 35776 10232 35788
rect 10284 35776 10290 35828
rect 13446 35816 13452 35828
rect 10612 35788 13452 35816
rect 6932 35720 8878 35748
rect 6932 35692 6960 35720
rect 4249 35683 4307 35689
rect 4249 35649 4261 35683
rect 4295 35649 4307 35683
rect 4249 35643 4307 35649
rect 5626 35640 5632 35692
rect 5684 35680 5690 35692
rect 6365 35683 6423 35689
rect 6365 35680 6377 35683
rect 5684 35652 6377 35680
rect 5684 35640 5690 35652
rect 6365 35649 6377 35652
rect 6411 35680 6423 35683
rect 6914 35680 6920 35692
rect 6411 35652 6920 35680
rect 6411 35649 6423 35652
rect 6365 35643 6423 35649
rect 6914 35640 6920 35652
rect 6972 35640 6978 35692
rect 10612 35680 10640 35788
rect 13446 35776 13452 35788
rect 13504 35776 13510 35828
rect 13538 35776 13544 35828
rect 13596 35816 13602 35828
rect 13909 35819 13967 35825
rect 13909 35816 13921 35819
rect 13596 35788 13921 35816
rect 13596 35776 13602 35788
rect 13909 35785 13921 35788
rect 13955 35785 13967 35819
rect 13909 35779 13967 35785
rect 14461 35819 14519 35825
rect 14461 35785 14473 35819
rect 14507 35816 14519 35819
rect 14642 35816 14648 35828
rect 14507 35788 14648 35816
rect 14507 35785 14519 35788
rect 14461 35779 14519 35785
rect 13924 35748 13952 35779
rect 14642 35776 14648 35788
rect 14700 35776 14706 35828
rect 17586 35776 17592 35828
rect 17644 35816 17650 35828
rect 20165 35819 20223 35825
rect 20165 35816 20177 35819
rect 17644 35788 20177 35816
rect 17644 35776 17650 35788
rect 20165 35785 20177 35788
rect 20211 35816 20223 35819
rect 20211 35788 21680 35816
rect 20211 35785 20223 35788
rect 20165 35779 20223 35785
rect 17402 35748 17408 35760
rect 13924 35720 17408 35748
rect 17402 35708 17408 35720
rect 17460 35708 17466 35760
rect 17770 35708 17776 35760
rect 17828 35748 17834 35760
rect 17865 35751 17923 35757
rect 17865 35748 17877 35751
rect 17828 35720 17877 35748
rect 17828 35708 17834 35720
rect 17865 35717 17877 35720
rect 17911 35717 17923 35751
rect 17865 35711 17923 35717
rect 18322 35708 18328 35760
rect 18380 35708 18386 35760
rect 19978 35708 19984 35760
rect 20036 35748 20042 35760
rect 20257 35751 20315 35757
rect 20257 35748 20269 35751
rect 20036 35720 20269 35748
rect 20036 35708 20042 35720
rect 20257 35717 20269 35720
rect 20303 35717 20315 35751
rect 20257 35711 20315 35717
rect 21542 35680 21548 35692
rect 9876 35652 10640 35680
rect 13110 35652 13860 35680
rect 4525 35615 4583 35621
rect 4525 35581 4537 35615
rect 4571 35612 4583 35615
rect 5810 35612 5816 35624
rect 4571 35584 5816 35612
rect 4571 35581 4583 35584
rect 4525 35575 4583 35581
rect 5810 35572 5816 35584
rect 5868 35572 5874 35624
rect 8113 35615 8171 35621
rect 8113 35581 8125 35615
rect 8159 35581 8171 35615
rect 8113 35575 8171 35581
rect 8389 35615 8447 35621
rect 8389 35581 8401 35615
rect 8435 35612 8447 35615
rect 9582 35612 9588 35624
rect 8435 35584 9588 35612
rect 8435 35581 8447 35584
rect 8389 35575 8447 35581
rect 1581 35479 1639 35485
rect 1581 35445 1593 35479
rect 1627 35476 1639 35479
rect 4062 35476 4068 35488
rect 1627 35448 4068 35476
rect 1627 35445 1639 35448
rect 1581 35439 1639 35445
rect 4062 35436 4068 35448
rect 4120 35436 4126 35488
rect 8128 35476 8156 35575
rect 9582 35572 9588 35584
rect 9640 35572 9646 35624
rect 8570 35476 8576 35488
rect 8128 35448 8576 35476
rect 8570 35436 8576 35448
rect 8628 35436 8634 35488
rect 9766 35436 9772 35488
rect 9824 35476 9830 35488
rect 9876 35485 9904 35652
rect 10962 35572 10968 35624
rect 11020 35612 11026 35624
rect 11701 35615 11759 35621
rect 11701 35612 11713 35615
rect 11020 35584 11713 35612
rect 11020 35572 11026 35584
rect 11701 35581 11713 35584
rect 11747 35581 11759 35615
rect 11701 35575 11759 35581
rect 11974 35572 11980 35624
rect 12032 35572 12038 35624
rect 9861 35479 9919 35485
rect 9861 35476 9873 35479
rect 9824 35448 9873 35476
rect 9824 35436 9830 35448
rect 9861 35445 9873 35448
rect 9907 35445 9919 35479
rect 9861 35439 9919 35445
rect 10226 35436 10232 35488
rect 10284 35476 10290 35488
rect 10778 35476 10784 35488
rect 10284 35448 10784 35476
rect 10284 35436 10290 35448
rect 10778 35436 10784 35448
rect 10836 35436 10842 35488
rect 11698 35436 11704 35488
rect 11756 35476 11762 35488
rect 13449 35479 13507 35485
rect 13449 35476 13461 35479
rect 11756 35448 13461 35476
rect 11756 35436 11762 35448
rect 13449 35445 13461 35448
rect 13495 35476 13507 35479
rect 13630 35476 13636 35488
rect 13495 35448 13636 35476
rect 13495 35445 13507 35448
rect 13449 35439 13507 35445
rect 13630 35436 13636 35448
rect 13688 35436 13694 35488
rect 13832 35485 13860 35652
rect 19352 35652 21548 35680
rect 15194 35572 15200 35624
rect 15252 35612 15258 35624
rect 17402 35612 17408 35624
rect 15252 35584 17408 35612
rect 15252 35572 15258 35584
rect 17402 35572 17408 35584
rect 17460 35572 17466 35624
rect 19352 35621 19380 35652
rect 21542 35640 21548 35652
rect 21600 35640 21606 35692
rect 17589 35615 17647 35621
rect 17589 35581 17601 35615
rect 17635 35581 17647 35615
rect 17589 35575 17647 35581
rect 19337 35615 19395 35621
rect 19337 35581 19349 35615
rect 19383 35581 19395 35615
rect 19337 35575 19395 35581
rect 20349 35615 20407 35621
rect 20349 35581 20361 35615
rect 20395 35581 20407 35615
rect 20349 35575 20407 35581
rect 13817 35479 13875 35485
rect 13817 35445 13829 35479
rect 13863 35476 13875 35479
rect 13906 35476 13912 35488
rect 13863 35448 13912 35476
rect 13863 35445 13875 35448
rect 13817 35439 13875 35445
rect 13906 35436 13912 35448
rect 13964 35436 13970 35488
rect 15930 35436 15936 35488
rect 15988 35476 15994 35488
rect 17604 35476 17632 35575
rect 19150 35504 19156 35556
rect 19208 35544 19214 35556
rect 19208 35516 20116 35544
rect 19208 35504 19214 35516
rect 17954 35476 17960 35488
rect 15988 35448 17960 35476
rect 15988 35436 15994 35448
rect 17954 35436 17960 35448
rect 18012 35436 18018 35488
rect 19794 35436 19800 35488
rect 19852 35436 19858 35488
rect 20088 35476 20116 35516
rect 20364 35476 20392 35575
rect 21652 35544 21680 35788
rect 22186 35776 22192 35828
rect 22244 35776 22250 35828
rect 23566 35776 23572 35828
rect 23624 35816 23630 35828
rect 24857 35819 24915 35825
rect 24857 35816 24869 35819
rect 23624 35788 24869 35816
rect 23624 35776 23630 35788
rect 24857 35785 24869 35788
rect 24903 35785 24915 35819
rect 24857 35779 24915 35785
rect 22204 35748 22232 35776
rect 24670 35748 24676 35760
rect 22112 35720 22232 35748
rect 24610 35720 24676 35748
rect 22112 35692 22140 35720
rect 24670 35708 24676 35720
rect 24728 35748 24734 35760
rect 25222 35748 25228 35760
rect 24728 35720 25228 35748
rect 24728 35708 24734 35720
rect 25222 35708 25228 35720
rect 25280 35708 25286 35760
rect 22094 35640 22100 35692
rect 22152 35640 22158 35692
rect 22186 35640 22192 35692
rect 22244 35680 22250 35692
rect 22830 35680 22836 35692
rect 22244 35652 22836 35680
rect 22244 35640 22250 35652
rect 22830 35640 22836 35652
rect 22888 35680 22894 35692
rect 23109 35683 23167 35689
rect 23109 35680 23121 35683
rect 22888 35652 23121 35680
rect 22888 35640 22894 35652
rect 23109 35649 23121 35652
rect 23155 35649 23167 35683
rect 23109 35643 23167 35649
rect 22462 35572 22468 35624
rect 22520 35572 22526 35624
rect 23382 35572 23388 35624
rect 23440 35572 23446 35624
rect 22370 35544 22376 35556
rect 21652 35516 22376 35544
rect 22370 35504 22376 35516
rect 22428 35504 22434 35556
rect 22554 35504 22560 35556
rect 22612 35544 22618 35556
rect 22830 35544 22836 35556
rect 22612 35516 22836 35544
rect 22612 35504 22618 35516
rect 22830 35504 22836 35516
rect 22888 35504 22894 35556
rect 20088 35448 20392 35476
rect 20714 35436 20720 35488
rect 20772 35476 20778 35488
rect 20809 35479 20867 35485
rect 20809 35476 20821 35479
rect 20772 35448 20821 35476
rect 20772 35436 20778 35448
rect 20809 35445 20821 35448
rect 20855 35445 20867 35479
rect 20809 35439 20867 35445
rect 25222 35436 25228 35488
rect 25280 35436 25286 35488
rect 25314 35436 25320 35488
rect 25372 35476 25378 35488
rect 25409 35479 25467 35485
rect 25409 35476 25421 35479
rect 25372 35448 25421 35476
rect 25372 35436 25378 35448
rect 25409 35445 25421 35448
rect 25455 35445 25467 35479
rect 25409 35439 25467 35445
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 7374 35232 7380 35284
rect 7432 35272 7438 35284
rect 7837 35275 7895 35281
rect 7837 35272 7849 35275
rect 7432 35244 7849 35272
rect 7432 35232 7438 35244
rect 7837 35241 7849 35244
rect 7883 35241 7895 35275
rect 7837 35235 7895 35241
rect 8754 35232 8760 35284
rect 8812 35272 8818 35284
rect 9309 35275 9367 35281
rect 9309 35272 9321 35275
rect 8812 35244 9321 35272
rect 8812 35232 8818 35244
rect 9309 35241 9321 35244
rect 9355 35241 9367 35275
rect 9309 35235 9367 35241
rect 9398 35232 9404 35284
rect 9456 35272 9462 35284
rect 12989 35275 13047 35281
rect 12989 35272 13001 35275
rect 9456 35244 13001 35272
rect 9456 35232 9462 35244
rect 12989 35241 13001 35244
rect 13035 35241 13047 35275
rect 12989 35235 13047 35241
rect 16114 35232 16120 35284
rect 16172 35272 16178 35284
rect 17129 35275 17187 35281
rect 17129 35272 17141 35275
rect 16172 35244 17141 35272
rect 16172 35232 16178 35244
rect 17129 35241 17141 35244
rect 17175 35241 17187 35275
rect 17129 35235 17187 35241
rect 17497 35275 17555 35281
rect 17497 35241 17509 35275
rect 17543 35272 17555 35275
rect 18322 35272 18328 35284
rect 17543 35244 18328 35272
rect 17543 35241 17555 35244
rect 17497 35235 17555 35241
rect 11974 35164 11980 35216
rect 12032 35204 12038 35216
rect 13814 35204 13820 35216
rect 12032 35176 13820 35204
rect 12032 35164 12038 35176
rect 13814 35164 13820 35176
rect 13872 35164 13878 35216
rect 5534 35096 5540 35148
rect 5592 35136 5598 35148
rect 6086 35136 6092 35148
rect 5592 35108 6092 35136
rect 5592 35096 5598 35108
rect 6086 35096 6092 35108
rect 6144 35096 6150 35148
rect 6365 35139 6423 35145
rect 6365 35105 6377 35139
rect 6411 35136 6423 35139
rect 9766 35136 9772 35148
rect 6411 35108 9772 35136
rect 6411 35105 6423 35108
rect 6365 35099 6423 35105
rect 9766 35096 9772 35108
rect 9824 35096 9830 35148
rect 9858 35096 9864 35148
rect 9916 35096 9922 35148
rect 11146 35096 11152 35148
rect 11204 35136 11210 35148
rect 13541 35139 13599 35145
rect 13541 35136 13553 35139
rect 11204 35108 13553 35136
rect 11204 35096 11210 35108
rect 13541 35105 13553 35108
rect 13587 35105 13599 35139
rect 13541 35099 13599 35105
rect 15381 35139 15439 35145
rect 15381 35105 15393 35139
rect 15427 35136 15439 35139
rect 15746 35136 15752 35148
rect 15427 35108 15752 35136
rect 15427 35105 15439 35108
rect 15381 35099 15439 35105
rect 15746 35096 15752 35108
rect 15804 35096 15810 35148
rect 13449 35071 13507 35077
rect 13449 35037 13461 35071
rect 13495 35068 13507 35071
rect 14550 35068 14556 35080
rect 13495 35040 14556 35068
rect 13495 35037 13507 35040
rect 13449 35031 13507 35037
rect 14550 35028 14556 35040
rect 14608 35028 14614 35080
rect 17512 35068 17540 35235
rect 18322 35232 18328 35244
rect 18380 35232 18386 35284
rect 19702 35232 19708 35284
rect 19760 35272 19766 35284
rect 20346 35272 20352 35284
rect 19760 35244 20352 35272
rect 19760 35232 19766 35244
rect 20346 35232 20352 35244
rect 20404 35232 20410 35284
rect 21634 35232 21640 35284
rect 21692 35232 21698 35284
rect 20714 35164 20720 35216
rect 20772 35204 20778 35216
rect 21729 35207 21787 35213
rect 21729 35204 21741 35207
rect 20772 35176 21741 35204
rect 20772 35164 20778 35176
rect 21729 35173 21741 35176
rect 21775 35204 21787 35207
rect 21775 35176 22094 35204
rect 21775 35173 21787 35176
rect 21729 35167 21787 35173
rect 17954 35096 17960 35148
rect 18012 35136 18018 35148
rect 18322 35136 18328 35148
rect 18012 35108 18328 35136
rect 18012 35096 18018 35108
rect 18322 35096 18328 35108
rect 18380 35136 18386 35148
rect 19429 35139 19487 35145
rect 19429 35136 19441 35139
rect 18380 35108 19441 35136
rect 18380 35096 18386 35108
rect 19429 35105 19441 35108
rect 19475 35136 19487 35139
rect 20162 35136 20168 35148
rect 19475 35108 20168 35136
rect 19475 35105 19487 35108
rect 19429 35099 19487 35105
rect 20162 35096 20168 35108
rect 20220 35096 20226 35148
rect 22066 35136 22094 35176
rect 22066 35108 23796 35136
rect 16790 35040 17540 35068
rect 22186 35028 22192 35080
rect 22244 35068 22250 35080
rect 22281 35071 22339 35077
rect 22281 35068 22293 35071
rect 22244 35040 22293 35068
rect 22244 35028 22250 35040
rect 22281 35037 22293 35040
rect 22327 35037 22339 35071
rect 22281 35031 22339 35037
rect 6914 34960 6920 35012
rect 6972 34960 6978 35012
rect 8662 34960 8668 35012
rect 8720 35000 8726 35012
rect 9677 35003 9735 35009
rect 9677 35000 9689 35003
rect 8720 34972 9689 35000
rect 8720 34960 8726 34972
rect 9677 34969 9689 34972
rect 9723 34969 9735 35003
rect 9677 34963 9735 34969
rect 9769 35003 9827 35009
rect 9769 34969 9781 35003
rect 9815 35000 9827 35003
rect 14182 35000 14188 35012
rect 9815 34972 14188 35000
rect 9815 34969 9827 34972
rect 9769 34963 9827 34969
rect 14182 34960 14188 34972
rect 14240 34960 14246 35012
rect 15657 35003 15715 35009
rect 15657 34969 15669 35003
rect 15703 34969 15715 35003
rect 15657 34963 15715 34969
rect 17052 34972 19656 35000
rect 7006 34892 7012 34944
rect 7064 34932 7070 34944
rect 8113 34935 8171 34941
rect 8113 34932 8125 34935
rect 7064 34904 8125 34932
rect 7064 34892 7070 34904
rect 8113 34901 8125 34904
rect 8159 34901 8171 34935
rect 8113 34895 8171 34901
rect 8294 34892 8300 34944
rect 8352 34932 8358 34944
rect 10686 34932 10692 34944
rect 8352 34904 10692 34932
rect 8352 34892 8358 34904
rect 10686 34892 10692 34904
rect 10744 34892 10750 34944
rect 13354 34892 13360 34944
rect 13412 34892 13418 34944
rect 15672 34932 15700 34963
rect 17052 34932 17080 34972
rect 15672 34904 17080 34932
rect 19628 34932 19656 34972
rect 19702 34960 19708 35012
rect 19760 35000 19766 35012
rect 19760 34972 20024 35000
rect 19760 34960 19766 34972
rect 19886 34932 19892 34944
rect 19628 34904 19892 34932
rect 19886 34892 19892 34904
rect 19944 34892 19950 34944
rect 19996 34932 20024 34972
rect 20714 34960 20720 35012
rect 20772 34960 20778 35012
rect 21266 34960 21272 35012
rect 21324 35000 21330 35012
rect 22557 35003 22615 35009
rect 22557 35000 22569 35003
rect 21324 34972 22569 35000
rect 21324 34960 21330 34972
rect 22557 34969 22569 34972
rect 22603 35000 22615 35003
rect 22646 35000 22652 35012
rect 22603 34972 22652 35000
rect 22603 34969 22615 34972
rect 22557 34963 22615 34969
rect 22646 34960 22652 34972
rect 22704 34960 22710 35012
rect 23768 35000 23796 35108
rect 25314 35028 25320 35080
rect 25372 35028 25378 35080
rect 25222 35000 25228 35012
rect 23768 34986 25228 35000
rect 23782 34972 25228 34986
rect 24320 34944 24348 34972
rect 25222 34960 25228 34972
rect 25280 34960 25286 35012
rect 20990 34932 20996 34944
rect 19996 34904 20996 34932
rect 20990 34892 20996 34904
rect 21048 34892 21054 34944
rect 21177 34935 21235 34941
rect 21177 34901 21189 34935
rect 21223 34932 21235 34935
rect 21358 34932 21364 34944
rect 21223 34904 21364 34932
rect 21223 34901 21235 34904
rect 21177 34895 21235 34901
rect 21358 34892 21364 34904
rect 21416 34892 21422 34944
rect 22370 34892 22376 34944
rect 22428 34932 22434 34944
rect 23198 34932 23204 34944
rect 22428 34904 23204 34932
rect 22428 34892 22434 34904
rect 23198 34892 23204 34904
rect 23256 34892 23262 34944
rect 23382 34892 23388 34944
rect 23440 34932 23446 34944
rect 24029 34935 24087 34941
rect 24029 34932 24041 34935
rect 23440 34904 24041 34932
rect 23440 34892 23446 34904
rect 24029 34901 24041 34904
rect 24075 34901 24087 34935
rect 24029 34895 24087 34901
rect 24302 34892 24308 34944
rect 24360 34932 24366 34944
rect 24397 34935 24455 34941
rect 24397 34932 24409 34935
rect 24360 34904 24409 34932
rect 24360 34892 24366 34904
rect 24397 34901 24409 34904
rect 24443 34901 24455 34935
rect 24397 34895 24455 34901
rect 24486 34892 24492 34944
rect 24544 34932 24550 34944
rect 25133 34935 25191 34941
rect 25133 34932 25145 34935
rect 24544 34904 25145 34932
rect 24544 34892 24550 34904
rect 25133 34901 25145 34904
rect 25179 34901 25191 34935
rect 25133 34895 25191 34901
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 7190 34688 7196 34740
rect 7248 34728 7254 34740
rect 8294 34728 8300 34740
rect 7248 34700 8300 34728
rect 7248 34688 7254 34700
rect 8294 34688 8300 34700
rect 8352 34688 8358 34740
rect 9490 34688 9496 34740
rect 9548 34728 9554 34740
rect 10597 34731 10655 34737
rect 10597 34728 10609 34731
rect 9548 34700 10609 34728
rect 9548 34688 9554 34700
rect 10597 34697 10609 34700
rect 10643 34697 10655 34731
rect 10597 34691 10655 34697
rect 10686 34688 10692 34740
rect 10744 34728 10750 34740
rect 12802 34728 12808 34740
rect 10744 34700 12808 34728
rect 10744 34688 10750 34700
rect 12802 34688 12808 34700
rect 12860 34728 12866 34740
rect 13722 34728 13728 34740
rect 12860 34700 13728 34728
rect 12860 34688 12866 34700
rect 13722 34688 13728 34700
rect 13780 34688 13786 34740
rect 15933 34731 15991 34737
rect 15933 34697 15945 34731
rect 15979 34728 15991 34731
rect 19794 34728 19800 34740
rect 15979 34700 19800 34728
rect 15979 34697 15991 34700
rect 15933 34691 15991 34697
rect 19794 34688 19800 34700
rect 19852 34688 19858 34740
rect 20254 34688 20260 34740
rect 20312 34688 20318 34740
rect 20717 34731 20775 34737
rect 20717 34697 20729 34731
rect 20763 34728 20775 34731
rect 20806 34728 20812 34740
rect 20763 34700 20812 34728
rect 20763 34697 20775 34700
rect 20717 34691 20775 34697
rect 20806 34688 20812 34700
rect 20864 34688 20870 34740
rect 21085 34731 21143 34737
rect 21085 34697 21097 34731
rect 21131 34728 21143 34731
rect 21174 34728 21180 34740
rect 21131 34700 21180 34728
rect 21131 34697 21143 34700
rect 21085 34691 21143 34697
rect 21174 34688 21180 34700
rect 21232 34688 21238 34740
rect 22278 34688 22284 34740
rect 22336 34728 22342 34740
rect 22373 34731 22431 34737
rect 22373 34728 22385 34731
rect 22336 34700 22385 34728
rect 22336 34688 22342 34700
rect 22373 34697 22385 34700
rect 22419 34697 22431 34731
rect 22373 34691 22431 34697
rect 23201 34731 23259 34737
rect 23201 34697 23213 34731
rect 23247 34728 23259 34731
rect 23658 34728 23664 34740
rect 23247 34700 23664 34728
rect 23247 34697 23259 34700
rect 23201 34691 23259 34697
rect 23658 34688 23664 34700
rect 23716 34688 23722 34740
rect 24397 34731 24455 34737
rect 24397 34697 24409 34731
rect 24443 34728 24455 34731
rect 24670 34728 24676 34740
rect 24443 34700 24676 34728
rect 24443 34697 24455 34700
rect 24397 34691 24455 34697
rect 24670 34688 24676 34700
rect 24728 34688 24734 34740
rect 5994 34620 6000 34672
rect 6052 34660 6058 34672
rect 6825 34663 6883 34669
rect 6825 34660 6837 34663
rect 6052 34632 6837 34660
rect 6052 34620 6058 34632
rect 6825 34629 6837 34632
rect 6871 34629 6883 34663
rect 6825 34623 6883 34629
rect 6914 34620 6920 34672
rect 6972 34660 6978 34672
rect 6972 34632 7314 34660
rect 6972 34620 6978 34632
rect 8478 34620 8484 34672
rect 8536 34660 8542 34672
rect 11977 34663 12035 34669
rect 8536 34632 9614 34660
rect 8536 34620 8542 34632
rect 11977 34629 11989 34663
rect 12023 34660 12035 34663
rect 12066 34660 12072 34672
rect 12023 34632 12072 34660
rect 12023 34629 12035 34632
rect 11977 34623 12035 34629
rect 12066 34620 12072 34632
rect 12124 34620 12130 34672
rect 13906 34660 13912 34672
rect 13202 34632 13912 34660
rect 13906 34620 13912 34632
rect 13964 34620 13970 34672
rect 16025 34663 16083 34669
rect 16025 34629 16037 34663
rect 16071 34660 16083 34663
rect 16574 34660 16580 34672
rect 16071 34632 16580 34660
rect 16071 34629 16083 34632
rect 16025 34623 16083 34629
rect 16574 34620 16580 34632
rect 16632 34620 16638 34672
rect 17954 34620 17960 34672
rect 18012 34660 18018 34672
rect 19702 34660 19708 34672
rect 18012 34632 19708 34660
rect 18012 34620 18018 34632
rect 19702 34620 19708 34632
rect 19760 34620 19766 34672
rect 22094 34620 22100 34672
rect 22152 34620 22158 34672
rect 22462 34620 22468 34672
rect 22520 34660 22526 34672
rect 23569 34663 23627 34669
rect 23569 34660 23581 34663
rect 22520 34632 23581 34660
rect 22520 34620 22526 34632
rect 23569 34629 23581 34632
rect 23615 34629 23627 34663
rect 23569 34623 23627 34629
rect 6086 34552 6092 34604
rect 6144 34592 6150 34604
rect 6549 34595 6607 34601
rect 6549 34592 6561 34595
rect 6144 34564 6561 34592
rect 6144 34552 6150 34564
rect 6549 34561 6561 34564
rect 6595 34561 6607 34595
rect 6549 34555 6607 34561
rect 8570 34552 8576 34604
rect 8628 34592 8634 34604
rect 8849 34595 8907 34601
rect 8849 34592 8861 34595
rect 8628 34564 8861 34592
rect 8628 34552 8634 34564
rect 8849 34561 8861 34564
rect 8895 34561 8907 34595
rect 8849 34555 8907 34561
rect 8864 34524 8892 34555
rect 13354 34552 13360 34604
rect 13412 34592 13418 34604
rect 17310 34592 17316 34604
rect 13412 34564 17316 34592
rect 13412 34552 13418 34564
rect 17310 34552 17316 34564
rect 17368 34552 17374 34604
rect 21177 34595 21235 34601
rect 21177 34561 21189 34595
rect 21223 34592 21235 34595
rect 21634 34592 21640 34604
rect 21223 34564 21640 34592
rect 21223 34561 21235 34564
rect 21177 34555 21235 34561
rect 21634 34552 21640 34564
rect 21692 34552 21698 34604
rect 22112 34592 22140 34620
rect 22112 34564 22508 34592
rect 22480 34536 22508 34564
rect 23290 34552 23296 34604
rect 23348 34592 23354 34604
rect 24581 34595 24639 34601
rect 24581 34592 24593 34595
rect 23348 34564 24593 34592
rect 23348 34552 23354 34564
rect 24581 34561 24593 34564
rect 24627 34561 24639 34595
rect 24581 34555 24639 34561
rect 25314 34552 25320 34604
rect 25372 34552 25378 34604
rect 9582 34524 9588 34536
rect 8864 34496 9588 34524
rect 9582 34484 9588 34496
rect 9640 34524 9646 34536
rect 10962 34524 10968 34536
rect 9640 34496 10968 34524
rect 9640 34484 9646 34496
rect 10962 34484 10968 34496
rect 11020 34524 11026 34536
rect 11701 34527 11759 34533
rect 11701 34524 11713 34527
rect 11020 34496 11713 34524
rect 11020 34484 11026 34496
rect 11701 34493 11713 34496
rect 11747 34493 11759 34527
rect 11701 34487 11759 34493
rect 13449 34527 13507 34533
rect 13449 34493 13461 34527
rect 13495 34524 13507 34527
rect 13814 34524 13820 34536
rect 13495 34496 13820 34524
rect 13495 34493 13507 34496
rect 13449 34487 13507 34493
rect 13814 34484 13820 34496
rect 13872 34524 13878 34536
rect 14826 34524 14832 34536
rect 13872 34496 14832 34524
rect 13872 34484 13878 34496
rect 14826 34484 14832 34496
rect 14884 34484 14890 34536
rect 16117 34527 16175 34533
rect 16117 34493 16129 34527
rect 16163 34493 16175 34527
rect 16117 34487 16175 34493
rect 21269 34527 21327 34533
rect 21269 34493 21281 34527
rect 21315 34493 21327 34527
rect 21269 34487 21327 34493
rect 11146 34456 11152 34468
rect 10704 34428 11152 34456
rect 9112 34391 9170 34397
rect 9112 34357 9124 34391
rect 9158 34388 9170 34391
rect 10134 34388 10140 34400
rect 9158 34360 10140 34388
rect 9158 34357 9170 34360
rect 9112 34351 9170 34357
rect 10134 34348 10140 34360
rect 10192 34388 10198 34400
rect 10704 34388 10732 34428
rect 11146 34416 11152 34428
rect 11204 34416 11210 34468
rect 13354 34416 13360 34468
rect 13412 34456 13418 34468
rect 13412 34428 15700 34456
rect 13412 34416 13418 34428
rect 10192 34360 10732 34388
rect 10192 34348 10198 34360
rect 10778 34348 10784 34400
rect 10836 34388 10842 34400
rect 10965 34391 11023 34397
rect 10965 34388 10977 34391
rect 10836 34360 10977 34388
rect 10836 34348 10842 34360
rect 10965 34357 10977 34360
rect 11011 34388 11023 34391
rect 11790 34388 11796 34400
rect 11011 34360 11796 34388
rect 11011 34357 11023 34360
rect 10965 34351 11023 34357
rect 11790 34348 11796 34360
rect 11848 34348 11854 34400
rect 13817 34391 13875 34397
rect 13817 34357 13829 34391
rect 13863 34388 13875 34391
rect 13906 34388 13912 34400
rect 13863 34360 13912 34388
rect 13863 34357 13875 34360
rect 13817 34351 13875 34357
rect 13906 34348 13912 34360
rect 13964 34388 13970 34400
rect 15470 34388 15476 34400
rect 13964 34360 15476 34388
rect 13964 34348 13970 34360
rect 15470 34348 15476 34360
rect 15528 34348 15534 34400
rect 15562 34348 15568 34400
rect 15620 34348 15626 34400
rect 15672 34388 15700 34428
rect 15838 34416 15844 34468
rect 15896 34456 15902 34468
rect 16132 34456 16160 34487
rect 15896 34428 16160 34456
rect 15896 34416 15902 34428
rect 19518 34416 19524 34468
rect 19576 34456 19582 34468
rect 21284 34456 21312 34487
rect 22462 34484 22468 34536
rect 22520 34484 22526 34536
rect 22646 34484 22652 34536
rect 22704 34484 22710 34536
rect 23474 34484 23480 34536
rect 23532 34524 23538 34536
rect 23661 34527 23719 34533
rect 23661 34524 23673 34527
rect 23532 34496 23673 34524
rect 23532 34484 23538 34496
rect 23661 34493 23673 34496
rect 23707 34493 23719 34527
rect 23661 34487 23719 34493
rect 23842 34484 23848 34536
rect 23900 34484 23906 34536
rect 25133 34459 25191 34465
rect 25133 34456 25145 34459
rect 19576 34428 21312 34456
rect 21376 34428 25145 34456
rect 19576 34416 19582 34428
rect 20162 34388 20168 34400
rect 15672 34360 20168 34388
rect 20162 34348 20168 34360
rect 20220 34388 20226 34400
rect 21376 34388 21404 34428
rect 25133 34425 25145 34428
rect 25179 34425 25191 34459
rect 25133 34419 25191 34425
rect 20220 34360 21404 34388
rect 20220 34348 20226 34360
rect 22002 34348 22008 34400
rect 22060 34348 22066 34400
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 6914 34144 6920 34196
rect 6972 34184 6978 34196
rect 7561 34187 7619 34193
rect 7561 34184 7573 34187
rect 6972 34156 7573 34184
rect 6972 34144 6978 34156
rect 7561 34153 7573 34156
rect 7607 34153 7619 34187
rect 7561 34147 7619 34153
rect 7576 34116 7604 34147
rect 7742 34144 7748 34196
rect 7800 34144 7806 34196
rect 7834 34144 7840 34196
rect 7892 34184 7898 34196
rect 9125 34187 9183 34193
rect 9125 34184 9137 34187
rect 7892 34156 9137 34184
rect 7892 34144 7898 34156
rect 9125 34153 9137 34156
rect 9171 34153 9183 34187
rect 9125 34147 9183 34153
rect 11146 34144 11152 34196
rect 11204 34184 11210 34196
rect 12161 34187 12219 34193
rect 12161 34184 12173 34187
rect 11204 34156 12173 34184
rect 11204 34144 11210 34156
rect 12161 34153 12173 34156
rect 12207 34184 12219 34187
rect 12207 34156 13584 34184
rect 12207 34153 12219 34156
rect 12161 34147 12219 34153
rect 8478 34116 8484 34128
rect 7576 34088 8484 34116
rect 8478 34076 8484 34088
rect 8536 34076 8542 34128
rect 5534 34008 5540 34060
rect 5592 34008 5598 34060
rect 5810 34008 5816 34060
rect 5868 34048 5874 34060
rect 7285 34051 7343 34057
rect 7285 34048 7297 34051
rect 5868 34020 7297 34048
rect 5868 34008 5874 34020
rect 7285 34017 7297 34020
rect 7331 34048 7343 34051
rect 9214 34048 9220 34060
rect 7331 34020 9220 34048
rect 7331 34017 7343 34020
rect 7285 34011 7343 34017
rect 9214 34008 9220 34020
rect 9272 34048 9278 34060
rect 9677 34051 9735 34057
rect 9677 34048 9689 34051
rect 9272 34020 9689 34048
rect 9272 34008 9278 34020
rect 9677 34017 9689 34020
rect 9723 34017 9735 34051
rect 9677 34011 9735 34017
rect 10689 34051 10747 34057
rect 10689 34017 10701 34051
rect 10735 34048 10747 34051
rect 11698 34048 11704 34060
rect 10735 34020 11704 34048
rect 10735 34017 10747 34020
rect 10689 34011 10747 34017
rect 11698 34008 11704 34020
rect 11756 34008 11762 34060
rect 12618 34008 12624 34060
rect 12676 34048 12682 34060
rect 13556 34057 13584 34156
rect 13906 34144 13912 34196
rect 13964 34144 13970 34196
rect 16942 34184 16948 34196
rect 14108 34156 16948 34184
rect 13449 34051 13507 34057
rect 13449 34048 13461 34051
rect 12676 34020 13461 34048
rect 12676 34008 12682 34020
rect 13449 34017 13461 34020
rect 13495 34017 13507 34051
rect 13449 34011 13507 34017
rect 13541 34051 13599 34057
rect 13541 34017 13553 34051
rect 13587 34017 13599 34051
rect 13541 34011 13599 34017
rect 6914 33940 6920 33992
rect 6972 33940 6978 33992
rect 9582 33940 9588 33992
rect 9640 33980 9646 33992
rect 10413 33983 10471 33989
rect 10413 33980 10425 33983
rect 9640 33952 10425 33980
rect 9640 33940 9646 33952
rect 10413 33949 10425 33952
rect 10459 33949 10471 33983
rect 10413 33943 10471 33949
rect 11790 33940 11796 33992
rect 11848 33980 11854 33992
rect 12529 33983 12587 33989
rect 12529 33980 12541 33983
rect 11848 33952 12541 33980
rect 11848 33940 11854 33952
rect 12529 33949 12541 33952
rect 12575 33980 12587 33983
rect 13924 33980 13952 34144
rect 12575 33952 13952 33980
rect 12575 33949 12587 33952
rect 12529 33943 12587 33949
rect 5813 33915 5871 33921
rect 5813 33881 5825 33915
rect 5859 33881 5871 33915
rect 5813 33875 5871 33881
rect 1210 33804 1216 33856
rect 1268 33844 1274 33856
rect 1397 33847 1455 33853
rect 1397 33844 1409 33847
rect 1268 33816 1409 33844
rect 1268 33804 1274 33816
rect 1397 33813 1409 33816
rect 1443 33813 1455 33847
rect 5828 33844 5856 33875
rect 7650 33872 7656 33924
rect 7708 33912 7714 33924
rect 9493 33915 9551 33921
rect 9493 33912 9505 33915
rect 7708 33884 9505 33912
rect 7708 33872 7714 33884
rect 9493 33881 9505 33884
rect 9539 33881 9551 33915
rect 9493 33875 9551 33881
rect 7742 33844 7748 33856
rect 5828 33816 7748 33844
rect 1397 33807 1455 33813
rect 7742 33804 7748 33816
rect 7800 33844 7806 33856
rect 8386 33844 8392 33856
rect 7800 33816 8392 33844
rect 7800 33804 7806 33816
rect 8386 33804 8392 33816
rect 8444 33804 8450 33856
rect 9585 33847 9643 33853
rect 9585 33813 9597 33847
rect 9631 33844 9643 33847
rect 10962 33844 10968 33856
rect 9631 33816 10968 33844
rect 9631 33813 9643 33816
rect 9585 33807 9643 33813
rect 10962 33804 10968 33816
rect 11020 33804 11026 33856
rect 12342 33804 12348 33856
rect 12400 33844 12406 33856
rect 12526 33844 12532 33856
rect 12400 33816 12532 33844
rect 12400 33804 12406 33816
rect 12526 33804 12532 33816
rect 12584 33804 12590 33856
rect 12802 33804 12808 33856
rect 12860 33844 12866 33856
rect 12989 33847 13047 33853
rect 12989 33844 13001 33847
rect 12860 33816 13001 33844
rect 12860 33804 12866 33816
rect 12989 33813 13001 33816
rect 13035 33813 13047 33847
rect 12989 33807 13047 33813
rect 13170 33804 13176 33856
rect 13228 33844 13234 33856
rect 14108 33853 14136 34156
rect 16942 34144 16948 34156
rect 17000 34144 17006 34196
rect 17681 34187 17739 34193
rect 17681 34153 17693 34187
rect 17727 34184 17739 34187
rect 17954 34184 17960 34196
rect 17727 34156 17960 34184
rect 17727 34153 17739 34156
rect 17681 34147 17739 34153
rect 17954 34144 17960 34156
rect 18012 34144 18018 34196
rect 18046 34144 18052 34196
rect 18104 34184 18110 34196
rect 18414 34184 18420 34196
rect 18104 34156 18420 34184
rect 18104 34144 18110 34156
rect 18414 34144 18420 34156
rect 18472 34184 18478 34196
rect 18782 34184 18788 34196
rect 18472 34156 18788 34184
rect 18472 34144 18478 34156
rect 18782 34144 18788 34156
rect 18840 34144 18846 34196
rect 20533 34187 20591 34193
rect 20533 34153 20545 34187
rect 20579 34184 20591 34187
rect 20714 34184 20720 34196
rect 20579 34156 20720 34184
rect 20579 34153 20591 34156
rect 20533 34147 20591 34153
rect 20714 34144 20720 34156
rect 20772 34144 20778 34196
rect 22462 34144 22468 34196
rect 22520 34184 22526 34196
rect 23293 34187 23351 34193
rect 23293 34184 23305 34187
rect 22520 34156 23305 34184
rect 22520 34144 22526 34156
rect 23293 34153 23305 34156
rect 23339 34153 23351 34187
rect 23293 34147 23351 34153
rect 25314 34144 25320 34196
rect 25372 34144 25378 34196
rect 17862 34076 17868 34128
rect 17920 34116 17926 34128
rect 19429 34119 19487 34125
rect 19429 34116 19441 34119
rect 17920 34088 19441 34116
rect 17920 34076 17926 34088
rect 19429 34085 19441 34088
rect 19475 34085 19487 34119
rect 19429 34079 19487 34085
rect 22281 34119 22339 34125
rect 22281 34085 22293 34119
rect 22327 34116 22339 34119
rect 23842 34116 23848 34128
rect 22327 34088 23848 34116
rect 22327 34085 22339 34088
rect 22281 34079 22339 34085
rect 23842 34076 23848 34088
rect 23900 34076 23906 34128
rect 15930 34008 15936 34060
rect 15988 34008 15994 34060
rect 18414 34008 18420 34060
rect 18472 34048 18478 34060
rect 19061 34051 19119 34057
rect 19061 34048 19073 34051
rect 18472 34020 19073 34048
rect 18472 34008 18478 34020
rect 19061 34017 19073 34020
rect 19107 34048 19119 34051
rect 19981 34051 20039 34057
rect 19981 34048 19993 34051
rect 19107 34020 19993 34048
rect 19107 34017 19119 34020
rect 19061 34011 19119 34017
rect 19981 34017 19993 34020
rect 20027 34017 20039 34051
rect 19981 34011 20039 34017
rect 21358 34008 21364 34060
rect 21416 34048 21422 34060
rect 21637 34051 21695 34057
rect 21637 34048 21649 34051
rect 21416 34020 21649 34048
rect 21416 34008 21422 34020
rect 21637 34017 21649 34020
rect 21683 34017 21695 34051
rect 21637 34011 21695 34017
rect 21910 34008 21916 34060
rect 21968 34048 21974 34060
rect 22741 34051 22799 34057
rect 22741 34048 22753 34051
rect 21968 34020 22753 34048
rect 21968 34008 21974 34020
rect 22741 34017 22753 34020
rect 22787 34017 22799 34051
rect 22741 34011 22799 34017
rect 22925 34051 22983 34057
rect 22925 34017 22937 34051
rect 22971 34048 22983 34051
rect 23382 34048 23388 34060
rect 22971 34020 23388 34048
rect 22971 34017 22983 34020
rect 22925 34011 22983 34017
rect 23382 34008 23388 34020
rect 23440 34008 23446 34060
rect 19797 33983 19855 33989
rect 19797 33949 19809 33983
rect 19843 33980 19855 33983
rect 20070 33980 20076 33992
rect 19843 33952 20076 33980
rect 19843 33949 19855 33952
rect 19797 33943 19855 33949
rect 20070 33940 20076 33952
rect 20128 33940 20134 33992
rect 21450 33940 21456 33992
rect 21508 33980 21514 33992
rect 21545 33983 21603 33989
rect 21545 33980 21557 33983
rect 21508 33952 21557 33980
rect 21508 33940 21514 33952
rect 21545 33949 21557 33952
rect 21591 33980 21603 33983
rect 21591 33952 22094 33980
rect 21591 33949 21603 33952
rect 21545 33943 21603 33949
rect 16206 33872 16212 33924
rect 16264 33872 16270 33924
rect 17586 33912 17592 33924
rect 17434 33884 17592 33912
rect 17586 33872 17592 33884
rect 17644 33912 17650 33924
rect 18046 33912 18052 33924
rect 17644 33884 18052 33912
rect 17644 33872 17650 33884
rect 18046 33872 18052 33884
rect 18104 33872 18110 33924
rect 19889 33915 19947 33921
rect 19889 33881 19901 33915
rect 19935 33912 19947 33915
rect 20254 33912 20260 33924
rect 19935 33884 20260 33912
rect 19935 33881 19947 33884
rect 19889 33875 19947 33881
rect 20254 33872 20260 33884
rect 20312 33872 20318 33924
rect 22066 33912 22094 33952
rect 24762 33940 24768 33992
rect 24820 33940 24826 33992
rect 23382 33912 23388 33924
rect 22066 33884 23388 33912
rect 23382 33872 23388 33884
rect 23440 33872 23446 33924
rect 24026 33872 24032 33924
rect 24084 33912 24090 33924
rect 24302 33912 24308 33924
rect 24084 33884 24308 33912
rect 24084 33872 24090 33884
rect 24302 33872 24308 33884
rect 24360 33912 24366 33924
rect 25409 33915 25467 33921
rect 25409 33912 25421 33915
rect 24360 33884 25421 33912
rect 24360 33872 24366 33884
rect 25409 33881 25421 33884
rect 25455 33881 25467 33915
rect 25409 33875 25467 33881
rect 13357 33847 13415 33853
rect 13357 33844 13369 33847
rect 13228 33816 13369 33844
rect 13228 33804 13234 33816
rect 13357 33813 13369 33816
rect 13403 33844 13415 33847
rect 14093 33847 14151 33853
rect 14093 33844 14105 33847
rect 13403 33816 14105 33844
rect 13403 33813 13415 33816
rect 13357 33807 13415 33813
rect 14093 33813 14105 33816
rect 14139 33813 14151 33847
rect 14093 33807 14151 33813
rect 16298 33804 16304 33856
rect 16356 33844 16362 33856
rect 19150 33844 19156 33856
rect 16356 33816 19156 33844
rect 16356 33804 16362 33816
rect 19150 33804 19156 33816
rect 19208 33804 19214 33856
rect 20622 33804 20628 33856
rect 20680 33804 20686 33856
rect 20714 33804 20720 33856
rect 20772 33844 20778 33856
rect 21085 33847 21143 33853
rect 21085 33844 21097 33847
rect 20772 33816 21097 33844
rect 20772 33804 20778 33816
rect 21085 33813 21097 33816
rect 21131 33813 21143 33847
rect 21085 33807 21143 33813
rect 21450 33804 21456 33856
rect 21508 33804 21514 33856
rect 22462 33804 22468 33856
rect 22520 33844 22526 33856
rect 22649 33847 22707 33853
rect 22649 33844 22661 33847
rect 22520 33816 22661 33844
rect 22520 33804 22526 33816
rect 22649 33813 22661 33816
rect 22695 33813 22707 33847
rect 22649 33807 22707 33813
rect 24578 33804 24584 33856
rect 24636 33804 24642 33856
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 6914 33600 6920 33652
rect 6972 33640 6978 33652
rect 7101 33643 7159 33649
rect 7101 33640 7113 33643
rect 6972 33612 7113 33640
rect 6972 33600 6978 33612
rect 7101 33609 7113 33612
rect 7147 33609 7159 33643
rect 7101 33603 7159 33609
rect 10410 33600 10416 33652
rect 10468 33600 10474 33652
rect 10870 33600 10876 33652
rect 10928 33600 10934 33652
rect 11330 33600 11336 33652
rect 11388 33640 11394 33652
rect 12897 33643 12955 33649
rect 12897 33640 12909 33643
rect 11388 33612 12909 33640
rect 11388 33600 11394 33612
rect 12897 33609 12909 33612
rect 12943 33609 12955 33643
rect 12897 33603 12955 33609
rect 13354 33600 13360 33652
rect 13412 33600 13418 33652
rect 14550 33640 14556 33652
rect 14108 33612 14556 33640
rect 10962 33532 10968 33584
rect 11020 33572 11026 33584
rect 12618 33572 12624 33584
rect 11020 33544 12624 33572
rect 11020 33532 11026 33544
rect 12618 33532 12624 33544
rect 12676 33532 12682 33584
rect 12805 33575 12863 33581
rect 12805 33541 12817 33575
rect 12851 33572 12863 33575
rect 13372 33572 13400 33600
rect 12851 33544 13400 33572
rect 12851 33541 12863 33544
rect 12805 33535 12863 33541
rect 1210 33464 1216 33516
rect 1268 33504 1274 33516
rect 1581 33507 1639 33513
rect 1581 33504 1593 33507
rect 1268 33476 1593 33504
rect 1268 33464 1274 33476
rect 1581 33473 1593 33476
rect 1627 33473 1639 33507
rect 1581 33467 1639 33473
rect 10781 33507 10839 33513
rect 10781 33473 10793 33507
rect 10827 33504 10839 33507
rect 11882 33504 11888 33516
rect 10827 33476 11888 33504
rect 10827 33473 10839 33476
rect 10781 33467 10839 33473
rect 11882 33464 11888 33476
rect 11940 33464 11946 33516
rect 12526 33464 12532 33516
rect 12584 33504 12590 33516
rect 14108 33513 14136 33612
rect 14550 33600 14556 33612
rect 14608 33640 14614 33652
rect 15930 33640 15936 33652
rect 14608 33612 15936 33640
rect 14608 33600 14614 33612
rect 15930 33600 15936 33612
rect 15988 33600 15994 33652
rect 16209 33643 16267 33649
rect 16209 33609 16221 33643
rect 16255 33640 16267 33643
rect 17586 33640 17592 33652
rect 16255 33612 17592 33640
rect 16255 33609 16267 33612
rect 16209 33603 16267 33609
rect 13265 33507 13323 33513
rect 13265 33504 13277 33507
rect 12584 33476 13277 33504
rect 12584 33464 12590 33476
rect 13265 33473 13277 33476
rect 13311 33473 13323 33507
rect 13265 33467 13323 33473
rect 14093 33507 14151 33513
rect 14093 33473 14105 33507
rect 14139 33473 14151 33507
rect 14093 33467 14151 33473
rect 15470 33464 15476 33516
rect 15528 33464 15534 33516
rect 15930 33464 15936 33516
rect 15988 33504 15994 33516
rect 16224 33504 16252 33603
rect 17586 33600 17592 33612
rect 17644 33600 17650 33652
rect 19797 33643 19855 33649
rect 19797 33609 19809 33643
rect 19843 33640 19855 33643
rect 19886 33640 19892 33652
rect 19843 33612 19892 33640
rect 19843 33609 19855 33612
rect 19797 33603 19855 33609
rect 19886 33600 19892 33612
rect 19944 33600 19950 33652
rect 21358 33640 21364 33652
rect 20088 33612 21364 33640
rect 18322 33572 18328 33584
rect 18064 33544 18328 33572
rect 18064 33513 18092 33544
rect 18322 33532 18328 33544
rect 18380 33532 18386 33584
rect 18782 33532 18788 33584
rect 18840 33532 18846 33584
rect 15988 33476 16252 33504
rect 18049 33507 18107 33513
rect 15988 33464 15994 33476
rect 18049 33473 18061 33507
rect 18095 33473 18107 33507
rect 18049 33467 18107 33473
rect 5350 33396 5356 33448
rect 5408 33396 5414 33448
rect 9766 33396 9772 33448
rect 9824 33396 9830 33448
rect 10965 33439 11023 33445
rect 10965 33405 10977 33439
rect 11011 33405 11023 33439
rect 10965 33399 11023 33405
rect 8294 33328 8300 33380
rect 8352 33368 8358 33380
rect 10980 33368 11008 33399
rect 13446 33396 13452 33448
rect 13504 33396 13510 33448
rect 14369 33439 14427 33445
rect 14369 33405 14381 33439
rect 14415 33436 14427 33439
rect 16298 33436 16304 33448
rect 14415 33408 16304 33436
rect 14415 33405 14427 33408
rect 14369 33399 14427 33405
rect 16298 33396 16304 33408
rect 16356 33396 16362 33448
rect 18325 33439 18383 33445
rect 18325 33405 18337 33439
rect 18371 33436 18383 33439
rect 20088 33436 20116 33612
rect 21358 33600 21364 33612
rect 21416 33600 21422 33652
rect 21450 33600 21456 33652
rect 21508 33640 21514 33652
rect 22649 33643 22707 33649
rect 22649 33640 22661 33643
rect 21508 33612 22661 33640
rect 21508 33600 21514 33612
rect 22649 33609 22661 33612
rect 22695 33609 22707 33643
rect 22649 33603 22707 33609
rect 25038 33600 25044 33652
rect 25096 33640 25102 33652
rect 25225 33643 25283 33649
rect 25225 33640 25237 33643
rect 25096 33612 25237 33640
rect 25096 33600 25102 33612
rect 25225 33609 25237 33612
rect 25271 33609 25283 33643
rect 25225 33603 25283 33609
rect 20254 33532 20260 33584
rect 20312 33572 20318 33584
rect 20312 33544 20760 33572
rect 20312 33532 20318 33544
rect 20622 33464 20628 33516
rect 20680 33464 20686 33516
rect 20732 33513 20760 33544
rect 24026 33532 24032 33584
rect 24084 33572 24090 33584
rect 24084 33544 24242 33572
rect 24084 33532 24090 33544
rect 20717 33507 20775 33513
rect 20717 33473 20729 33507
rect 20763 33473 20775 33507
rect 20717 33467 20775 33473
rect 21450 33464 21456 33516
rect 21508 33504 21514 33516
rect 22094 33504 22100 33516
rect 21508 33476 22100 33504
rect 21508 33464 21514 33476
rect 22094 33464 22100 33476
rect 22152 33464 22158 33516
rect 22186 33464 22192 33516
rect 22244 33504 22250 33516
rect 23477 33507 23535 33513
rect 23477 33504 23489 33507
rect 22244 33476 23489 33504
rect 22244 33464 22250 33476
rect 23477 33473 23489 33476
rect 23523 33473 23535 33507
rect 23477 33467 23535 33473
rect 18371 33408 20116 33436
rect 18371 33405 18383 33408
rect 18325 33399 18383 33405
rect 20438 33396 20444 33448
rect 20496 33436 20502 33448
rect 20809 33439 20867 33445
rect 20809 33436 20821 33439
rect 20496 33408 20821 33436
rect 20496 33396 20502 33408
rect 20809 33405 20821 33408
rect 20855 33405 20867 33439
rect 20809 33399 20867 33405
rect 21174 33396 21180 33448
rect 21232 33436 21238 33448
rect 22005 33439 22063 33445
rect 22005 33436 22017 33439
rect 21232 33408 22017 33436
rect 21232 33396 21238 33408
rect 22005 33405 22017 33408
rect 22051 33405 22063 33439
rect 22005 33399 22063 33405
rect 23750 33396 23756 33448
rect 23808 33396 23814 33448
rect 8352 33340 11008 33368
rect 8352 33328 8358 33340
rect 15470 33328 15476 33380
rect 15528 33368 15534 33380
rect 15930 33368 15936 33380
rect 15528 33340 15936 33368
rect 15528 33328 15534 33340
rect 15930 33328 15936 33340
rect 15988 33328 15994 33380
rect 20257 33371 20315 33377
rect 20257 33337 20269 33371
rect 20303 33368 20315 33371
rect 23474 33368 23480 33380
rect 20303 33340 20760 33368
rect 20303 33337 20315 33340
rect 20257 33331 20315 33337
rect 1762 33260 1768 33312
rect 1820 33300 1826 33312
rect 2225 33303 2283 33309
rect 2225 33300 2237 33303
rect 1820 33272 2237 33300
rect 1820 33260 1826 33272
rect 2225 33269 2237 33272
rect 2271 33269 2283 33303
rect 2225 33263 2283 33269
rect 7098 33260 7104 33312
rect 7156 33300 7162 33312
rect 10594 33300 10600 33312
rect 7156 33272 10600 33300
rect 7156 33260 7162 33272
rect 10594 33260 10600 33272
rect 10652 33260 10658 33312
rect 12526 33260 12532 33312
rect 12584 33260 12590 33312
rect 13170 33260 13176 33312
rect 13228 33300 13234 33312
rect 13446 33300 13452 33312
rect 13228 33272 13452 33300
rect 13228 33260 13234 33272
rect 13446 33260 13452 33272
rect 13504 33260 13510 33312
rect 13538 33260 13544 33312
rect 13596 33300 13602 33312
rect 15838 33300 15844 33312
rect 13596 33272 15844 33300
rect 13596 33260 13602 33272
rect 15838 33260 15844 33272
rect 15896 33260 15902 33312
rect 20732 33300 20760 33340
rect 20916 33340 23480 33368
rect 20916 33300 20944 33340
rect 23474 33328 23480 33340
rect 23532 33328 23538 33380
rect 20732 33272 20944 33300
rect 21358 33260 21364 33312
rect 21416 33300 21422 33312
rect 22278 33300 22284 33312
rect 21416 33272 22284 33300
rect 21416 33260 21422 33272
rect 22278 33260 22284 33272
rect 22336 33260 22342 33312
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 7466 33056 7472 33108
rect 7524 33056 7530 33108
rect 9306 33056 9312 33108
rect 9364 33096 9370 33108
rect 9401 33099 9459 33105
rect 9401 33096 9413 33099
rect 9364 33068 9413 33096
rect 9364 33056 9370 33068
rect 9401 33065 9413 33068
rect 9447 33065 9459 33099
rect 9401 33059 9459 33065
rect 10594 33056 10600 33108
rect 10652 33056 10658 33108
rect 11054 33056 11060 33108
rect 11112 33096 11118 33108
rect 11149 33099 11207 33105
rect 11149 33096 11161 33099
rect 11112 33068 11161 33096
rect 11112 33056 11118 33068
rect 11149 33065 11161 33068
rect 11195 33065 11207 33099
rect 11149 33059 11207 33065
rect 12250 33056 12256 33108
rect 12308 33056 12314 33108
rect 12434 33056 12440 33108
rect 12492 33096 12498 33108
rect 13906 33096 13912 33108
rect 12492 33068 13912 33096
rect 12492 33056 12498 33068
rect 13906 33056 13912 33068
rect 13964 33056 13970 33108
rect 13998 33056 14004 33108
rect 14056 33096 14062 33108
rect 19429 33099 19487 33105
rect 19429 33096 19441 33099
rect 14056 33068 19441 33096
rect 14056 33056 14062 33068
rect 19429 33065 19441 33068
rect 19475 33065 19487 33099
rect 19429 33059 19487 33065
rect 19797 33099 19855 33105
rect 19797 33065 19809 33099
rect 19843 33096 19855 33099
rect 22462 33096 22468 33108
rect 19843 33068 22468 33096
rect 19843 33065 19855 33068
rect 19797 33059 19855 33065
rect 7009 33031 7067 33037
rect 7009 32997 7021 33031
rect 7055 33028 7067 33031
rect 7558 33028 7564 33040
rect 7055 33000 7564 33028
rect 7055 32997 7067 33000
rect 7009 32991 7067 32997
rect 7558 32988 7564 33000
rect 7616 32988 7622 33040
rect 5261 32963 5319 32969
rect 5261 32929 5273 32963
rect 5307 32960 5319 32963
rect 5534 32960 5540 32972
rect 5307 32932 5540 32960
rect 5307 32929 5319 32932
rect 5261 32923 5319 32929
rect 5534 32920 5540 32932
rect 5592 32920 5598 32972
rect 8113 32963 8171 32969
rect 8113 32929 8125 32963
rect 8159 32960 8171 32963
rect 8294 32960 8300 32972
rect 8159 32932 8300 32960
rect 8159 32929 8171 32932
rect 8113 32923 8171 32929
rect 1762 32852 1768 32904
rect 1820 32852 1826 32904
rect 6914 32892 6920 32904
rect 6670 32864 6920 32892
rect 6914 32852 6920 32864
rect 6972 32852 6978 32904
rect 8128 32892 8156 32923
rect 8294 32920 8300 32932
rect 8352 32920 8358 32972
rect 10045 32963 10103 32969
rect 10045 32929 10057 32963
rect 10091 32960 10103 32963
rect 10134 32960 10140 32972
rect 10091 32932 10140 32960
rect 10091 32929 10103 32932
rect 10045 32923 10103 32929
rect 10134 32920 10140 32932
rect 10192 32920 10198 32972
rect 10873 32963 10931 32969
rect 10873 32929 10885 32963
rect 10919 32960 10931 32963
rect 11606 32960 11612 32972
rect 10919 32932 11612 32960
rect 10919 32929 10931 32932
rect 10873 32923 10931 32929
rect 11606 32920 11612 32932
rect 11664 32920 11670 32972
rect 11793 32963 11851 32969
rect 11793 32929 11805 32963
rect 11839 32960 11851 32963
rect 12268 32960 12296 33056
rect 14918 32988 14924 33040
rect 14976 33028 14982 33040
rect 14976 33000 19380 33028
rect 14976 32988 14982 33000
rect 11839 32932 12296 32960
rect 11839 32929 11851 32932
rect 11793 32923 11851 32929
rect 14274 32920 14280 32972
rect 14332 32960 14338 32972
rect 14737 32963 14795 32969
rect 14737 32960 14749 32963
rect 14332 32932 14749 32960
rect 14332 32920 14338 32932
rect 14737 32929 14749 32932
rect 14783 32929 14795 32963
rect 14737 32923 14795 32929
rect 14826 32920 14832 32972
rect 14884 32920 14890 32972
rect 16482 32920 16488 32972
rect 16540 32960 16546 32972
rect 16669 32963 16727 32969
rect 16669 32960 16681 32963
rect 16540 32932 16681 32960
rect 16540 32920 16546 32932
rect 16669 32929 16681 32932
rect 16715 32960 16727 32963
rect 18506 32960 18512 32972
rect 16715 32932 18512 32960
rect 16715 32929 16727 32932
rect 16669 32923 16727 32929
rect 18506 32920 18512 32932
rect 18564 32920 18570 32972
rect 7668 32864 8156 32892
rect 5537 32827 5595 32833
rect 5537 32793 5549 32827
rect 5583 32793 5595 32827
rect 5537 32787 5595 32793
rect 1578 32716 1584 32768
rect 1636 32716 1642 32768
rect 5552 32756 5580 32787
rect 7668 32756 7696 32864
rect 9766 32852 9772 32904
rect 9824 32852 9830 32904
rect 10594 32852 10600 32904
rect 10652 32892 10658 32904
rect 11517 32895 11575 32901
rect 11517 32892 11529 32895
rect 10652 32864 11529 32892
rect 10652 32852 10658 32864
rect 11517 32861 11529 32864
rect 11563 32892 11575 32895
rect 11974 32892 11980 32904
rect 11563 32864 11980 32892
rect 11563 32861 11575 32864
rect 11517 32855 11575 32861
rect 11974 32852 11980 32864
rect 12032 32852 12038 32904
rect 12526 32852 12532 32904
rect 12584 32892 12590 32904
rect 13630 32892 13636 32904
rect 12584 32864 13636 32892
rect 12584 32852 12590 32864
rect 13630 32852 13636 32864
rect 13688 32892 13694 32904
rect 15749 32895 15807 32901
rect 15749 32892 15761 32895
rect 13688 32864 15761 32892
rect 13688 32852 13694 32864
rect 15749 32861 15761 32864
rect 15795 32892 15807 32895
rect 16577 32895 16635 32901
rect 15795 32864 15976 32892
rect 15795 32861 15807 32864
rect 15749 32855 15807 32861
rect 7742 32784 7748 32836
rect 7800 32824 7806 32836
rect 7929 32827 7987 32833
rect 7929 32824 7941 32827
rect 7800 32796 7941 32824
rect 7800 32784 7806 32796
rect 7929 32793 7941 32796
rect 7975 32793 7987 32827
rect 15838 32824 15844 32836
rect 7929 32787 7987 32793
rect 14292 32796 15844 32824
rect 5552 32728 7696 32756
rect 7834 32716 7840 32768
rect 7892 32716 7898 32768
rect 9490 32716 9496 32768
rect 9548 32756 9554 32768
rect 9861 32759 9919 32765
rect 9861 32756 9873 32759
rect 9548 32728 9873 32756
rect 9548 32716 9554 32728
rect 9861 32725 9873 32728
rect 9907 32725 9919 32759
rect 9861 32719 9919 32725
rect 11606 32716 11612 32768
rect 11664 32756 11670 32768
rect 13998 32756 14004 32768
rect 11664 32728 14004 32756
rect 11664 32716 11670 32728
rect 13998 32716 14004 32728
rect 14056 32716 14062 32768
rect 14292 32765 14320 32796
rect 15838 32784 15844 32796
rect 15896 32784 15902 32836
rect 15948 32824 15976 32864
rect 16577 32861 16589 32895
rect 16623 32892 16635 32895
rect 16758 32892 16764 32904
rect 16623 32864 16764 32892
rect 16623 32861 16635 32864
rect 16577 32855 16635 32861
rect 16758 32852 16764 32864
rect 16816 32892 16822 32904
rect 17313 32895 17371 32901
rect 17313 32892 17325 32895
rect 16816 32864 17325 32892
rect 16816 32852 16822 32864
rect 17313 32861 17325 32864
rect 17359 32861 17371 32895
rect 17313 32855 17371 32861
rect 17221 32827 17279 32833
rect 15948 32796 16252 32824
rect 14277 32759 14335 32765
rect 14277 32725 14289 32759
rect 14323 32725 14335 32759
rect 14277 32719 14335 32725
rect 14642 32716 14648 32768
rect 14700 32716 14706 32768
rect 16114 32716 16120 32768
rect 16172 32716 16178 32768
rect 16224 32756 16252 32796
rect 17221 32793 17233 32827
rect 17267 32824 17279 32827
rect 17586 32824 17592 32836
rect 17267 32796 17592 32824
rect 17267 32793 17279 32796
rect 17221 32787 17279 32793
rect 17586 32784 17592 32796
rect 17644 32784 17650 32836
rect 19352 32824 19380 33000
rect 19444 32960 19472 33059
rect 22462 33056 22468 33068
rect 22520 33056 22526 33108
rect 23566 33056 23572 33108
rect 23624 33096 23630 33108
rect 25133 33099 25191 33105
rect 25133 33096 25145 33099
rect 23624 33068 25145 33096
rect 23624 33056 23630 33068
rect 25133 33065 25145 33068
rect 25179 33065 25191 33099
rect 25133 33059 25191 33065
rect 20993 33031 21051 33037
rect 20993 32997 21005 33031
rect 21039 33028 21051 33031
rect 22094 33028 22100 33040
rect 21039 33000 22100 33028
rect 21039 32997 21051 33000
rect 20993 32991 21051 32997
rect 22094 32988 22100 33000
rect 22152 32988 22158 33040
rect 22278 33028 22284 33040
rect 22204 33000 22284 33028
rect 20257 32963 20315 32969
rect 20257 32960 20269 32963
rect 19444 32932 20269 32960
rect 20257 32929 20269 32932
rect 20303 32929 20315 32963
rect 20257 32923 20315 32929
rect 20441 32963 20499 32969
rect 20441 32929 20453 32963
rect 20487 32960 20499 32963
rect 21266 32960 21272 32972
rect 20487 32932 21272 32960
rect 20487 32929 20499 32932
rect 20441 32923 20499 32929
rect 21266 32920 21272 32932
rect 21324 32920 21330 32972
rect 21542 32920 21548 32972
rect 21600 32920 21606 32972
rect 22204 32960 22232 33000
rect 22278 32988 22284 33000
rect 22336 33028 22342 33040
rect 22925 33031 22983 33037
rect 22925 33028 22937 33031
rect 22336 33000 22937 33028
rect 22336 32988 22342 33000
rect 22925 32997 22937 33000
rect 22971 33028 22983 33031
rect 23658 33028 23664 33040
rect 22971 33000 23664 33028
rect 22971 32997 22983 33000
rect 22925 32991 22983 32997
rect 23658 32988 23664 33000
rect 23716 32988 23722 33040
rect 24026 32960 24032 32972
rect 21836 32932 22232 32960
rect 22296 32932 24032 32960
rect 20165 32895 20223 32901
rect 20165 32861 20177 32895
rect 20211 32892 20223 32895
rect 21174 32892 21180 32904
rect 20211 32864 21180 32892
rect 20211 32861 20223 32864
rect 20165 32855 20223 32861
rect 21174 32852 21180 32864
rect 21232 32852 21238 32904
rect 21836 32892 21864 32932
rect 22296 32892 22324 32932
rect 24026 32920 24032 32932
rect 24084 32920 24090 32972
rect 21468 32888 21864 32892
rect 21376 32864 21864 32888
rect 22204 32864 22324 32892
rect 21376 32860 21496 32864
rect 20622 32824 20628 32836
rect 19352 32796 20628 32824
rect 20622 32784 20628 32796
rect 20680 32784 20686 32836
rect 16485 32759 16543 32765
rect 16485 32756 16497 32759
rect 16224 32728 16497 32756
rect 16485 32725 16497 32728
rect 16531 32725 16543 32759
rect 16485 32719 16543 32725
rect 17957 32759 18015 32765
rect 17957 32725 17969 32759
rect 18003 32756 18015 32759
rect 18598 32756 18604 32768
rect 18003 32728 18604 32756
rect 18003 32725 18015 32728
rect 17957 32719 18015 32725
rect 18598 32716 18604 32728
rect 18656 32716 18662 32768
rect 21376 32765 21404 32860
rect 21361 32759 21419 32765
rect 21361 32725 21373 32759
rect 21407 32725 21419 32759
rect 21361 32719 21419 32725
rect 21453 32759 21511 32765
rect 21453 32725 21465 32759
rect 21499 32756 21511 32759
rect 21910 32756 21916 32768
rect 21499 32728 21916 32756
rect 21499 32725 21511 32728
rect 21453 32719 21511 32725
rect 21910 32716 21916 32728
rect 21968 32716 21974 32768
rect 22204 32765 22232 32864
rect 22370 32852 22376 32904
rect 22428 32852 22434 32904
rect 24857 32895 24915 32901
rect 24857 32861 24869 32895
rect 24903 32892 24915 32895
rect 25314 32892 25320 32904
rect 24903 32864 25320 32892
rect 24903 32861 24915 32864
rect 24857 32855 24915 32861
rect 25314 32852 25320 32864
rect 25372 32852 25378 32904
rect 22373 32851 22431 32852
rect 22189 32759 22247 32765
rect 22189 32725 22201 32759
rect 22235 32725 22247 32759
rect 22189 32719 22247 32725
rect 22738 32716 22744 32768
rect 22796 32716 22802 32768
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 4614 32512 4620 32564
rect 4672 32512 4678 32564
rect 4982 32512 4988 32564
rect 5040 32512 5046 32564
rect 5350 32512 5356 32564
rect 5408 32512 5414 32564
rect 6917 32555 6975 32561
rect 6917 32521 6929 32555
rect 6963 32552 6975 32555
rect 7834 32552 7840 32564
rect 6963 32524 7840 32552
rect 6963 32521 6975 32524
rect 6917 32515 6975 32521
rect 7834 32512 7840 32524
rect 7892 32512 7898 32564
rect 11977 32555 12035 32561
rect 11977 32521 11989 32555
rect 12023 32552 12035 32555
rect 14642 32552 14648 32564
rect 12023 32524 14648 32552
rect 12023 32521 12035 32524
rect 11977 32515 12035 32521
rect 14642 32512 14648 32524
rect 14700 32512 14706 32564
rect 14734 32512 14740 32564
rect 14792 32552 14798 32564
rect 18417 32555 18475 32561
rect 18417 32552 18429 32555
rect 14792 32524 18429 32552
rect 14792 32512 14798 32524
rect 18417 32521 18429 32524
rect 18463 32521 18475 32555
rect 18417 32515 18475 32521
rect 4632 32484 4660 32512
rect 5442 32484 5448 32496
rect 4632 32456 5448 32484
rect 5442 32444 5448 32456
rect 5500 32444 5506 32496
rect 5534 32444 5540 32496
rect 5592 32444 5598 32496
rect 9122 32484 9128 32496
rect 9062 32456 9128 32484
rect 9122 32444 9128 32456
rect 9180 32484 9186 32496
rect 9180 32456 9674 32484
rect 9180 32444 9186 32456
rect 5552 32416 5580 32444
rect 6178 32416 6184 32428
rect 5552 32388 6184 32416
rect 6178 32376 6184 32388
rect 6236 32416 6242 32428
rect 7561 32419 7619 32425
rect 7561 32416 7573 32419
rect 6236 32388 7573 32416
rect 6236 32376 6242 32388
rect 7561 32385 7573 32388
rect 7607 32385 7619 32419
rect 7561 32379 7619 32385
rect 5258 32308 5264 32360
rect 5316 32348 5322 32360
rect 5537 32351 5595 32357
rect 5537 32348 5549 32351
rect 5316 32320 5549 32348
rect 5316 32308 5322 32320
rect 5537 32317 5549 32320
rect 5583 32317 5595 32351
rect 7837 32351 7895 32357
rect 7837 32348 7849 32351
rect 5537 32311 5595 32317
rect 7576 32320 7849 32348
rect 7576 32292 7604 32320
rect 7837 32317 7849 32320
rect 7883 32317 7895 32351
rect 7837 32311 7895 32317
rect 8386 32308 8392 32360
rect 8444 32348 8450 32360
rect 9398 32348 9404 32360
rect 8444 32320 9404 32348
rect 8444 32308 8450 32320
rect 9398 32308 9404 32320
rect 9456 32308 9462 32360
rect 7558 32240 7564 32292
rect 7616 32240 7622 32292
rect 9306 32172 9312 32224
rect 9364 32172 9370 32224
rect 9646 32212 9674 32456
rect 13722 32444 13728 32496
rect 13780 32484 13786 32496
rect 15102 32484 15108 32496
rect 13780 32456 15108 32484
rect 13780 32444 13786 32456
rect 15102 32444 15108 32456
rect 15160 32444 15166 32496
rect 17218 32444 17224 32496
rect 17276 32444 17282 32496
rect 12345 32419 12403 32425
rect 12345 32385 12357 32419
rect 12391 32416 12403 32419
rect 13173 32419 13231 32425
rect 13173 32416 13185 32419
rect 12391 32388 13185 32416
rect 12391 32385 12403 32388
rect 12345 32379 12403 32385
rect 13173 32385 13185 32388
rect 13219 32385 13231 32419
rect 13173 32379 13231 32385
rect 14550 32376 14556 32428
rect 14608 32376 14614 32428
rect 15930 32376 15936 32428
rect 15988 32376 15994 32428
rect 18432 32416 18460 32515
rect 18506 32512 18512 32564
rect 18564 32552 18570 32564
rect 19061 32555 19119 32561
rect 19061 32552 19073 32555
rect 18564 32524 19073 32552
rect 18564 32512 18570 32524
rect 19061 32521 19073 32524
rect 19107 32521 19119 32555
rect 19061 32515 19119 32521
rect 21082 32512 21088 32564
rect 21140 32512 21146 32564
rect 21174 32512 21180 32564
rect 21232 32552 21238 32564
rect 21910 32552 21916 32564
rect 21232 32524 21916 32552
rect 21232 32512 21238 32524
rect 21910 32512 21916 32524
rect 21968 32512 21974 32564
rect 22370 32512 22376 32564
rect 22428 32552 22434 32564
rect 22738 32552 22744 32564
rect 22428 32524 22744 32552
rect 22428 32512 22434 32524
rect 22738 32512 22744 32524
rect 22796 32512 22802 32564
rect 21100 32484 21128 32512
rect 21100 32456 22048 32484
rect 20162 32416 20168 32428
rect 18432 32388 20168 32416
rect 9858 32308 9864 32360
rect 9916 32308 9922 32360
rect 11701 32351 11759 32357
rect 11701 32317 11713 32351
rect 11747 32348 11759 32351
rect 12250 32348 12256 32360
rect 11747 32320 12256 32348
rect 11747 32317 11759 32320
rect 11701 32311 11759 32317
rect 12250 32308 12256 32320
rect 12308 32348 12314 32360
rect 12437 32351 12495 32357
rect 12437 32348 12449 32351
rect 12308 32320 12449 32348
rect 12308 32308 12314 32320
rect 12437 32317 12449 32320
rect 12483 32317 12495 32351
rect 12437 32311 12495 32317
rect 12529 32351 12587 32357
rect 12529 32317 12541 32351
rect 12575 32317 12587 32351
rect 12529 32311 12587 32317
rect 12066 32240 12072 32292
rect 12124 32280 12130 32292
rect 12544 32280 12572 32311
rect 14826 32308 14832 32360
rect 14884 32308 14890 32360
rect 16298 32308 16304 32360
rect 16356 32308 16362 32360
rect 17313 32351 17371 32357
rect 17313 32317 17325 32351
rect 17359 32317 17371 32351
rect 17313 32311 17371 32317
rect 12124 32252 12572 32280
rect 12124 32240 12130 32252
rect 16114 32240 16120 32292
rect 16172 32280 16178 32292
rect 17328 32280 17356 32311
rect 17494 32308 17500 32360
rect 17552 32308 17558 32360
rect 18598 32308 18604 32360
rect 18656 32308 18662 32360
rect 19260 32357 19288 32388
rect 20162 32376 20168 32388
rect 20220 32376 20226 32428
rect 20257 32419 20315 32425
rect 20257 32385 20269 32419
rect 20303 32385 20315 32419
rect 20257 32379 20315 32385
rect 19245 32351 19303 32357
rect 19245 32317 19257 32351
rect 19291 32348 19303 32351
rect 20272 32348 20300 32379
rect 21082 32376 21088 32428
rect 21140 32416 21146 32428
rect 21450 32416 21456 32428
rect 21140 32388 21456 32416
rect 21140 32376 21146 32388
rect 21450 32376 21456 32388
rect 21508 32416 21514 32428
rect 22020 32416 22048 32456
rect 22094 32444 22100 32496
rect 22152 32484 22158 32496
rect 22278 32484 22284 32496
rect 22152 32456 22284 32484
rect 22152 32444 22158 32456
rect 22278 32444 22284 32456
rect 22336 32444 22342 32496
rect 22373 32419 22431 32425
rect 22373 32416 22385 32419
rect 21508 32388 21956 32416
rect 22020 32388 22385 32416
rect 21508 32376 21514 32388
rect 19291 32320 19325 32348
rect 19996 32320 20300 32348
rect 19291 32317 19303 32320
rect 19245 32311 19303 32317
rect 16172 32252 17356 32280
rect 16172 32240 16178 32252
rect 17586 32240 17592 32292
rect 17644 32280 17650 32292
rect 19996 32280 20024 32320
rect 21358 32308 21364 32360
rect 21416 32308 21422 32360
rect 21928 32348 21956 32388
rect 22373 32385 22385 32388
rect 22419 32385 22431 32419
rect 22373 32379 22431 32385
rect 22554 32376 22560 32428
rect 22612 32416 22618 32428
rect 23017 32419 23075 32425
rect 23017 32416 23029 32419
rect 22612 32388 23029 32416
rect 22612 32376 22618 32388
rect 23017 32385 23029 32388
rect 23063 32385 23075 32419
rect 23017 32379 23075 32385
rect 24857 32419 24915 32425
rect 24857 32385 24869 32419
rect 24903 32416 24915 32419
rect 25317 32419 25375 32425
rect 25317 32416 25329 32419
rect 24903 32388 25329 32416
rect 24903 32385 24915 32388
rect 24857 32379 24915 32385
rect 25317 32385 25329 32388
rect 25363 32416 25375 32419
rect 25406 32416 25412 32428
rect 25363 32388 25412 32416
rect 25363 32385 25375 32388
rect 25317 32379 25375 32385
rect 25406 32376 25412 32388
rect 25464 32376 25470 32428
rect 23293 32351 23351 32357
rect 23293 32348 23305 32351
rect 21928 32320 23305 32348
rect 23293 32317 23305 32320
rect 23339 32317 23351 32351
rect 23293 32311 23351 32317
rect 17644 32252 20024 32280
rect 17644 32240 17650 32252
rect 25130 32240 25136 32292
rect 25188 32240 25194 32292
rect 10413 32215 10471 32221
rect 10413 32212 10425 32215
rect 9646 32184 10425 32212
rect 10413 32181 10425 32184
rect 10459 32212 10471 32215
rect 10962 32212 10968 32224
rect 10459 32184 10968 32212
rect 10459 32181 10471 32184
rect 10413 32175 10471 32181
rect 10962 32172 10968 32184
rect 11020 32172 11026 32224
rect 12342 32172 12348 32224
rect 12400 32212 12406 32224
rect 13446 32212 13452 32224
rect 12400 32184 13452 32212
rect 12400 32172 12406 32184
rect 13446 32172 13452 32184
rect 13504 32172 13510 32224
rect 14550 32172 14556 32224
rect 14608 32212 14614 32224
rect 15194 32212 15200 32224
rect 14608 32184 15200 32212
rect 14608 32172 14614 32184
rect 15194 32172 15200 32184
rect 15252 32172 15258 32224
rect 16666 32172 16672 32224
rect 16724 32212 16730 32224
rect 16853 32215 16911 32221
rect 16853 32212 16865 32215
rect 16724 32184 16865 32212
rect 16724 32172 16730 32184
rect 16853 32181 16865 32184
rect 16899 32181 16911 32215
rect 16853 32175 16911 32181
rect 18049 32215 18107 32221
rect 18049 32181 18061 32215
rect 18095 32212 18107 32215
rect 18322 32212 18328 32224
rect 18095 32184 18328 32212
rect 18095 32181 18107 32184
rect 18049 32175 18107 32181
rect 18322 32172 18328 32184
rect 18380 32172 18386 32224
rect 20073 32215 20131 32221
rect 20073 32181 20085 32215
rect 20119 32212 20131 32215
rect 20622 32212 20628 32224
rect 20119 32184 20628 32212
rect 20119 32181 20131 32184
rect 20073 32175 20131 32181
rect 20622 32172 20628 32184
rect 20680 32172 20686 32224
rect 20717 32215 20775 32221
rect 20717 32181 20729 32215
rect 20763 32212 20775 32215
rect 20990 32212 20996 32224
rect 20763 32184 20996 32212
rect 20763 32181 20775 32184
rect 20717 32175 20775 32181
rect 20990 32172 20996 32184
rect 21048 32172 21054 32224
rect 21358 32172 21364 32224
rect 21416 32212 21422 32224
rect 21542 32212 21548 32224
rect 21416 32184 21548 32212
rect 21416 32172 21422 32184
rect 21542 32172 21548 32184
rect 21600 32172 21606 32224
rect 22189 32215 22247 32221
rect 22189 32181 22201 32215
rect 22235 32212 22247 32215
rect 22554 32212 22560 32224
rect 22235 32184 22560 32212
rect 22235 32181 22247 32184
rect 22189 32175 22247 32181
rect 22554 32172 22560 32184
rect 22612 32172 22618 32224
rect 22738 32172 22744 32224
rect 22796 32212 22802 32224
rect 22833 32215 22891 32221
rect 22833 32212 22845 32215
rect 22796 32184 22845 32212
rect 22796 32172 22802 32184
rect 22833 32181 22845 32184
rect 22879 32181 22891 32215
rect 22833 32175 22891 32181
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 7929 32011 7987 32017
rect 7929 31977 7941 32011
rect 7975 32008 7987 32011
rect 8294 32008 8300 32020
rect 7975 31980 8300 32008
rect 7975 31977 7987 31980
rect 7929 31971 7987 31977
rect 8294 31968 8300 31980
rect 8352 31968 8358 32020
rect 8386 31968 8392 32020
rect 8444 31968 8450 32020
rect 8573 32011 8631 32017
rect 8573 31977 8585 32011
rect 8619 32008 8631 32011
rect 9122 32008 9128 32020
rect 8619 31980 9128 32008
rect 8619 31977 8631 31980
rect 8573 31971 8631 31977
rect 8588 31940 8616 31971
rect 9122 31968 9128 31980
rect 9180 31968 9186 32020
rect 9398 31968 9404 32020
rect 9456 32008 9462 32020
rect 9674 32008 9680 32020
rect 9456 31980 9680 32008
rect 9456 31968 9462 31980
rect 9674 31968 9680 31980
rect 9732 31968 9738 32020
rect 10134 31968 10140 32020
rect 10192 32008 10198 32020
rect 11149 32011 11207 32017
rect 11149 32008 11161 32011
rect 10192 31980 11161 32008
rect 10192 31968 10198 31980
rect 11149 31977 11161 31980
rect 11195 31977 11207 32011
rect 11149 31971 11207 31977
rect 11882 31968 11888 32020
rect 11940 32008 11946 32020
rect 16393 32011 16451 32017
rect 16393 32008 16405 32011
rect 11940 31980 16405 32008
rect 11940 31968 11946 31980
rect 16393 31977 16405 31980
rect 16439 31977 16451 32011
rect 16393 31971 16451 31977
rect 17586 31968 17592 32020
rect 17644 32008 17650 32020
rect 18049 32011 18107 32017
rect 18049 32008 18061 32011
rect 17644 31980 18061 32008
rect 17644 31968 17650 31980
rect 18049 31977 18061 31980
rect 18095 32008 18107 32011
rect 18230 32008 18236 32020
rect 18095 31980 18236 32008
rect 18095 31977 18107 31980
rect 18049 31971 18107 31977
rect 18230 31968 18236 31980
rect 18288 31968 18294 32020
rect 18598 31968 18604 32020
rect 18656 32008 18662 32020
rect 18656 31980 20116 32008
rect 18656 31968 18662 31980
rect 7576 31912 8616 31940
rect 6178 31832 6184 31884
rect 6236 31832 6242 31884
rect 6457 31875 6515 31881
rect 6457 31841 6469 31875
rect 6503 31872 6515 31875
rect 7190 31872 7196 31884
rect 6503 31844 7196 31872
rect 6503 31841 6515 31844
rect 6457 31835 6515 31841
rect 7190 31832 7196 31844
rect 7248 31832 7254 31884
rect 7576 31790 7604 31912
rect 9306 31900 9312 31952
rect 9364 31940 9370 31952
rect 9364 31912 9444 31940
rect 9364 31900 9370 31912
rect 9416 31872 9444 31912
rect 12158 31900 12164 31952
rect 12216 31940 12222 31952
rect 13633 31943 13691 31949
rect 13633 31940 13645 31943
rect 12216 31912 13645 31940
rect 12216 31900 12222 31912
rect 13633 31909 13645 31912
rect 13679 31940 13691 31943
rect 13814 31940 13820 31952
rect 13679 31912 13820 31940
rect 13679 31909 13691 31912
rect 13633 31903 13691 31909
rect 13814 31900 13820 31912
rect 13872 31900 13878 31952
rect 13906 31900 13912 31952
rect 13964 31940 13970 31952
rect 13964 31912 14136 31940
rect 13964 31900 13970 31912
rect 9677 31875 9735 31881
rect 9677 31872 9689 31875
rect 9416 31844 9689 31872
rect 9677 31841 9689 31844
rect 9723 31872 9735 31875
rect 9766 31872 9772 31884
rect 9723 31844 9772 31872
rect 9723 31841 9735 31844
rect 9677 31835 9735 31841
rect 9766 31832 9772 31844
rect 9824 31832 9830 31884
rect 9390 31807 9448 31813
rect 9390 31804 9402 31807
rect 9324 31776 9402 31804
rect 9324 31736 9352 31776
rect 9390 31773 9402 31776
rect 9436 31773 9448 31807
rect 14108 31804 14136 31912
rect 14182 31900 14188 31952
rect 14240 31940 14246 31952
rect 14277 31943 14335 31949
rect 14277 31940 14289 31943
rect 14240 31912 14289 31940
rect 14240 31900 14246 31912
rect 14277 31909 14289 31912
rect 14323 31909 14335 31943
rect 18782 31940 18788 31952
rect 14277 31903 14335 31909
rect 14752 31912 18788 31940
rect 14752 31881 14780 31912
rect 18782 31900 18788 31912
rect 18840 31900 18846 31952
rect 19426 31900 19432 31952
rect 19484 31900 19490 31952
rect 19886 31900 19892 31952
rect 19944 31940 19950 31952
rect 19944 31912 20024 31940
rect 19944 31900 19950 31912
rect 14737 31875 14795 31881
rect 14737 31841 14749 31875
rect 14783 31841 14795 31875
rect 14737 31835 14795 31841
rect 14829 31875 14887 31881
rect 14829 31841 14841 31875
rect 14875 31841 14887 31875
rect 14829 31835 14887 31841
rect 14844 31804 14872 31835
rect 15102 31832 15108 31884
rect 15160 31872 15166 31884
rect 19996 31881 20024 31912
rect 16945 31875 17003 31881
rect 16945 31872 16957 31875
rect 15160 31844 16957 31872
rect 15160 31832 15166 31844
rect 16945 31841 16957 31844
rect 16991 31841 17003 31875
rect 19981 31875 20039 31881
rect 16945 31835 17003 31841
rect 17328 31844 19748 31872
rect 14108 31776 14872 31804
rect 9390 31767 9448 31773
rect 15654 31764 15660 31816
rect 15712 31804 15718 31816
rect 16758 31804 16764 31816
rect 15712 31776 16764 31804
rect 15712 31764 15718 31776
rect 16758 31764 16764 31776
rect 16816 31764 16822 31816
rect 9582 31736 9588 31748
rect 9324 31708 9588 31736
rect 9582 31696 9588 31708
rect 9640 31696 9646 31748
rect 10962 31736 10968 31748
rect 10902 31708 10968 31736
rect 10962 31696 10968 31708
rect 11020 31736 11026 31748
rect 16853 31739 16911 31745
rect 11020 31708 11560 31736
rect 11020 31696 11026 31708
rect 9122 31628 9128 31680
rect 9180 31628 9186 31680
rect 11532 31677 11560 31708
rect 16853 31705 16865 31739
rect 16899 31736 16911 31739
rect 17328 31736 17356 31844
rect 16899 31708 17356 31736
rect 16899 31705 16911 31708
rect 16853 31699 16911 31705
rect 17402 31696 17408 31748
rect 17460 31736 17466 31748
rect 18417 31739 18475 31745
rect 18417 31736 18429 31739
rect 17460 31708 18429 31736
rect 17460 31696 17466 31708
rect 18417 31705 18429 31708
rect 18463 31736 18475 31739
rect 18874 31736 18880 31748
rect 18463 31708 18880 31736
rect 18463 31705 18475 31708
rect 18417 31699 18475 31705
rect 18874 31696 18880 31708
rect 18932 31696 18938 31748
rect 11517 31671 11575 31677
rect 11517 31637 11529 31671
rect 11563 31668 11575 31671
rect 11698 31668 11704 31680
rect 11563 31640 11704 31668
rect 11563 31637 11575 31640
rect 11517 31631 11575 31637
rect 11698 31628 11704 31640
rect 11756 31628 11762 31680
rect 12434 31628 12440 31680
rect 12492 31668 12498 31680
rect 12710 31668 12716 31680
rect 12492 31640 12716 31668
rect 12492 31628 12498 31640
rect 12710 31628 12716 31640
rect 12768 31628 12774 31680
rect 13814 31628 13820 31680
rect 13872 31668 13878 31680
rect 14645 31671 14703 31677
rect 14645 31668 14657 31671
rect 13872 31640 14657 31668
rect 13872 31628 13878 31640
rect 14645 31637 14657 31640
rect 14691 31668 14703 31671
rect 14918 31668 14924 31680
rect 14691 31640 14924 31668
rect 14691 31637 14703 31640
rect 14645 31631 14703 31637
rect 14918 31628 14924 31640
rect 14976 31628 14982 31680
rect 16761 31671 16819 31677
rect 16761 31637 16773 31671
rect 16807 31668 16819 31671
rect 17218 31668 17224 31680
rect 16807 31640 17224 31668
rect 16807 31637 16819 31640
rect 16761 31631 16819 31637
rect 17218 31628 17224 31640
rect 17276 31628 17282 31680
rect 18230 31668 18236 31680
rect 18191 31640 18236 31668
rect 18230 31628 18236 31640
rect 18288 31668 18294 31680
rect 19150 31668 19156 31680
rect 18288 31640 19156 31668
rect 18288 31628 18294 31640
rect 19150 31628 19156 31640
rect 19208 31628 19214 31680
rect 19720 31668 19748 31844
rect 19981 31841 19993 31875
rect 20027 31841 20039 31875
rect 20088 31872 20116 31980
rect 22554 31968 22560 32020
rect 22612 32008 22618 32020
rect 24302 32008 24308 32020
rect 22612 31980 24308 32008
rect 22612 31968 22618 31980
rect 24302 31968 24308 31980
rect 24360 31968 24366 32020
rect 20254 31900 20260 31952
rect 20312 31940 20318 31952
rect 20625 31943 20683 31949
rect 20625 31940 20637 31943
rect 20312 31912 20637 31940
rect 20312 31900 20318 31912
rect 20625 31909 20637 31912
rect 20671 31909 20683 31943
rect 20625 31903 20683 31909
rect 20990 31900 20996 31952
rect 21048 31940 21054 31952
rect 21913 31943 21971 31949
rect 21048 31912 21588 31940
rect 21048 31900 21054 31912
rect 21177 31875 21235 31881
rect 21177 31872 21189 31875
rect 20088 31844 21189 31872
rect 19981 31835 20039 31841
rect 21177 31841 21189 31844
rect 21223 31841 21235 31875
rect 21560 31872 21588 31912
rect 21913 31909 21925 31943
rect 21959 31940 21971 31943
rect 23382 31940 23388 31952
rect 21959 31912 23388 31940
rect 21959 31909 21971 31912
rect 21913 31903 21971 31909
rect 23382 31900 23388 31912
rect 23440 31900 23446 31952
rect 23566 31900 23572 31952
rect 23624 31940 23630 31952
rect 25133 31943 25191 31949
rect 25133 31940 25145 31943
rect 23624 31912 25145 31940
rect 23624 31900 23630 31912
rect 25133 31909 25145 31912
rect 25179 31909 25191 31943
rect 25133 31903 25191 31909
rect 22373 31875 22431 31881
rect 22373 31872 22385 31875
rect 21560 31844 22385 31872
rect 21177 31835 21235 31841
rect 22373 31841 22385 31844
rect 22419 31841 22431 31875
rect 22373 31835 22431 31841
rect 22557 31875 22615 31881
rect 22557 31841 22569 31875
rect 22603 31872 22615 31875
rect 23474 31872 23480 31884
rect 22603 31844 23480 31872
rect 22603 31841 22615 31844
rect 22557 31835 22615 31841
rect 23474 31832 23480 31844
rect 23532 31832 23538 31884
rect 19889 31807 19947 31813
rect 19889 31773 19901 31807
rect 19935 31804 19947 31807
rect 20898 31804 20904 31816
rect 19935 31776 20904 31804
rect 19935 31773 19947 31776
rect 19889 31767 19947 31773
rect 20898 31764 20904 31776
rect 20956 31764 20962 31816
rect 21085 31807 21143 31813
rect 21085 31773 21097 31807
rect 21131 31804 21143 31807
rect 21634 31804 21640 31816
rect 21131 31776 21640 31804
rect 21131 31773 21143 31776
rect 21085 31767 21143 31773
rect 21634 31764 21640 31776
rect 21692 31764 21698 31816
rect 23934 31764 23940 31816
rect 23992 31804 23998 31816
rect 24029 31807 24087 31813
rect 24029 31804 24041 31807
rect 23992 31776 24041 31804
rect 23992 31764 23998 31776
rect 24029 31773 24041 31776
rect 24075 31773 24087 31807
rect 24029 31767 24087 31773
rect 24857 31807 24915 31813
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 25314 31804 25320 31816
rect 24903 31776 25320 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 19797 31739 19855 31745
rect 19797 31705 19809 31739
rect 19843 31736 19855 31739
rect 20714 31736 20720 31748
rect 19843 31708 20720 31736
rect 19843 31705 19855 31708
rect 19797 31699 19855 31705
rect 20714 31696 20720 31708
rect 20772 31696 20778 31748
rect 20993 31739 21051 31745
rect 20993 31705 21005 31739
rect 21039 31736 21051 31739
rect 21818 31736 21824 31748
rect 21039 31708 21824 31736
rect 21039 31705 21051 31708
rect 20993 31699 21051 31705
rect 21008 31668 21036 31699
rect 21818 31696 21824 31708
rect 21876 31696 21882 31748
rect 22278 31696 22284 31748
rect 22336 31696 22342 31748
rect 19720 31640 21036 31668
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 7469 31467 7527 31473
rect 7469 31433 7481 31467
rect 7515 31464 7527 31467
rect 7650 31464 7656 31476
rect 7515 31436 7656 31464
rect 7515 31433 7527 31436
rect 7469 31427 7527 31433
rect 7650 31424 7656 31436
rect 7708 31424 7714 31476
rect 8662 31424 8668 31476
rect 8720 31424 8726 31476
rect 9033 31467 9091 31473
rect 9033 31433 9045 31467
rect 9079 31464 9091 31467
rect 9858 31464 9864 31476
rect 9079 31436 9864 31464
rect 9079 31433 9091 31436
rect 9033 31427 9091 31433
rect 9858 31424 9864 31436
rect 9916 31424 9922 31476
rect 12710 31424 12716 31476
rect 12768 31464 12774 31476
rect 13354 31464 13360 31476
rect 12768 31436 13360 31464
rect 12768 31424 12774 31436
rect 13354 31424 13360 31436
rect 13412 31424 13418 31476
rect 14642 31424 14648 31476
rect 14700 31464 14706 31476
rect 16206 31464 16212 31476
rect 14700 31436 16212 31464
rect 14700 31424 14706 31436
rect 16206 31424 16212 31436
rect 16264 31424 16270 31476
rect 17310 31424 17316 31476
rect 17368 31464 17374 31476
rect 18325 31467 18383 31473
rect 18325 31464 18337 31467
rect 17368 31436 18337 31464
rect 17368 31424 17374 31436
rect 18325 31433 18337 31436
rect 18371 31433 18383 31467
rect 18325 31427 18383 31433
rect 19521 31467 19579 31473
rect 19521 31433 19533 31467
rect 19567 31464 19579 31467
rect 21450 31464 21456 31476
rect 19567 31436 21456 31464
rect 19567 31433 19579 31436
rect 19521 31427 19579 31433
rect 21450 31424 21456 31436
rect 21508 31424 21514 31476
rect 21545 31467 21603 31473
rect 21545 31433 21557 31467
rect 21591 31464 21603 31467
rect 21634 31464 21640 31476
rect 21591 31436 21640 31464
rect 21591 31433 21603 31436
rect 21545 31427 21603 31433
rect 21634 31424 21640 31436
rect 21692 31424 21698 31476
rect 23290 31424 23296 31476
rect 23348 31464 23354 31476
rect 25133 31467 25191 31473
rect 25133 31464 25145 31467
rect 23348 31436 25145 31464
rect 23348 31424 23354 31436
rect 25133 31433 25145 31436
rect 25179 31433 25191 31467
rect 25133 31427 25191 31433
rect 9674 31396 9680 31408
rect 8128 31368 9680 31396
rect 1765 31331 1823 31337
rect 1765 31297 1777 31331
rect 1811 31328 1823 31331
rect 1946 31328 1952 31340
rect 1811 31300 1952 31328
rect 1811 31297 1823 31300
rect 1765 31291 1823 31297
rect 1946 31288 1952 31300
rect 2004 31288 2010 31340
rect 7834 31288 7840 31340
rect 7892 31288 7898 31340
rect 1302 31220 1308 31272
rect 1360 31260 1366 31272
rect 8128 31269 8156 31368
rect 9674 31356 9680 31368
rect 9732 31396 9738 31408
rect 11330 31396 11336 31408
rect 9732 31368 11336 31396
rect 9732 31356 9738 31368
rect 11330 31356 11336 31368
rect 11388 31356 11394 31408
rect 15378 31356 15384 31408
rect 15436 31396 15442 31408
rect 19889 31399 19947 31405
rect 19889 31396 19901 31399
rect 15436 31368 19901 31396
rect 15436 31356 15442 31368
rect 19889 31365 19901 31368
rect 19935 31396 19947 31399
rect 20533 31399 20591 31405
rect 20533 31396 20545 31399
rect 19935 31368 20545 31396
rect 19935 31365 19947 31368
rect 19889 31359 19947 31365
rect 20533 31365 20545 31368
rect 20579 31365 20591 31399
rect 20533 31359 20591 31365
rect 20622 31356 20628 31408
rect 20680 31396 20686 31408
rect 21358 31396 21364 31408
rect 20680 31368 21364 31396
rect 20680 31356 20686 31368
rect 21358 31356 21364 31368
rect 21416 31356 21422 31408
rect 22465 31399 22523 31405
rect 22465 31396 22477 31399
rect 21560 31368 22477 31396
rect 21560 31340 21588 31368
rect 22465 31365 22477 31368
rect 22511 31365 22523 31399
rect 23934 31396 23940 31408
rect 23690 31368 23940 31396
rect 22465 31359 22523 31365
rect 23934 31356 23940 31368
rect 23992 31356 23998 31408
rect 8754 31288 8760 31340
rect 8812 31328 8818 31340
rect 8812 31300 9260 31328
rect 8812 31288 8818 31300
rect 9232 31269 9260 31300
rect 9582 31288 9588 31340
rect 9640 31328 9646 31340
rect 9640 31300 12940 31328
rect 9640 31288 9646 31300
rect 12912 31269 12940 31300
rect 14274 31288 14280 31340
rect 14332 31328 14338 31340
rect 15013 31331 15071 31337
rect 15013 31328 15025 31331
rect 14332 31300 15025 31328
rect 14332 31288 14338 31300
rect 15013 31297 15025 31300
rect 15059 31328 15071 31331
rect 15930 31328 15936 31340
rect 15059 31300 15936 31328
rect 15059 31297 15071 31300
rect 15013 31291 15071 31297
rect 15930 31288 15936 31300
rect 15988 31288 15994 31340
rect 17497 31331 17555 31337
rect 17497 31328 17509 31331
rect 16776 31300 17509 31328
rect 2041 31263 2099 31269
rect 2041 31260 2053 31263
rect 1360 31232 2053 31260
rect 1360 31220 1366 31232
rect 2041 31229 2053 31232
rect 2087 31229 2099 31263
rect 2041 31223 2099 31229
rect 7929 31263 7987 31269
rect 7929 31229 7941 31263
rect 7975 31229 7987 31263
rect 7929 31223 7987 31229
rect 8113 31263 8171 31269
rect 8113 31229 8125 31263
rect 8159 31229 8171 31263
rect 8113 31223 8171 31229
rect 9125 31263 9183 31269
rect 9125 31229 9137 31263
rect 9171 31229 9183 31263
rect 9125 31223 9183 31229
rect 9217 31263 9275 31269
rect 9217 31229 9229 31263
rect 9263 31260 9275 31263
rect 9677 31263 9735 31269
rect 9677 31260 9689 31263
rect 9263 31232 9689 31260
rect 9263 31229 9275 31232
rect 9217 31223 9275 31229
rect 9677 31229 9689 31232
rect 9723 31229 9735 31263
rect 9677 31223 9735 31229
rect 12897 31263 12955 31269
rect 12897 31229 12909 31263
rect 12943 31229 12955 31263
rect 12897 31223 12955 31229
rect 13173 31263 13231 31269
rect 13173 31229 13185 31263
rect 13219 31260 13231 31263
rect 13262 31260 13268 31272
rect 13219 31232 13268 31260
rect 13219 31229 13231 31232
rect 13173 31223 13231 31229
rect 4798 31152 4804 31204
rect 4856 31192 4862 31204
rect 7193 31195 7251 31201
rect 7193 31192 7205 31195
rect 4856 31164 7205 31192
rect 4856 31152 4862 31164
rect 7193 31161 7205 31164
rect 7239 31192 7251 31195
rect 7944 31192 7972 31223
rect 8662 31192 8668 31204
rect 7239 31164 8668 31192
rect 7239 31161 7251 31164
rect 7193 31155 7251 31161
rect 8662 31152 8668 31164
rect 8720 31152 8726 31204
rect 8754 31152 8760 31204
rect 8812 31192 8818 31204
rect 9140 31192 9168 31223
rect 8812 31164 9168 31192
rect 8812 31152 8818 31164
rect 5718 31084 5724 31136
rect 5776 31124 5782 31136
rect 8772 31124 8800 31152
rect 5776 31096 8800 31124
rect 12912 31124 12940 31223
rect 13262 31220 13268 31232
rect 13320 31260 13326 31272
rect 13538 31260 13544 31272
rect 13320 31232 13544 31260
rect 13320 31220 13326 31232
rect 13538 31220 13544 31232
rect 13596 31220 13602 31272
rect 14458 31124 14464 31136
rect 12912 31096 14464 31124
rect 5776 31084 5782 31096
rect 14458 31084 14464 31096
rect 14516 31084 14522 31136
rect 15286 31084 15292 31136
rect 15344 31124 15350 31136
rect 16776 31133 16804 31300
rect 17497 31297 17509 31300
rect 17543 31297 17555 31331
rect 17497 31291 17555 31297
rect 17589 31331 17647 31337
rect 17589 31297 17601 31331
rect 17635 31328 17647 31331
rect 18693 31331 18751 31337
rect 17635 31300 18276 31328
rect 17635 31297 17647 31300
rect 17589 31291 17647 31297
rect 17034 31220 17040 31272
rect 17092 31260 17098 31272
rect 17681 31263 17739 31269
rect 17681 31260 17693 31263
rect 17092 31232 17693 31260
rect 17092 31220 17098 31232
rect 17604 31204 17632 31232
rect 17681 31229 17693 31232
rect 17727 31229 17739 31263
rect 17681 31223 17739 31229
rect 17586 31152 17592 31204
rect 17644 31152 17650 31204
rect 16761 31127 16819 31133
rect 16761 31124 16773 31127
rect 15344 31096 16773 31124
rect 15344 31084 15350 31096
rect 16761 31093 16773 31096
rect 16807 31093 16819 31127
rect 16761 31087 16819 31093
rect 17126 31084 17132 31136
rect 17184 31084 17190 31136
rect 18248 31124 18276 31300
rect 18693 31297 18705 31331
rect 18739 31328 18751 31331
rect 19242 31328 19248 31340
rect 18739 31300 19248 31328
rect 18739 31297 18751 31300
rect 18693 31291 18751 31297
rect 19242 31288 19248 31300
rect 19300 31288 19306 31340
rect 20717 31331 20775 31337
rect 20717 31328 20729 31331
rect 19996 31300 20729 31328
rect 19996 31272 20024 31300
rect 20717 31297 20729 31300
rect 20763 31297 20775 31331
rect 20717 31291 20775 31297
rect 21542 31288 21548 31340
rect 21600 31288 21606 31340
rect 24394 31288 24400 31340
rect 24452 31328 24458 31340
rect 24581 31331 24639 31337
rect 24581 31328 24593 31331
rect 24452 31300 24593 31328
rect 24452 31288 24458 31300
rect 24581 31297 24593 31300
rect 24627 31297 24639 31331
rect 24581 31291 24639 31297
rect 25314 31288 25320 31340
rect 25372 31288 25378 31340
rect 18785 31263 18843 31269
rect 18785 31229 18797 31263
rect 18831 31229 18843 31263
rect 18785 31223 18843 31229
rect 18800 31192 18828 31223
rect 18874 31220 18880 31272
rect 18932 31220 18938 31272
rect 19978 31220 19984 31272
rect 20036 31220 20042 31272
rect 20165 31263 20223 31269
rect 20165 31229 20177 31263
rect 20211 31260 20223 31263
rect 20211 31232 20668 31260
rect 20211 31229 20223 31232
rect 20165 31223 20223 31229
rect 20438 31192 20444 31204
rect 18800 31164 20444 31192
rect 20438 31152 20444 31164
rect 20496 31152 20502 31204
rect 20640 31136 20668 31232
rect 22186 31220 22192 31272
rect 22244 31220 22250 31272
rect 19150 31124 19156 31136
rect 18248 31096 19156 31124
rect 19150 31084 19156 31096
rect 19208 31084 19214 31136
rect 20162 31084 20168 31136
rect 20220 31124 20226 31136
rect 20346 31124 20352 31136
rect 20220 31096 20352 31124
rect 20220 31084 20226 31096
rect 20346 31084 20352 31096
rect 20404 31084 20410 31136
rect 20622 31084 20628 31136
rect 20680 31124 20686 31136
rect 22646 31124 22652 31136
rect 20680 31096 22652 31124
rect 20680 31084 20686 31096
rect 22646 31084 22652 31096
rect 22704 31084 22710 31136
rect 23566 31084 23572 31136
rect 23624 31124 23630 31136
rect 23937 31127 23995 31133
rect 23937 31124 23949 31127
rect 23624 31096 23949 31124
rect 23624 31084 23630 31096
rect 23937 31093 23949 31096
rect 23983 31093 23995 31127
rect 23937 31087 23995 31093
rect 24394 31084 24400 31136
rect 24452 31084 24458 31136
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 12618 30880 12624 30932
rect 12676 30920 12682 30932
rect 12805 30923 12863 30929
rect 12805 30920 12817 30923
rect 12676 30892 12817 30920
rect 12676 30880 12682 30892
rect 12805 30889 12817 30892
rect 12851 30889 12863 30923
rect 18690 30920 18696 30932
rect 12805 30883 12863 30889
rect 14752 30892 18696 30920
rect 11698 30852 11704 30864
rect 10980 30824 11704 30852
rect 1854 30744 1860 30796
rect 1912 30784 1918 30796
rect 4065 30787 4123 30793
rect 4065 30784 4077 30787
rect 1912 30756 4077 30784
rect 1912 30744 1918 30756
rect 4065 30753 4077 30756
rect 4111 30753 4123 30787
rect 4065 30747 4123 30753
rect 4614 30744 4620 30796
rect 4672 30744 4678 30796
rect 7834 30744 7840 30796
rect 7892 30784 7898 30796
rect 7929 30787 7987 30793
rect 7929 30784 7941 30787
rect 7892 30756 7941 30784
rect 7892 30744 7898 30756
rect 7929 30753 7941 30756
rect 7975 30753 7987 30787
rect 7929 30747 7987 30753
rect 9582 30744 9588 30796
rect 9640 30744 9646 30796
rect 9861 30787 9919 30793
rect 9861 30753 9873 30787
rect 9907 30784 9919 30787
rect 10870 30784 10876 30796
rect 9907 30756 10876 30784
rect 9907 30753 9919 30756
rect 9861 30747 9919 30753
rect 10870 30744 10876 30756
rect 10928 30744 10934 30796
rect 10980 30702 11008 30824
rect 11698 30812 11704 30824
rect 11756 30852 11762 30864
rect 14274 30852 14280 30864
rect 11756 30824 14280 30852
rect 11756 30812 11762 30824
rect 14274 30812 14280 30824
rect 14332 30812 14338 30864
rect 11330 30744 11336 30796
rect 11388 30784 11394 30796
rect 12529 30787 12587 30793
rect 12529 30784 12541 30787
rect 11388 30756 12541 30784
rect 11388 30744 11394 30756
rect 12529 30753 12541 30756
rect 12575 30784 12587 30787
rect 13357 30787 13415 30793
rect 13357 30784 13369 30787
rect 12575 30756 13369 30784
rect 12575 30753 12587 30756
rect 12529 30747 12587 30753
rect 13357 30753 13369 30756
rect 13403 30753 13415 30787
rect 13357 30747 13415 30753
rect 11422 30676 11428 30728
rect 11480 30716 11486 30728
rect 12253 30719 12311 30725
rect 12253 30716 12265 30719
rect 11480 30688 12265 30716
rect 11480 30676 11486 30688
rect 12253 30685 12265 30688
rect 12299 30716 12311 30719
rect 13173 30719 13231 30725
rect 13173 30716 13185 30719
rect 12299 30688 13185 30716
rect 12299 30685 12311 30688
rect 12253 30679 12311 30685
rect 13173 30685 13185 30688
rect 13219 30716 13231 30719
rect 14752 30716 14780 30892
rect 18690 30880 18696 30892
rect 18748 30880 18754 30932
rect 19610 30880 19616 30932
rect 19668 30920 19674 30932
rect 20346 30920 20352 30932
rect 19668 30892 20352 30920
rect 19668 30880 19674 30892
rect 20346 30880 20352 30892
rect 20404 30920 20410 30932
rect 24857 30923 24915 30929
rect 20404 30892 22094 30920
rect 20404 30880 20410 30892
rect 15930 30812 15936 30864
rect 15988 30812 15994 30864
rect 17678 30812 17684 30864
rect 17736 30852 17742 30864
rect 18233 30855 18291 30861
rect 18233 30852 18245 30855
rect 17736 30824 18245 30852
rect 17736 30812 17742 30824
rect 18233 30821 18245 30824
rect 18279 30821 18291 30855
rect 20441 30855 20499 30861
rect 20441 30852 20453 30855
rect 18233 30815 18291 30821
rect 19904 30824 20453 30852
rect 19904 30796 19932 30824
rect 20441 30821 20453 30824
rect 20487 30821 20499 30855
rect 22066 30852 22094 30892
rect 24857 30889 24869 30923
rect 24903 30920 24915 30923
rect 25314 30920 25320 30932
rect 24903 30892 25320 30920
rect 24903 30889 24915 30892
rect 24857 30883 24915 30889
rect 25314 30880 25320 30892
rect 25372 30880 25378 30932
rect 25133 30855 25191 30861
rect 25133 30852 25145 30855
rect 22066 30824 25145 30852
rect 20441 30815 20499 30821
rect 25133 30821 25145 30824
rect 25179 30821 25191 30855
rect 25133 30815 25191 30821
rect 15194 30744 15200 30796
rect 15252 30784 15258 30796
rect 16209 30787 16267 30793
rect 16209 30784 16221 30787
rect 15252 30756 16221 30784
rect 15252 30744 15258 30756
rect 16209 30753 16221 30756
rect 16255 30753 16267 30787
rect 16209 30747 16267 30753
rect 16482 30744 16488 30796
rect 16540 30784 16546 30796
rect 19058 30784 19064 30796
rect 16540 30756 19064 30784
rect 16540 30744 16546 30756
rect 19058 30744 19064 30756
rect 19116 30744 19122 30796
rect 19886 30744 19892 30796
rect 19944 30744 19950 30796
rect 19978 30744 19984 30796
rect 20036 30744 20042 30796
rect 20530 30744 20536 30796
rect 20588 30784 20594 30796
rect 22557 30787 22615 30793
rect 22557 30784 22569 30787
rect 20588 30756 22569 30784
rect 20588 30744 20594 30756
rect 22557 30753 22569 30756
rect 22603 30753 22615 30787
rect 22557 30747 22615 30753
rect 13219 30688 14780 30716
rect 13219 30685 13231 30688
rect 13173 30679 13231 30685
rect 15470 30676 15476 30728
rect 15528 30716 15534 30728
rect 15930 30716 15936 30728
rect 15528 30688 15936 30716
rect 15528 30676 15534 30688
rect 15930 30676 15936 30688
rect 15988 30716 15994 30728
rect 19797 30719 19855 30725
rect 15988 30688 16252 30716
rect 15988 30676 15994 30688
rect 3786 30608 3792 30660
rect 3844 30648 3850 30660
rect 4157 30651 4215 30657
rect 4157 30648 4169 30651
rect 3844 30620 4169 30648
rect 3844 30608 3850 30620
rect 4157 30617 4169 30620
rect 4203 30617 4215 30651
rect 4157 30611 4215 30617
rect 13265 30651 13323 30657
rect 13265 30617 13277 30651
rect 13311 30648 13323 30651
rect 13909 30651 13967 30657
rect 13909 30648 13921 30651
rect 13311 30620 13921 30648
rect 13311 30617 13323 30620
rect 13265 30611 13323 30617
rect 13909 30617 13921 30620
rect 13955 30648 13967 30651
rect 16114 30648 16120 30660
rect 13955 30620 16120 30648
rect 13955 30617 13967 30620
rect 13909 30611 13967 30617
rect 16114 30608 16120 30620
rect 16172 30608 16178 30660
rect 16224 30648 16252 30688
rect 19797 30685 19809 30719
rect 19843 30716 19855 30719
rect 20070 30716 20076 30728
rect 19843 30688 20076 30716
rect 19843 30685 19855 30688
rect 19797 30679 19855 30685
rect 20070 30676 20076 30688
rect 20128 30676 20134 30728
rect 20438 30676 20444 30728
rect 20496 30716 20502 30728
rect 20496 30688 22094 30716
rect 20496 30676 20502 30688
rect 22066 30648 22094 30688
rect 22462 30676 22468 30728
rect 22520 30716 22526 30728
rect 23017 30719 23075 30725
rect 23017 30716 23029 30719
rect 22520 30688 23029 30716
rect 22520 30676 22526 30688
rect 23017 30685 23029 30688
rect 23063 30685 23075 30719
rect 23017 30679 23075 30685
rect 23842 30676 23848 30728
rect 23900 30676 23906 30728
rect 25317 30719 25375 30725
rect 25317 30685 25329 30719
rect 25363 30716 25375 30719
rect 25498 30716 25504 30728
rect 25363 30688 25504 30716
rect 25363 30685 25375 30688
rect 25317 30679 25375 30685
rect 25498 30676 25504 30688
rect 25556 30676 25562 30728
rect 22373 30651 22431 30657
rect 22373 30648 22385 30651
rect 16224 30620 16974 30648
rect 22066 30620 22385 30648
rect 22373 30617 22385 30620
rect 22419 30648 22431 30651
rect 24486 30648 24492 30660
rect 22419 30620 24492 30648
rect 22419 30617 22431 30620
rect 22373 30611 22431 30617
rect 24486 30608 24492 30620
rect 24544 30608 24550 30660
rect 8573 30583 8631 30589
rect 8573 30549 8585 30583
rect 8619 30580 8631 30583
rect 8754 30580 8760 30592
rect 8619 30552 8760 30580
rect 8619 30549 8631 30552
rect 8573 30543 8631 30549
rect 8754 30540 8760 30552
rect 8812 30540 8818 30592
rect 11330 30540 11336 30592
rect 11388 30540 11394 30592
rect 14090 30540 14096 30592
rect 14148 30580 14154 30592
rect 15378 30580 15384 30592
rect 14148 30552 15384 30580
rect 14148 30540 14154 30552
rect 15378 30540 15384 30552
rect 15436 30540 15442 30592
rect 17494 30540 17500 30592
rect 17552 30580 17558 30592
rect 17957 30583 18015 30589
rect 17957 30580 17969 30583
rect 17552 30552 17969 30580
rect 17552 30540 17558 30552
rect 17957 30549 17969 30552
rect 18003 30549 18015 30583
rect 17957 30543 18015 30549
rect 19426 30540 19432 30592
rect 19484 30540 19490 30592
rect 21818 30540 21824 30592
rect 21876 30580 21882 30592
rect 22005 30583 22063 30589
rect 22005 30580 22017 30583
rect 21876 30552 22017 30580
rect 21876 30540 21882 30552
rect 22005 30549 22017 30552
rect 22051 30549 22063 30583
rect 22005 30543 22063 30549
rect 23661 30583 23719 30589
rect 23661 30549 23673 30583
rect 23707 30580 23719 30583
rect 25130 30580 25136 30592
rect 23707 30552 25136 30580
rect 23707 30549 23719 30552
rect 23661 30543 23719 30549
rect 25130 30540 25136 30552
rect 25188 30540 25194 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 10042 30336 10048 30388
rect 10100 30376 10106 30388
rect 10318 30376 10324 30388
rect 10100 30348 10324 30376
rect 10100 30336 10106 30348
rect 10318 30336 10324 30348
rect 10376 30376 10382 30388
rect 10873 30379 10931 30385
rect 10873 30376 10885 30379
rect 10376 30348 10885 30376
rect 10376 30336 10382 30348
rect 10873 30345 10885 30348
rect 10919 30345 10931 30379
rect 10873 30339 10931 30345
rect 15120 30348 16068 30376
rect 6270 30268 6276 30320
rect 6328 30308 6334 30320
rect 8941 30311 8999 30317
rect 8941 30308 8953 30311
rect 6328 30280 8953 30308
rect 6328 30268 6334 30280
rect 8941 30277 8953 30280
rect 8987 30308 8999 30311
rect 9582 30308 9588 30320
rect 8987 30280 9588 30308
rect 8987 30277 8999 30280
rect 8941 30271 8999 30277
rect 9582 30268 9588 30280
rect 9640 30268 9646 30320
rect 14366 30308 14372 30320
rect 12268 30280 14372 30308
rect 10781 30243 10839 30249
rect 10781 30209 10793 30243
rect 10827 30240 10839 30243
rect 11701 30243 11759 30249
rect 11701 30240 11713 30243
rect 10827 30212 11713 30240
rect 10827 30209 10839 30212
rect 10781 30203 10839 30209
rect 11701 30209 11713 30212
rect 11747 30209 11759 30243
rect 11701 30203 11759 30209
rect 11057 30175 11115 30181
rect 11057 30141 11069 30175
rect 11103 30172 11115 30175
rect 11146 30172 11152 30184
rect 11103 30144 11152 30172
rect 11103 30141 11115 30144
rect 11057 30135 11115 30141
rect 11146 30132 11152 30144
rect 11204 30132 11210 30184
rect 10410 29996 10416 30048
rect 10468 29996 10474 30048
rect 11882 29996 11888 30048
rect 11940 30036 11946 30048
rect 12268 30045 12296 30280
rect 14366 30268 14372 30280
rect 14424 30308 14430 30320
rect 15120 30308 15148 30348
rect 14424 30280 15148 30308
rect 14424 30268 14430 30280
rect 15470 30268 15476 30320
rect 15528 30268 15534 30320
rect 14458 30200 14464 30252
rect 14516 30200 14522 30252
rect 16040 30240 16068 30348
rect 16114 30336 16120 30388
rect 16172 30376 16178 30388
rect 17954 30376 17960 30388
rect 16172 30348 17960 30376
rect 16172 30336 16178 30348
rect 17954 30336 17960 30348
rect 18012 30336 18018 30388
rect 18874 30336 18880 30388
rect 18932 30376 18938 30388
rect 21082 30376 21088 30388
rect 18932 30348 21088 30376
rect 18932 30336 18938 30348
rect 21082 30336 21088 30348
rect 21140 30336 21146 30388
rect 23934 30336 23940 30388
rect 23992 30376 23998 30388
rect 23992 30348 24992 30376
rect 23992 30336 23998 30348
rect 16298 30268 16304 30320
rect 16356 30308 16362 30320
rect 16356 30280 19656 30308
rect 16356 30268 16362 30280
rect 17957 30243 18015 30249
rect 17957 30240 17969 30243
rect 16040 30212 17969 30240
rect 17957 30209 17969 30212
rect 18003 30240 18015 30243
rect 18601 30243 18659 30249
rect 18601 30240 18613 30243
rect 18003 30212 18613 30240
rect 18003 30209 18015 30212
rect 17957 30203 18015 30209
rect 18601 30209 18613 30212
rect 18647 30209 18659 30243
rect 18601 30203 18659 30209
rect 18690 30200 18696 30252
rect 18748 30240 18754 30252
rect 19628 30249 19656 30280
rect 23566 30268 23572 30320
rect 23624 30308 23630 30320
rect 23661 30311 23719 30317
rect 23661 30308 23673 30311
rect 23624 30280 23673 30308
rect 23624 30268 23630 30280
rect 23661 30277 23673 30280
rect 23707 30277 23719 30311
rect 24964 30308 24992 30348
rect 25409 30311 25467 30317
rect 25409 30308 25421 30311
rect 24886 30280 25421 30308
rect 23661 30271 23719 30277
rect 25409 30277 25421 30280
rect 25455 30277 25467 30311
rect 25409 30271 25467 30277
rect 18785 30243 18843 30249
rect 18785 30240 18797 30243
rect 18748 30212 18797 30240
rect 18748 30200 18754 30212
rect 18785 30209 18797 30212
rect 18831 30209 18843 30243
rect 18785 30203 18843 30209
rect 19613 30243 19671 30249
rect 19613 30209 19625 30243
rect 19659 30209 19671 30243
rect 19613 30203 19671 30209
rect 22186 30200 22192 30252
rect 22244 30240 22250 30252
rect 23385 30243 23443 30249
rect 23385 30240 23397 30243
rect 22244 30212 23397 30240
rect 22244 30200 22250 30212
rect 23385 30209 23397 30212
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 12434 30132 12440 30184
rect 12492 30172 12498 30184
rect 12618 30172 12624 30184
rect 12492 30144 12624 30172
rect 12492 30132 12498 30144
rect 12618 30132 12624 30144
rect 12676 30132 12682 30184
rect 14826 30132 14832 30184
rect 14884 30172 14890 30184
rect 16206 30172 16212 30184
rect 14884 30144 16212 30172
rect 14884 30132 14890 30144
rect 16206 30132 16212 30144
rect 16264 30132 16270 30184
rect 16945 30175 17003 30181
rect 16945 30141 16957 30175
rect 16991 30172 17003 30175
rect 17218 30172 17224 30184
rect 16991 30144 17224 30172
rect 16991 30141 17003 30144
rect 16945 30135 17003 30141
rect 17218 30132 17224 30144
rect 17276 30132 17282 30184
rect 18046 30132 18052 30184
rect 18104 30132 18110 30184
rect 18233 30175 18291 30181
rect 18233 30141 18245 30175
rect 18279 30172 18291 30175
rect 19518 30172 19524 30184
rect 18279 30144 19524 30172
rect 18279 30141 18291 30144
rect 18233 30135 18291 30141
rect 19518 30132 19524 30144
rect 19576 30132 19582 30184
rect 23750 30132 23756 30184
rect 23808 30172 23814 30184
rect 25133 30175 25191 30181
rect 25133 30172 25145 30175
rect 23808 30144 25145 30172
rect 23808 30132 23814 30144
rect 25133 30141 25145 30144
rect 25179 30141 25191 30175
rect 25133 30135 25191 30141
rect 15838 30064 15844 30116
rect 15896 30104 15902 30116
rect 17678 30104 17684 30116
rect 15896 30076 17684 30104
rect 15896 30064 15902 30076
rect 17678 30064 17684 30076
rect 17736 30064 17742 30116
rect 17954 30064 17960 30116
rect 18012 30104 18018 30116
rect 18690 30104 18696 30116
rect 18012 30076 18696 30104
rect 18012 30064 18018 30076
rect 18690 30064 18696 30076
rect 18748 30104 18754 30116
rect 21634 30104 21640 30116
rect 18748 30076 21640 30104
rect 18748 30064 18754 30076
rect 21634 30064 21640 30076
rect 21692 30064 21698 30116
rect 12253 30039 12311 30045
rect 12253 30036 12265 30039
rect 11940 30008 12265 30036
rect 11940 29996 11946 30008
rect 12253 30005 12265 30008
rect 12299 30005 12311 30039
rect 12253 29999 12311 30005
rect 12342 29996 12348 30048
rect 12400 30036 12406 30048
rect 12529 30039 12587 30045
rect 12529 30036 12541 30039
rect 12400 30008 12541 30036
rect 12400 29996 12406 30008
rect 12529 30005 12541 30008
rect 12575 30036 12587 30039
rect 14458 30036 14464 30048
rect 12575 30008 14464 30036
rect 12575 30005 12587 30008
rect 12529 29999 12587 30005
rect 14458 29996 14464 30008
rect 14516 29996 14522 30048
rect 14724 30039 14782 30045
rect 14724 30005 14736 30039
rect 14770 30036 14782 30039
rect 17494 30036 17500 30048
rect 14770 30008 17500 30036
rect 14770 30005 14782 30008
rect 14724 29999 14782 30005
rect 17494 29996 17500 30008
rect 17552 29996 17558 30048
rect 17586 29996 17592 30048
rect 17644 29996 17650 30048
rect 19429 30039 19487 30045
rect 19429 30005 19441 30039
rect 19475 30036 19487 30039
rect 21726 30036 21732 30048
rect 19475 30008 21732 30036
rect 19475 30005 19487 30008
rect 19429 29999 19487 30005
rect 21726 29996 21732 30008
rect 21784 29996 21790 30048
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 4246 29792 4252 29844
rect 4304 29832 4310 29844
rect 7285 29835 7343 29841
rect 7285 29832 7297 29835
rect 4304 29804 7297 29832
rect 4304 29792 4310 29804
rect 7285 29801 7297 29804
rect 7331 29832 7343 29835
rect 7650 29832 7656 29844
rect 7331 29804 7656 29832
rect 7331 29801 7343 29804
rect 7285 29795 7343 29801
rect 7650 29792 7656 29804
rect 7708 29792 7714 29844
rect 7742 29792 7748 29844
rect 7800 29832 7806 29844
rect 7837 29835 7895 29841
rect 7837 29832 7849 29835
rect 7800 29804 7849 29832
rect 7800 29792 7806 29804
rect 7837 29801 7849 29804
rect 7883 29801 7895 29835
rect 7837 29795 7895 29801
rect 9490 29792 9496 29844
rect 9548 29792 9554 29844
rect 14458 29792 14464 29844
rect 14516 29832 14522 29844
rect 14516 29804 14688 29832
rect 14516 29792 14522 29804
rect 11330 29724 11336 29776
rect 11388 29764 11394 29776
rect 12621 29767 12679 29773
rect 11388 29736 12434 29764
rect 11388 29724 11394 29736
rect 2682 29656 2688 29708
rect 2740 29696 2746 29708
rect 4341 29699 4399 29705
rect 4341 29696 4353 29699
rect 2740 29668 4353 29696
rect 2740 29656 2746 29668
rect 4341 29665 4353 29668
rect 4387 29665 4399 29699
rect 4341 29659 4399 29665
rect 7190 29656 7196 29708
rect 7248 29696 7254 29708
rect 8389 29699 8447 29705
rect 8389 29696 8401 29699
rect 7248 29668 8401 29696
rect 7248 29656 7254 29668
rect 8389 29665 8401 29668
rect 8435 29665 8447 29699
rect 8389 29659 8447 29665
rect 9122 29656 9128 29708
rect 9180 29696 9186 29708
rect 9217 29699 9275 29705
rect 9217 29696 9229 29699
rect 9180 29668 9229 29696
rect 9180 29656 9186 29668
rect 9217 29665 9229 29668
rect 9263 29696 9275 29699
rect 10045 29699 10103 29705
rect 10045 29696 10057 29699
rect 9263 29668 10057 29696
rect 9263 29665 9275 29668
rect 9217 29659 9275 29665
rect 10045 29665 10057 29668
rect 10091 29665 10103 29699
rect 11977 29699 12035 29705
rect 11977 29696 11989 29699
rect 10045 29659 10103 29665
rect 10152 29668 11989 29696
rect 7282 29588 7288 29640
rect 7340 29588 7346 29640
rect 7834 29588 7840 29640
rect 7892 29628 7898 29640
rect 10152 29628 10180 29668
rect 11977 29665 11989 29668
rect 12023 29665 12035 29699
rect 12406 29696 12434 29736
rect 12621 29733 12633 29767
rect 12667 29764 12679 29767
rect 14550 29764 14556 29776
rect 12667 29736 14556 29764
rect 12667 29733 12679 29736
rect 12621 29727 12679 29733
rect 14550 29724 14556 29736
rect 14608 29724 14614 29776
rect 14660 29764 14688 29804
rect 16022 29792 16028 29844
rect 16080 29832 16086 29844
rect 16482 29832 16488 29844
rect 16080 29804 16488 29832
rect 16080 29792 16086 29804
rect 16482 29792 16488 29804
rect 16540 29792 16546 29844
rect 16574 29792 16580 29844
rect 16632 29832 16638 29844
rect 18966 29832 18972 29844
rect 16632 29804 18972 29832
rect 16632 29792 16638 29804
rect 18966 29792 18972 29804
rect 19024 29792 19030 29844
rect 19794 29792 19800 29844
rect 19852 29832 19858 29844
rect 21545 29835 21603 29841
rect 19852 29804 21312 29832
rect 19852 29792 19858 29804
rect 16758 29764 16764 29776
rect 14660 29736 16764 29764
rect 16758 29724 16764 29736
rect 16816 29724 16822 29776
rect 17586 29724 17592 29776
rect 17644 29764 17650 29776
rect 17644 29736 20116 29764
rect 17644 29724 17650 29736
rect 13173 29699 13231 29705
rect 13173 29696 13185 29699
rect 12406 29668 13185 29696
rect 11977 29659 12035 29665
rect 13173 29665 13185 29668
rect 13219 29665 13231 29699
rect 13173 29659 13231 29665
rect 14458 29656 14464 29708
rect 14516 29696 14522 29708
rect 17497 29699 17555 29705
rect 17497 29696 17509 29699
rect 14516 29668 17509 29696
rect 14516 29656 14522 29668
rect 17497 29665 17509 29668
rect 17543 29665 17555 29699
rect 17497 29659 17555 29665
rect 18785 29699 18843 29705
rect 18785 29665 18797 29699
rect 18831 29696 18843 29699
rect 19058 29696 19064 29708
rect 18831 29668 19064 29696
rect 18831 29665 18843 29668
rect 18785 29659 18843 29665
rect 19058 29656 19064 29668
rect 19116 29656 19122 29708
rect 20088 29705 20116 29736
rect 20073 29699 20131 29705
rect 20073 29665 20085 29699
rect 20119 29665 20131 29699
rect 20073 29659 20131 29665
rect 20257 29699 20315 29705
rect 20257 29665 20269 29699
rect 20303 29696 20315 29699
rect 21174 29696 21180 29708
rect 20303 29668 21180 29696
rect 20303 29665 20315 29668
rect 20257 29659 20315 29665
rect 21174 29656 21180 29668
rect 21232 29656 21238 29708
rect 21284 29696 21312 29804
rect 21545 29801 21557 29835
rect 21591 29832 21603 29835
rect 25682 29832 25688 29844
rect 21591 29804 25688 29832
rect 21591 29801 21603 29804
rect 21545 29795 21603 29801
rect 25682 29792 25688 29804
rect 25740 29792 25746 29844
rect 21634 29724 21640 29776
rect 21692 29764 21698 29776
rect 22830 29764 22836 29776
rect 21692 29736 22836 29764
rect 21692 29724 21698 29736
rect 22830 29724 22836 29736
rect 22888 29724 22894 29776
rect 22925 29767 22983 29773
rect 22925 29733 22937 29767
rect 22971 29764 22983 29767
rect 24762 29764 24768 29776
rect 22971 29736 24768 29764
rect 22971 29733 22983 29736
rect 22925 29727 22983 29733
rect 24762 29724 24768 29736
rect 24820 29724 24826 29776
rect 22189 29699 22247 29705
rect 21284 29668 22140 29696
rect 7892 29600 10180 29628
rect 7892 29588 7898 29600
rect 10410 29588 10416 29640
rect 10468 29628 10474 29640
rect 12989 29631 13047 29637
rect 12989 29628 13001 29631
rect 10468 29600 13001 29628
rect 10468 29588 10474 29600
rect 12989 29597 13001 29600
rect 13035 29597 13047 29631
rect 12989 29591 13047 29597
rect 13998 29588 14004 29640
rect 14056 29628 14062 29640
rect 15286 29628 15292 29640
rect 14056 29600 15292 29628
rect 14056 29588 14062 29600
rect 15286 29588 15292 29600
rect 15344 29588 15350 29640
rect 16298 29588 16304 29640
rect 16356 29628 16362 29640
rect 17405 29631 17463 29637
rect 17405 29628 17417 29631
rect 16356 29600 17417 29628
rect 16356 29588 16362 29600
rect 17405 29597 17417 29600
rect 17451 29597 17463 29631
rect 17405 29591 17463 29597
rect 18046 29588 18052 29640
rect 18104 29628 18110 29640
rect 18966 29628 18972 29640
rect 18104 29600 18972 29628
rect 18104 29588 18110 29600
rect 18966 29588 18972 29600
rect 19024 29588 19030 29640
rect 19981 29631 20039 29637
rect 19981 29597 19993 29631
rect 20027 29628 20039 29631
rect 20806 29628 20812 29640
rect 20027 29600 20812 29628
rect 20027 29597 20039 29600
rect 19981 29591 20039 29597
rect 20806 29588 20812 29600
rect 20864 29588 20870 29640
rect 21913 29631 21971 29637
rect 21913 29597 21925 29631
rect 21959 29628 21971 29631
rect 22002 29628 22008 29640
rect 21959 29600 22008 29628
rect 21959 29597 21971 29600
rect 21913 29591 21971 29597
rect 22002 29588 22008 29600
rect 22060 29588 22066 29640
rect 22112 29628 22140 29668
rect 22189 29665 22201 29699
rect 22235 29696 22247 29699
rect 22554 29696 22560 29708
rect 22235 29668 22560 29696
rect 22235 29665 22247 29668
rect 22189 29659 22247 29665
rect 22554 29656 22560 29668
rect 22612 29656 22618 29708
rect 23382 29656 23388 29708
rect 23440 29656 23446 29708
rect 23569 29699 23627 29705
rect 23569 29665 23581 29699
rect 23615 29696 23627 29699
rect 23750 29696 23756 29708
rect 23615 29668 23756 29696
rect 23615 29665 23627 29668
rect 23569 29659 23627 29665
rect 23750 29656 23756 29668
rect 23808 29656 23814 29708
rect 22278 29628 22284 29640
rect 22112 29600 22284 29628
rect 22278 29588 22284 29600
rect 22336 29588 22342 29640
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 3418 29520 3424 29572
rect 3476 29560 3482 29572
rect 4433 29563 4491 29569
rect 4433 29560 4445 29563
rect 3476 29532 4445 29560
rect 3476 29520 3482 29532
rect 4433 29529 4445 29532
rect 4479 29529 4491 29563
rect 4433 29523 4491 29529
rect 5258 29520 5264 29572
rect 5316 29560 5322 29572
rect 5353 29563 5411 29569
rect 5353 29560 5365 29563
rect 5316 29532 5365 29560
rect 5316 29520 5322 29532
rect 5353 29529 5365 29532
rect 5399 29529 5411 29563
rect 5353 29523 5411 29529
rect 7006 29520 7012 29572
rect 7064 29560 7070 29572
rect 7300 29560 7328 29588
rect 7469 29563 7527 29569
rect 7469 29560 7481 29563
rect 7064 29532 7481 29560
rect 7064 29520 7070 29532
rect 7469 29529 7481 29532
rect 7515 29560 7527 29563
rect 8297 29563 8355 29569
rect 8297 29560 8309 29563
rect 7515 29532 8309 29560
rect 7515 29529 7527 29532
rect 7469 29523 7527 29529
rect 8297 29529 8309 29532
rect 8343 29529 8355 29563
rect 8297 29523 8355 29529
rect 9306 29520 9312 29572
rect 9364 29560 9370 29572
rect 9582 29560 9588 29572
rect 9364 29532 9588 29560
rect 9364 29520 9370 29532
rect 9582 29520 9588 29532
rect 9640 29560 9646 29572
rect 9861 29563 9919 29569
rect 9861 29560 9873 29563
rect 9640 29532 9873 29560
rect 9640 29520 9646 29532
rect 9861 29529 9873 29532
rect 9907 29529 9919 29563
rect 9861 29523 9919 29529
rect 11793 29563 11851 29569
rect 11793 29529 11805 29563
rect 11839 29560 11851 29563
rect 12342 29560 12348 29572
rect 11839 29532 12348 29560
rect 11839 29529 11851 29532
rect 11793 29523 11851 29529
rect 12342 29520 12348 29532
rect 12400 29520 12406 29572
rect 12802 29520 12808 29572
rect 12860 29560 12866 29572
rect 13081 29563 13139 29569
rect 13081 29560 13093 29563
rect 12860 29532 13093 29560
rect 12860 29520 12866 29532
rect 13081 29529 13093 29532
rect 13127 29529 13139 29563
rect 13081 29523 13139 29529
rect 14734 29520 14740 29572
rect 14792 29520 14798 29572
rect 16574 29560 16580 29572
rect 15028 29532 16580 29560
rect 7650 29452 7656 29504
rect 7708 29492 7714 29504
rect 8205 29495 8263 29501
rect 8205 29492 8217 29495
rect 7708 29464 8217 29492
rect 7708 29452 7714 29464
rect 8205 29461 8217 29464
rect 8251 29461 8263 29495
rect 8205 29455 8263 29461
rect 9033 29495 9091 29501
rect 9033 29461 9045 29495
rect 9079 29492 9091 29495
rect 9953 29495 10011 29501
rect 9953 29492 9965 29495
rect 9079 29464 9965 29492
rect 9079 29461 9091 29464
rect 9033 29455 9091 29461
rect 9953 29461 9965 29464
rect 9999 29492 10011 29495
rect 10042 29492 10048 29504
rect 9999 29464 10048 29492
rect 9999 29461 10011 29464
rect 9953 29455 10011 29461
rect 10042 29452 10048 29464
rect 10100 29452 10106 29504
rect 10778 29452 10784 29504
rect 10836 29492 10842 29504
rect 11425 29495 11483 29501
rect 11425 29492 11437 29495
rect 10836 29464 11437 29492
rect 10836 29452 10842 29464
rect 11425 29461 11437 29464
rect 11471 29461 11483 29495
rect 11425 29455 11483 29461
rect 11882 29452 11888 29504
rect 11940 29452 11946 29504
rect 12894 29452 12900 29504
rect 12952 29492 12958 29504
rect 13725 29495 13783 29501
rect 13725 29492 13737 29495
rect 12952 29464 13737 29492
rect 12952 29452 12958 29464
rect 13725 29461 13737 29464
rect 13771 29492 13783 29495
rect 15028 29492 15056 29532
rect 16574 29520 16580 29532
rect 16632 29520 16638 29572
rect 17313 29563 17371 29569
rect 17313 29529 17325 29563
rect 17359 29560 17371 29563
rect 17586 29560 17592 29572
rect 17359 29532 17592 29560
rect 17359 29529 17371 29532
rect 17313 29523 17371 29529
rect 17586 29520 17592 29532
rect 17644 29520 17650 29572
rect 18601 29563 18659 29569
rect 18601 29529 18613 29563
rect 18647 29560 18659 29563
rect 19334 29560 19340 29572
rect 18647 29532 19340 29560
rect 18647 29529 18659 29532
rect 18601 29523 18659 29529
rect 19334 29520 19340 29532
rect 19392 29560 19398 29572
rect 19392 29532 25176 29560
rect 19392 29520 19398 29532
rect 13771 29464 15056 29492
rect 13771 29461 13783 29464
rect 13725 29455 13783 29461
rect 15102 29452 15108 29504
rect 15160 29492 15166 29504
rect 16945 29495 17003 29501
rect 16945 29492 16957 29495
rect 15160 29464 16957 29492
rect 15160 29452 15166 29464
rect 16945 29461 16957 29464
rect 16991 29461 17003 29495
rect 16945 29455 17003 29461
rect 17494 29452 17500 29504
rect 17552 29492 17558 29504
rect 18141 29495 18199 29501
rect 18141 29492 18153 29495
rect 17552 29464 18153 29492
rect 17552 29452 17558 29464
rect 18141 29461 18153 29464
rect 18187 29461 18199 29495
rect 18141 29455 18199 29461
rect 18230 29452 18236 29504
rect 18288 29492 18294 29504
rect 18414 29492 18420 29504
rect 18288 29464 18420 29492
rect 18288 29452 18294 29464
rect 18414 29452 18420 29464
rect 18472 29452 18478 29504
rect 18506 29452 18512 29504
rect 18564 29452 18570 29504
rect 19613 29495 19671 29501
rect 19613 29461 19625 29495
rect 19659 29492 19671 29495
rect 20346 29492 20352 29504
rect 19659 29464 20352 29492
rect 19659 29461 19671 29464
rect 19613 29455 19671 29461
rect 20346 29452 20352 29464
rect 20404 29452 20410 29504
rect 20898 29452 20904 29504
rect 20956 29452 20962 29504
rect 21450 29452 21456 29504
rect 21508 29492 21514 29504
rect 22005 29495 22063 29501
rect 22005 29492 22017 29495
rect 21508 29464 22017 29492
rect 21508 29452 21514 29464
rect 22005 29461 22017 29464
rect 22051 29461 22063 29495
rect 22005 29455 22063 29461
rect 23290 29452 23296 29504
rect 23348 29452 23354 29504
rect 25148 29501 25176 29532
rect 25133 29495 25191 29501
rect 25133 29461 25145 29495
rect 25179 29461 25191 29495
rect 25133 29455 25191 29461
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 7742 29248 7748 29300
rect 7800 29288 7806 29300
rect 7800 29260 12434 29288
rect 7800 29248 7806 29260
rect 9490 29220 9496 29232
rect 9246 29192 9496 29220
rect 9490 29180 9496 29192
rect 9548 29220 9554 29232
rect 9769 29223 9827 29229
rect 9769 29220 9781 29223
rect 9548 29192 9781 29220
rect 9548 29180 9554 29192
rect 9769 29189 9781 29192
rect 9815 29189 9827 29223
rect 12406 29220 12434 29260
rect 12894 29248 12900 29300
rect 12952 29248 12958 29300
rect 14185 29291 14243 29297
rect 14185 29257 14197 29291
rect 14231 29288 14243 29291
rect 15562 29288 15568 29300
rect 14231 29260 15568 29288
rect 14231 29257 14243 29260
rect 14185 29251 14243 29257
rect 15562 29248 15568 29260
rect 15620 29248 15626 29300
rect 16025 29291 16083 29297
rect 16025 29257 16037 29291
rect 16071 29288 16083 29291
rect 16390 29288 16396 29300
rect 16071 29260 16396 29288
rect 16071 29257 16083 29260
rect 16025 29251 16083 29257
rect 12406 29192 15516 29220
rect 9769 29183 9827 29189
rect 12989 29155 13047 29161
rect 9508 29124 12756 29152
rect 6546 29044 6552 29096
rect 6604 29084 6610 29096
rect 7745 29087 7803 29093
rect 7745 29084 7757 29087
rect 6604 29056 7757 29084
rect 6604 29044 6610 29056
rect 7745 29053 7757 29056
rect 7791 29053 7803 29087
rect 7745 29047 7803 29053
rect 9398 29044 9404 29096
rect 9456 29084 9462 29096
rect 9508 29093 9536 29124
rect 9493 29087 9551 29093
rect 9493 29084 9505 29087
rect 9456 29056 9505 29084
rect 9456 29044 9462 29056
rect 9493 29053 9505 29056
rect 9539 29053 9551 29087
rect 9493 29047 9551 29053
rect 10870 28976 10876 29028
rect 10928 29016 10934 29028
rect 12529 29019 12587 29025
rect 12529 29016 12541 29019
rect 10928 28988 12541 29016
rect 10928 28976 10934 28988
rect 12529 28985 12541 28988
rect 12575 28985 12587 29019
rect 12728 29016 12756 29124
rect 12989 29121 13001 29155
rect 13035 29152 13047 29155
rect 13998 29152 14004 29164
rect 13035 29124 14004 29152
rect 13035 29121 13047 29124
rect 12989 29115 13047 29121
rect 13998 29112 14004 29124
rect 14056 29112 14062 29164
rect 14090 29112 14096 29164
rect 14148 29112 14154 29164
rect 15289 29155 15347 29161
rect 15289 29121 15301 29155
rect 15335 29121 15347 29155
rect 15289 29115 15347 29121
rect 13081 29087 13139 29093
rect 13081 29053 13093 29087
rect 13127 29053 13139 29087
rect 13081 29047 13139 29053
rect 13096 29016 13124 29047
rect 13538 29044 13544 29096
rect 13596 29084 13602 29096
rect 14369 29087 14427 29093
rect 13596 29056 13860 29084
rect 13596 29044 13602 29056
rect 12728 28988 13124 29016
rect 12529 28979 12587 28985
rect 13630 28976 13636 29028
rect 13688 29016 13694 29028
rect 13725 29019 13783 29025
rect 13725 29016 13737 29019
rect 13688 28988 13737 29016
rect 13688 28976 13694 28988
rect 13725 28985 13737 28988
rect 13771 28985 13783 29019
rect 13832 29016 13860 29056
rect 14369 29053 14381 29087
rect 14415 29084 14427 29087
rect 14642 29084 14648 29096
rect 14415 29056 14648 29084
rect 14415 29053 14427 29056
rect 14369 29047 14427 29053
rect 14642 29044 14648 29056
rect 14700 29044 14706 29096
rect 14921 29019 14979 29025
rect 14921 29016 14933 29019
rect 13832 28988 14933 29016
rect 13725 28979 13783 28985
rect 14921 28985 14933 28988
rect 14967 28985 14979 29019
rect 15304 29016 15332 29115
rect 15378 29044 15384 29096
rect 15436 29044 15442 29096
rect 15488 29093 15516 29192
rect 15473 29087 15531 29093
rect 15473 29053 15485 29087
rect 15519 29053 15531 29087
rect 15473 29047 15531 29053
rect 16040 29016 16068 29251
rect 16390 29248 16396 29260
rect 16448 29248 16454 29300
rect 17218 29248 17224 29300
rect 17276 29248 17282 29300
rect 17313 29291 17371 29297
rect 17313 29257 17325 29291
rect 17359 29288 17371 29291
rect 17494 29288 17500 29300
rect 17359 29260 17500 29288
rect 17359 29257 17371 29260
rect 17313 29251 17371 29257
rect 17494 29248 17500 29260
rect 17552 29248 17558 29300
rect 17586 29248 17592 29300
rect 17644 29288 17650 29300
rect 17957 29291 18015 29297
rect 17957 29288 17969 29291
rect 17644 29260 17969 29288
rect 17644 29248 17650 29260
rect 17957 29257 17969 29260
rect 18003 29288 18015 29291
rect 19794 29288 19800 29300
rect 18003 29260 19800 29288
rect 18003 29257 18015 29260
rect 17957 29251 18015 29257
rect 19794 29248 19800 29260
rect 19852 29248 19858 29300
rect 20162 29248 20168 29300
rect 20220 29288 20226 29300
rect 20220 29260 20852 29288
rect 20220 29248 20226 29260
rect 16209 29223 16267 29229
rect 16209 29189 16221 29223
rect 16255 29220 16267 29223
rect 18874 29220 18880 29232
rect 16255 29192 18880 29220
rect 16255 29189 16267 29192
rect 16209 29183 16267 29189
rect 15304 28988 16068 29016
rect 14921 28979 14979 28985
rect 8008 28951 8066 28957
rect 8008 28917 8020 28951
rect 8054 28948 8066 28951
rect 9674 28948 9680 28960
rect 8054 28920 9680 28948
rect 8054 28917 8066 28920
rect 8008 28911 8066 28917
rect 9674 28908 9680 28920
rect 9732 28908 9738 28960
rect 15194 28908 15200 28960
rect 15252 28948 15258 28960
rect 16022 28948 16028 28960
rect 15252 28920 16028 28948
rect 15252 28908 15258 28920
rect 16022 28908 16028 28920
rect 16080 28948 16086 28960
rect 16224 28948 16252 29183
rect 18874 29180 18880 29192
rect 18932 29180 18938 29232
rect 20070 29220 20076 29232
rect 18984 29192 20076 29220
rect 16758 29112 16764 29164
rect 16816 29152 16822 29164
rect 18984 29152 19012 29192
rect 20070 29180 20076 29192
rect 20128 29180 20134 29232
rect 20530 29180 20536 29232
rect 20588 29180 20594 29232
rect 20824 29220 20852 29260
rect 20898 29248 20904 29300
rect 20956 29288 20962 29300
rect 22373 29291 22431 29297
rect 22373 29288 22385 29291
rect 20956 29260 22385 29288
rect 20956 29248 20962 29260
rect 22373 29257 22385 29260
rect 22419 29257 22431 29291
rect 22373 29251 22431 29257
rect 22830 29248 22836 29300
rect 22888 29288 22894 29300
rect 23937 29291 23995 29297
rect 23937 29288 23949 29291
rect 22888 29260 23949 29288
rect 22888 29248 22894 29260
rect 23937 29257 23949 29260
rect 23983 29257 23995 29291
rect 23937 29251 23995 29257
rect 25314 29248 25320 29300
rect 25372 29248 25378 29300
rect 25498 29248 25504 29300
rect 25556 29248 25562 29300
rect 21085 29223 21143 29229
rect 21085 29220 21097 29223
rect 20824 29192 21097 29220
rect 21085 29189 21097 29192
rect 21131 29189 21143 29223
rect 21085 29183 21143 29189
rect 20441 29155 20499 29161
rect 20441 29152 20453 29155
rect 16816 29124 19012 29152
rect 19720 29124 20453 29152
rect 16816 29112 16822 29124
rect 17402 29044 17408 29096
rect 17460 29044 17466 29096
rect 19720 29093 19748 29124
rect 20441 29121 20453 29124
rect 20487 29121 20499 29155
rect 20548 29152 20576 29180
rect 21100 29152 21128 29183
rect 21542 29180 21548 29232
rect 21600 29220 21606 29232
rect 22465 29223 22523 29229
rect 22465 29220 22477 29223
rect 21600 29192 22477 29220
rect 21600 29180 21606 29192
rect 22465 29189 22477 29192
rect 22511 29189 22523 29223
rect 22465 29183 22523 29189
rect 24578 29180 24584 29232
rect 24636 29220 24642 29232
rect 24673 29223 24731 29229
rect 24673 29220 24685 29223
rect 24636 29192 24685 29220
rect 24636 29180 24642 29192
rect 24673 29189 24685 29192
rect 24719 29189 24731 29223
rect 24673 29183 24731 29189
rect 22738 29152 22744 29164
rect 20548 29124 20668 29152
rect 21100 29124 22744 29152
rect 20441 29115 20499 29121
rect 19705 29087 19763 29093
rect 19705 29084 19717 29087
rect 17696 29056 19717 29084
rect 16390 28976 16396 29028
rect 16448 29016 16454 29028
rect 17696 29016 17724 29056
rect 19705 29053 19717 29056
rect 19751 29053 19763 29087
rect 19705 29047 19763 29053
rect 20162 29044 20168 29096
rect 20220 29084 20226 29096
rect 20640 29093 20668 29124
rect 22738 29112 22744 29124
rect 22796 29112 22802 29164
rect 23661 29155 23719 29161
rect 23661 29121 23673 29155
rect 23707 29152 23719 29155
rect 24118 29152 24124 29164
rect 23707 29124 24124 29152
rect 23707 29121 23719 29124
rect 23661 29115 23719 29121
rect 24118 29112 24124 29124
rect 24176 29112 24182 29164
rect 20533 29087 20591 29093
rect 20533 29084 20545 29087
rect 20220 29056 20545 29084
rect 20220 29044 20226 29056
rect 20533 29053 20545 29056
rect 20579 29053 20591 29087
rect 20533 29047 20591 29053
rect 20625 29087 20683 29093
rect 20625 29053 20637 29087
rect 20671 29053 20683 29087
rect 22462 29084 22468 29096
rect 20625 29047 20683 29053
rect 21100 29056 22468 29084
rect 16448 28988 17724 29016
rect 18141 29019 18199 29025
rect 16448 28976 16454 28988
rect 18141 28985 18153 29019
rect 18187 29016 18199 29019
rect 18506 29016 18512 29028
rect 18187 28988 18512 29016
rect 18187 28985 18199 28988
rect 18141 28979 18199 28985
rect 18506 28976 18512 28988
rect 18564 28976 18570 29028
rect 20073 29019 20131 29025
rect 20073 28985 20085 29019
rect 20119 29016 20131 29019
rect 21100 29016 21128 29056
rect 22462 29044 22468 29056
rect 22520 29044 22526 29096
rect 22649 29087 22707 29093
rect 22649 29053 22661 29087
rect 22695 29084 22707 29087
rect 23566 29084 23572 29096
rect 22695 29056 23572 29084
rect 22695 29053 22707 29056
rect 22649 29047 22707 29053
rect 23566 29044 23572 29056
rect 23624 29044 23630 29096
rect 20119 28988 21128 29016
rect 22005 29019 22063 29025
rect 20119 28985 20131 28988
rect 20073 28979 20131 28985
rect 22005 28985 22017 29019
rect 22051 29016 22063 29019
rect 23290 29016 23296 29028
rect 22051 28988 23296 29016
rect 22051 28985 22063 28988
rect 22005 28979 22063 28985
rect 23290 28976 23296 28988
rect 23348 28976 23354 29028
rect 23382 28976 23388 29028
rect 23440 29016 23446 29028
rect 24857 29019 24915 29025
rect 24857 29016 24869 29019
rect 23440 28988 24869 29016
rect 23440 28976 23446 28988
rect 24857 28985 24869 28988
rect 24903 28985 24915 29019
rect 24857 28979 24915 28985
rect 16080 28920 16252 28948
rect 16080 28908 16086 28920
rect 16850 28908 16856 28960
rect 16908 28908 16914 28960
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 8110 28704 8116 28756
rect 8168 28744 8174 28756
rect 8665 28747 8723 28753
rect 8665 28744 8677 28747
rect 8168 28716 8677 28744
rect 8168 28704 8174 28716
rect 8665 28713 8677 28716
rect 8711 28744 8723 28747
rect 9490 28744 9496 28756
rect 8711 28716 9496 28744
rect 8711 28713 8723 28716
rect 8665 28707 8723 28713
rect 9490 28704 9496 28716
rect 9548 28704 9554 28756
rect 12805 28747 12863 28753
rect 12805 28713 12817 28747
rect 12851 28744 12863 28747
rect 14090 28744 14096 28756
rect 12851 28716 14096 28744
rect 12851 28713 12863 28716
rect 12805 28707 12863 28713
rect 14090 28704 14096 28716
rect 14148 28704 14154 28756
rect 18782 28704 18788 28756
rect 18840 28744 18846 28756
rect 18966 28744 18972 28756
rect 18840 28716 18972 28744
rect 18840 28704 18846 28716
rect 18966 28704 18972 28716
rect 19024 28744 19030 28756
rect 19024 28716 20760 28744
rect 19024 28704 19030 28716
rect 8297 28679 8355 28685
rect 8297 28645 8309 28679
rect 8343 28676 8355 28679
rect 9858 28676 9864 28688
rect 8343 28648 9864 28676
rect 8343 28645 8355 28648
rect 8297 28639 8355 28645
rect 9858 28636 9864 28648
rect 9916 28636 9922 28688
rect 16390 28636 16396 28688
rect 16448 28676 16454 28688
rect 18322 28676 18328 28688
rect 16448 28648 18328 28676
rect 16448 28636 16454 28648
rect 18322 28636 18328 28648
rect 18380 28636 18386 28688
rect 20732 28676 20760 28716
rect 21174 28704 21180 28756
rect 21232 28704 21238 28756
rect 23845 28679 23903 28685
rect 23845 28676 23857 28679
rect 20732 28648 23857 28676
rect 23845 28645 23857 28648
rect 23891 28645 23903 28679
rect 23845 28639 23903 28645
rect 1302 28568 1308 28620
rect 1360 28608 1366 28620
rect 2041 28611 2099 28617
rect 2041 28608 2053 28611
rect 1360 28580 2053 28608
rect 1360 28568 1366 28580
rect 2041 28577 2053 28580
rect 2087 28577 2099 28611
rect 2041 28571 2099 28577
rect 4062 28568 4068 28620
rect 4120 28608 4126 28620
rect 4341 28611 4399 28617
rect 4341 28608 4353 28611
rect 4120 28580 4353 28608
rect 4120 28568 4126 28580
rect 4341 28577 4353 28580
rect 4387 28577 4399 28611
rect 4341 28571 4399 28577
rect 5166 28568 5172 28620
rect 5224 28568 5230 28620
rect 6546 28568 6552 28620
rect 6604 28568 6610 28620
rect 6825 28611 6883 28617
rect 6825 28577 6837 28611
rect 6871 28608 6883 28611
rect 9398 28608 9404 28620
rect 6871 28580 9404 28608
rect 6871 28577 6883 28580
rect 6825 28571 6883 28577
rect 9398 28568 9404 28580
rect 9456 28568 9462 28620
rect 10873 28611 10931 28617
rect 10873 28577 10885 28611
rect 10919 28608 10931 28611
rect 11330 28608 11336 28620
rect 10919 28580 11336 28608
rect 10919 28577 10931 28580
rect 10873 28571 10931 28577
rect 11330 28568 11336 28580
rect 11388 28568 11394 28620
rect 13354 28568 13360 28620
rect 13412 28568 13418 28620
rect 14826 28568 14832 28620
rect 14884 28568 14890 28620
rect 16206 28568 16212 28620
rect 16264 28568 16270 28620
rect 17126 28568 17132 28620
rect 17184 28608 17190 28620
rect 17681 28611 17739 28617
rect 17681 28608 17693 28611
rect 17184 28580 17693 28608
rect 17184 28568 17190 28580
rect 17681 28577 17693 28580
rect 17727 28577 17739 28611
rect 17681 28571 17739 28577
rect 17770 28568 17776 28620
rect 17828 28568 17834 28620
rect 19429 28611 19487 28617
rect 19429 28577 19441 28611
rect 19475 28608 19487 28611
rect 22002 28608 22008 28620
rect 19475 28580 22008 28608
rect 19475 28577 19487 28580
rect 19429 28571 19487 28577
rect 22002 28568 22008 28580
rect 22060 28568 22066 28620
rect 1762 28500 1768 28552
rect 1820 28500 1826 28552
rect 9950 28500 9956 28552
rect 10008 28540 10014 28552
rect 10597 28543 10655 28549
rect 10597 28540 10609 28543
rect 10008 28512 10609 28540
rect 10008 28500 10014 28512
rect 10597 28509 10609 28512
rect 10643 28509 10655 28543
rect 10597 28503 10655 28509
rect 14645 28543 14703 28549
rect 14645 28509 14657 28543
rect 14691 28540 14703 28543
rect 15194 28540 15200 28552
rect 14691 28512 15200 28540
rect 14691 28509 14703 28512
rect 14645 28503 14703 28509
rect 15194 28500 15200 28512
rect 15252 28500 15258 28552
rect 16025 28543 16083 28549
rect 16025 28509 16037 28543
rect 16071 28540 16083 28543
rect 16850 28540 16856 28552
rect 16071 28512 16856 28540
rect 16071 28509 16083 28512
rect 16025 28503 16083 28509
rect 16850 28500 16856 28512
rect 16908 28500 16914 28552
rect 17589 28543 17647 28549
rect 17589 28509 17601 28543
rect 17635 28540 17647 28543
rect 17862 28540 17868 28552
rect 17635 28512 17868 28540
rect 17635 28509 17647 28512
rect 17589 28503 17647 28509
rect 17862 28500 17868 28512
rect 17920 28500 17926 28552
rect 24029 28543 24087 28549
rect 24029 28509 24041 28543
rect 24075 28509 24087 28543
rect 24029 28503 24087 28509
rect 4433 28475 4491 28481
rect 4433 28441 4445 28475
rect 4479 28441 4491 28475
rect 8110 28472 8116 28484
rect 8050 28444 8116 28472
rect 4433 28435 4491 28441
rect 3970 28364 3976 28416
rect 4028 28404 4034 28416
rect 4448 28404 4476 28435
rect 8110 28432 8116 28444
rect 8168 28432 8174 28484
rect 12526 28472 12532 28484
rect 12098 28444 12532 28472
rect 12526 28432 12532 28444
rect 12584 28472 12590 28484
rect 13354 28472 13360 28484
rect 12584 28444 13360 28472
rect 12584 28432 12590 28444
rect 13354 28432 13360 28444
rect 13412 28472 13418 28484
rect 15470 28472 15476 28484
rect 13412 28444 15476 28472
rect 13412 28432 13418 28444
rect 15470 28432 15476 28444
rect 15528 28432 15534 28484
rect 16117 28475 16175 28481
rect 16117 28441 16129 28475
rect 16163 28472 16175 28475
rect 16666 28472 16672 28484
rect 16163 28444 16672 28472
rect 16163 28441 16175 28444
rect 16117 28435 16175 28441
rect 16666 28432 16672 28444
rect 16724 28432 16730 28484
rect 19610 28432 19616 28484
rect 19668 28472 19674 28484
rect 19705 28475 19763 28481
rect 19705 28472 19717 28475
rect 19668 28444 19717 28472
rect 19668 28432 19674 28444
rect 19705 28441 19717 28444
rect 19751 28441 19763 28475
rect 21453 28475 21511 28481
rect 21453 28472 21465 28475
rect 20930 28444 21465 28472
rect 19705 28435 19763 28441
rect 21453 28441 21465 28444
rect 21499 28472 21511 28475
rect 22186 28472 22192 28484
rect 21499 28444 22192 28472
rect 21499 28441 21511 28444
rect 21453 28435 21511 28441
rect 22186 28432 22192 28444
rect 22244 28432 22250 28484
rect 24044 28472 24072 28503
rect 24762 28500 24768 28552
rect 24820 28500 24826 28552
rect 24210 28472 24216 28484
rect 24044 28444 24216 28472
rect 24210 28432 24216 28444
rect 24268 28472 24274 28484
rect 24854 28472 24860 28484
rect 24268 28444 24860 28472
rect 24268 28432 24274 28444
rect 24854 28432 24860 28444
rect 24912 28432 24918 28484
rect 4028 28376 4476 28404
rect 12345 28407 12403 28413
rect 4028 28364 4034 28376
rect 12345 28373 12357 28407
rect 12391 28404 12403 28407
rect 12802 28404 12808 28416
rect 12391 28376 12808 28404
rect 12391 28373 12403 28376
rect 12345 28367 12403 28373
rect 12802 28364 12808 28376
rect 12860 28364 12866 28416
rect 13170 28364 13176 28416
rect 13228 28364 13234 28416
rect 13262 28364 13268 28416
rect 13320 28364 13326 28416
rect 13909 28407 13967 28413
rect 13909 28373 13921 28407
rect 13955 28404 13967 28407
rect 13998 28404 14004 28416
rect 13955 28376 14004 28404
rect 13955 28373 13967 28376
rect 13909 28367 13967 28373
rect 13998 28364 14004 28376
rect 14056 28364 14062 28416
rect 14274 28364 14280 28416
rect 14332 28364 14338 28416
rect 14737 28407 14795 28413
rect 14737 28373 14749 28407
rect 14783 28404 14795 28407
rect 14918 28404 14924 28416
rect 14783 28376 14924 28404
rect 14783 28373 14795 28376
rect 14737 28367 14795 28373
rect 14918 28364 14924 28376
rect 14976 28364 14982 28416
rect 15286 28364 15292 28416
rect 15344 28364 15350 28416
rect 15657 28407 15715 28413
rect 15657 28373 15669 28407
rect 15703 28404 15715 28407
rect 15746 28404 15752 28416
rect 15703 28376 15752 28404
rect 15703 28373 15715 28376
rect 15657 28367 15715 28373
rect 15746 28364 15752 28376
rect 15804 28364 15810 28416
rect 16758 28364 16764 28416
rect 16816 28364 16822 28416
rect 16942 28364 16948 28416
rect 17000 28404 17006 28416
rect 17221 28407 17279 28413
rect 17221 28404 17233 28407
rect 17000 28376 17233 28404
rect 17000 28364 17006 28376
rect 17221 28373 17233 28376
rect 17267 28373 17279 28407
rect 17221 28367 17279 28373
rect 24578 28364 24584 28416
rect 24636 28364 24642 28416
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 1946 28160 1952 28212
rect 2004 28200 2010 28212
rect 3786 28209 3792 28212
rect 2041 28203 2099 28209
rect 2041 28200 2053 28203
rect 2004 28172 2053 28200
rect 2004 28160 2010 28172
rect 2041 28169 2053 28172
rect 2087 28169 2099 28203
rect 2041 28163 2099 28169
rect 3743 28203 3792 28209
rect 3743 28169 3755 28203
rect 3789 28169 3792 28203
rect 3743 28163 3792 28169
rect 3786 28160 3792 28163
rect 3844 28160 3850 28212
rect 12621 28203 12679 28209
rect 12621 28169 12633 28203
rect 12667 28200 12679 28203
rect 13170 28200 13176 28212
rect 12667 28172 13176 28200
rect 12667 28169 12679 28172
rect 12621 28163 12679 28169
rect 13170 28160 13176 28172
rect 13228 28160 13234 28212
rect 13354 28160 13360 28212
rect 13412 28160 13418 28212
rect 15470 28160 15476 28212
rect 15528 28200 15534 28212
rect 15930 28200 15936 28212
rect 15528 28172 15936 28200
rect 15528 28160 15534 28172
rect 15930 28160 15936 28172
rect 15988 28200 15994 28212
rect 16853 28203 16911 28209
rect 16853 28200 16865 28203
rect 15988 28172 16865 28200
rect 15988 28160 15994 28172
rect 16853 28169 16865 28172
rect 16899 28169 16911 28203
rect 16853 28163 16911 28169
rect 18322 28160 18328 28212
rect 18380 28160 18386 28212
rect 19058 28160 19064 28212
rect 19116 28200 19122 28212
rect 23753 28203 23811 28209
rect 23753 28200 23765 28203
rect 19116 28172 23765 28200
rect 19116 28160 19122 28172
rect 23753 28169 23765 28172
rect 23799 28169 23811 28203
rect 23753 28163 23811 28169
rect 16390 28092 16396 28144
rect 16448 28132 16454 28144
rect 16669 28135 16727 28141
rect 16669 28132 16681 28135
rect 16448 28104 16681 28132
rect 16448 28092 16454 28104
rect 16669 28101 16681 28104
rect 16715 28101 16727 28135
rect 21082 28132 21088 28144
rect 16669 28095 16727 28101
rect 17052 28104 21088 28132
rect 2225 28067 2283 28073
rect 2225 28033 2237 28067
rect 2271 28064 2283 28067
rect 3326 28064 3332 28076
rect 2271 28036 3332 28064
rect 2271 28033 2283 28036
rect 2225 28027 2283 28033
rect 3326 28024 3332 28036
rect 3384 28024 3390 28076
rect 3602 28024 3608 28076
rect 3660 28073 3666 28076
rect 3660 28067 3698 28073
rect 3686 28033 3698 28067
rect 13173 28067 13231 28073
rect 9706 28036 10732 28064
rect 3660 28027 3698 28033
rect 3660 28024 3666 28027
rect 8297 27999 8355 28005
rect 8297 27965 8309 27999
rect 8343 27996 8355 27999
rect 8343 27968 8432 27996
rect 8343 27965 8355 27968
rect 8297 27959 8355 27965
rect 8404 27860 8432 27968
rect 8570 27956 8576 28008
rect 8628 27956 8634 28008
rect 9674 27888 9680 27940
rect 9732 27928 9738 27940
rect 10045 27931 10103 27937
rect 10045 27928 10057 27931
rect 9732 27900 10057 27928
rect 9732 27888 9738 27900
rect 10045 27897 10057 27900
rect 10091 27928 10103 27931
rect 10594 27928 10600 27940
rect 10091 27900 10600 27928
rect 10091 27897 10103 27900
rect 10045 27891 10103 27897
rect 10594 27888 10600 27900
rect 10652 27888 10658 27940
rect 10704 27872 10732 28036
rect 13173 28033 13185 28067
rect 13219 28064 13231 28067
rect 13262 28064 13268 28076
rect 13219 28036 13268 28064
rect 13219 28033 13231 28036
rect 13173 28027 13231 28033
rect 13262 28024 13268 28036
rect 13320 28024 13326 28076
rect 15930 28024 15936 28076
rect 15988 28064 15994 28076
rect 16408 28064 16436 28092
rect 15988 28036 16436 28064
rect 15988 28024 15994 28036
rect 16022 27956 16028 28008
rect 16080 27956 16086 28008
rect 16209 27999 16267 28005
rect 16209 27965 16221 27999
rect 16255 27996 16267 27999
rect 16408 27996 16436 28036
rect 16255 27968 16436 27996
rect 16255 27965 16267 27968
rect 16209 27959 16267 27965
rect 16040 27928 16068 27956
rect 17052 27937 17080 28104
rect 21082 28092 21088 28104
rect 21140 28092 21146 28144
rect 22186 28092 22192 28144
rect 22244 28132 22250 28144
rect 22244 28104 22770 28132
rect 22244 28092 22250 28104
rect 24670 28092 24676 28144
rect 24728 28092 24734 28144
rect 18233 28067 18291 28073
rect 18233 28064 18245 28067
rect 17512 28036 18245 28064
rect 17037 27931 17095 27937
rect 17037 27928 17049 27931
rect 15120 27900 15700 27928
rect 16040 27900 17049 27928
rect 9950 27860 9956 27872
rect 8404 27832 9956 27860
rect 9950 27820 9956 27832
rect 10008 27820 10014 27872
rect 10413 27863 10471 27869
rect 10413 27829 10425 27863
rect 10459 27860 10471 27863
rect 10686 27860 10692 27872
rect 10459 27832 10692 27860
rect 10459 27829 10471 27832
rect 10413 27823 10471 27829
rect 10686 27820 10692 27832
rect 10744 27820 10750 27872
rect 14918 27820 14924 27872
rect 14976 27860 14982 27872
rect 15120 27869 15148 27900
rect 15105 27863 15163 27869
rect 15105 27860 15117 27863
rect 14976 27832 15117 27860
rect 14976 27820 14982 27832
rect 15105 27829 15117 27832
rect 15151 27829 15163 27863
rect 15105 27823 15163 27829
rect 15562 27820 15568 27872
rect 15620 27820 15626 27872
rect 15672 27860 15700 27900
rect 17037 27897 17049 27900
rect 17083 27897 17095 27931
rect 17037 27891 17095 27897
rect 15838 27860 15844 27872
rect 15672 27832 15844 27860
rect 15838 27820 15844 27832
rect 15896 27860 15902 27872
rect 17512 27869 17540 28036
rect 18233 28033 18245 28036
rect 18279 28033 18291 28067
rect 18233 28027 18291 28033
rect 19334 28024 19340 28076
rect 19392 28064 19398 28076
rect 19429 28067 19487 28073
rect 19429 28064 19441 28067
rect 19392 28036 19441 28064
rect 19392 28024 19398 28036
rect 19429 28033 19441 28036
rect 19475 28033 19487 28067
rect 19429 28027 19487 28033
rect 22002 28024 22008 28076
rect 22060 28024 22066 28076
rect 18509 27999 18567 28005
rect 18509 27965 18521 27999
rect 18555 27996 18567 27999
rect 18598 27996 18604 28008
rect 18555 27968 18604 27996
rect 18555 27965 18567 27968
rect 18509 27959 18567 27965
rect 18598 27956 18604 27968
rect 18656 27996 18662 28008
rect 18782 27996 18788 28008
rect 18656 27968 18788 27996
rect 18656 27956 18662 27968
rect 18782 27956 18788 27968
rect 18840 27956 18846 28008
rect 19521 27999 19579 28005
rect 19521 27965 19533 27999
rect 19567 27965 19579 27999
rect 19521 27959 19579 27965
rect 19705 27999 19763 28005
rect 19705 27965 19717 27999
rect 19751 27996 19763 27999
rect 19978 27996 19984 28008
rect 19751 27968 19984 27996
rect 19751 27965 19763 27968
rect 19705 27959 19763 27965
rect 17497 27863 17555 27869
rect 17497 27860 17509 27863
rect 15896 27832 17509 27860
rect 15896 27820 15902 27832
rect 17497 27829 17509 27832
rect 17543 27829 17555 27863
rect 17497 27823 17555 27829
rect 17862 27820 17868 27872
rect 17920 27820 17926 27872
rect 19058 27820 19064 27872
rect 19116 27820 19122 27872
rect 19536 27860 19564 27959
rect 19978 27956 19984 27968
rect 20036 27956 20042 28008
rect 22281 27999 22339 28005
rect 22281 27965 22293 27999
rect 22327 27996 22339 27999
rect 24670 27996 24676 28008
rect 22327 27968 24676 27996
rect 22327 27965 22339 27968
rect 22281 27959 22339 27965
rect 24670 27956 24676 27968
rect 24728 27956 24734 28008
rect 24857 27931 24915 27937
rect 24857 27928 24869 27931
rect 23308 27900 24869 27928
rect 20070 27860 20076 27872
rect 19536 27832 20076 27860
rect 20070 27820 20076 27832
rect 20128 27820 20134 27872
rect 22738 27820 22744 27872
rect 22796 27860 22802 27872
rect 23308 27860 23336 27900
rect 24857 27897 24869 27900
rect 24903 27897 24915 27931
rect 24857 27891 24915 27897
rect 22796 27832 23336 27860
rect 22796 27820 22802 27832
rect 23382 27820 23388 27872
rect 23440 27860 23446 27872
rect 24121 27863 24179 27869
rect 24121 27860 24133 27863
rect 23440 27832 24133 27860
rect 23440 27820 23446 27832
rect 24121 27829 24133 27832
rect 24167 27829 24179 27863
rect 24121 27823 24179 27829
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 6444 27659 6502 27665
rect 6444 27625 6456 27659
rect 6490 27656 6502 27659
rect 9858 27656 9864 27668
rect 6490 27628 9864 27656
rect 6490 27625 6502 27628
rect 6444 27619 6502 27625
rect 9858 27616 9864 27628
rect 9916 27616 9922 27668
rect 12526 27616 12532 27668
rect 12584 27656 12590 27668
rect 13173 27659 13231 27665
rect 13173 27656 13185 27659
rect 12584 27628 13185 27656
rect 12584 27616 12590 27628
rect 13173 27625 13185 27628
rect 13219 27656 13231 27659
rect 13262 27656 13268 27668
rect 13219 27628 13268 27656
rect 13219 27625 13231 27628
rect 13173 27619 13231 27625
rect 13262 27616 13268 27628
rect 13320 27616 13326 27668
rect 18322 27616 18328 27668
rect 18380 27656 18386 27668
rect 18598 27656 18604 27668
rect 18380 27628 18604 27656
rect 18380 27616 18386 27628
rect 18598 27616 18604 27628
rect 18656 27656 18662 27668
rect 18693 27659 18751 27665
rect 18693 27656 18705 27659
rect 18656 27628 18705 27656
rect 18656 27616 18662 27628
rect 18693 27625 18705 27628
rect 18739 27625 18751 27659
rect 18693 27619 18751 27625
rect 21634 27616 21640 27668
rect 21692 27656 21698 27668
rect 22186 27656 22192 27668
rect 21692 27628 22192 27656
rect 21692 27616 21698 27628
rect 22186 27616 22192 27628
rect 22244 27656 22250 27668
rect 22830 27656 22836 27668
rect 22244 27628 22836 27656
rect 22244 27616 22250 27628
rect 22830 27616 22836 27628
rect 22888 27656 22894 27668
rect 23382 27656 23388 27668
rect 22888 27628 23388 27656
rect 22888 27616 22894 27628
rect 23382 27616 23388 27628
rect 23440 27616 23446 27668
rect 24210 27616 24216 27668
rect 24268 27616 24274 27668
rect 7834 27548 7840 27600
rect 7892 27588 7898 27600
rect 7929 27591 7987 27597
rect 7929 27588 7941 27591
rect 7892 27560 7941 27588
rect 7892 27548 7898 27560
rect 7929 27557 7941 27560
rect 7975 27557 7987 27591
rect 7929 27551 7987 27557
rect 8294 27548 8300 27600
rect 8352 27588 8358 27600
rect 8389 27591 8447 27597
rect 8389 27588 8401 27591
rect 8352 27560 8401 27588
rect 8352 27548 8358 27560
rect 8389 27557 8401 27560
rect 8435 27557 8447 27591
rect 8389 27551 8447 27557
rect 18141 27591 18199 27597
rect 18141 27557 18153 27591
rect 18187 27588 18199 27591
rect 21542 27588 21548 27600
rect 18187 27560 21548 27588
rect 18187 27557 18199 27560
rect 18141 27551 18199 27557
rect 21542 27548 21548 27560
rect 21600 27548 21606 27600
rect 6181 27523 6239 27529
rect 6181 27489 6193 27523
rect 6227 27520 6239 27523
rect 6546 27520 6552 27532
rect 6227 27492 6552 27520
rect 6227 27489 6239 27492
rect 6181 27483 6239 27489
rect 6546 27480 6552 27492
rect 6604 27480 6610 27532
rect 12066 27520 12072 27532
rect 11164 27492 12072 27520
rect 9950 27412 9956 27464
rect 10008 27452 10014 27464
rect 11164 27461 11192 27492
rect 12066 27480 12072 27492
rect 12124 27480 12130 27532
rect 12802 27480 12808 27532
rect 12860 27520 12866 27532
rect 15657 27523 15715 27529
rect 15657 27520 15669 27523
rect 12860 27492 15669 27520
rect 12860 27480 12866 27492
rect 15657 27489 15669 27492
rect 15703 27489 15715 27523
rect 15657 27483 15715 27489
rect 16393 27523 16451 27529
rect 16393 27489 16405 27523
rect 16439 27520 16451 27523
rect 16439 27492 18460 27520
rect 16439 27489 16451 27492
rect 16393 27483 16451 27489
rect 11149 27455 11207 27461
rect 11149 27452 11161 27455
rect 10008 27424 11161 27452
rect 10008 27412 10014 27424
rect 11149 27421 11161 27424
rect 11195 27421 11207 27455
rect 11149 27415 11207 27421
rect 12526 27412 12532 27464
rect 12584 27412 12590 27464
rect 15473 27455 15531 27461
rect 15473 27421 15485 27455
rect 15519 27452 15531 27455
rect 15838 27452 15844 27464
rect 15519 27424 15844 27452
rect 15519 27421 15531 27424
rect 15473 27415 15531 27421
rect 15838 27412 15844 27424
rect 15896 27452 15902 27464
rect 16408 27452 16436 27483
rect 15896 27424 16436 27452
rect 15896 27412 15902 27424
rect 17678 27412 17684 27464
rect 17736 27452 17742 27464
rect 18325 27455 18383 27461
rect 18325 27452 18337 27455
rect 17736 27424 18337 27452
rect 17736 27412 17742 27424
rect 18325 27421 18337 27424
rect 18371 27421 18383 27455
rect 18432 27452 18460 27492
rect 20438 27480 20444 27532
rect 20496 27520 20502 27532
rect 20533 27523 20591 27529
rect 20533 27520 20545 27523
rect 20496 27492 20545 27520
rect 20496 27480 20502 27492
rect 20533 27489 20545 27492
rect 20579 27489 20591 27523
rect 20533 27483 20591 27489
rect 20622 27480 20628 27532
rect 20680 27480 20686 27532
rect 21910 27480 21916 27532
rect 21968 27480 21974 27532
rect 22646 27480 22652 27532
rect 22704 27520 22710 27532
rect 22704 27492 24716 27520
rect 22704 27480 22710 27492
rect 21266 27452 21272 27464
rect 18432 27424 21272 27452
rect 18325 27415 18383 27421
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 24688 27461 24716 27492
rect 24673 27455 24731 27461
rect 24673 27421 24685 27455
rect 24719 27421 24731 27455
rect 24673 27415 24731 27421
rect 8294 27384 8300 27396
rect 7682 27356 8300 27384
rect 8294 27344 8300 27356
rect 8352 27344 8358 27396
rect 11422 27344 11428 27396
rect 11480 27344 11486 27396
rect 15378 27344 15384 27396
rect 15436 27384 15442 27396
rect 15565 27387 15623 27393
rect 15565 27384 15577 27387
rect 15436 27356 15577 27384
rect 15436 27344 15442 27356
rect 15565 27353 15577 27356
rect 15611 27384 15623 27387
rect 16117 27387 16175 27393
rect 16117 27384 16129 27387
rect 15611 27356 16129 27384
rect 15611 27353 15623 27356
rect 15565 27347 15623 27353
rect 16117 27353 16129 27356
rect 16163 27384 16175 27387
rect 16163 27356 17080 27384
rect 16163 27353 16175 27356
rect 16117 27347 16175 27353
rect 10226 27276 10232 27328
rect 10284 27316 10290 27328
rect 12894 27316 12900 27328
rect 10284 27288 12900 27316
rect 10284 27276 10290 27288
rect 12894 27276 12900 27288
rect 12952 27276 12958 27328
rect 15010 27276 15016 27328
rect 15068 27316 15074 27328
rect 15105 27319 15163 27325
rect 15105 27316 15117 27319
rect 15068 27288 15117 27316
rect 15068 27276 15074 27288
rect 15105 27285 15117 27288
rect 15151 27285 15163 27319
rect 17052 27316 17080 27356
rect 17218 27344 17224 27396
rect 17276 27384 17282 27396
rect 19705 27387 19763 27393
rect 19705 27384 19717 27387
rect 17276 27356 19717 27384
rect 17276 27344 17282 27356
rect 19705 27353 19717 27356
rect 19751 27384 19763 27387
rect 20441 27387 20499 27393
rect 20441 27384 20453 27387
rect 19751 27356 20453 27384
rect 19751 27353 19763 27356
rect 19705 27347 19763 27353
rect 20441 27353 20453 27356
rect 20487 27353 20499 27387
rect 22094 27384 22100 27396
rect 20441 27347 20499 27353
rect 21100 27356 22100 27384
rect 17126 27316 17132 27328
rect 17052 27288 17132 27316
rect 15105 27279 15163 27285
rect 17126 27276 17132 27288
rect 17184 27316 17190 27328
rect 18877 27319 18935 27325
rect 18877 27316 18889 27319
rect 17184 27288 18889 27316
rect 17184 27276 17190 27288
rect 18877 27285 18889 27288
rect 18923 27316 18935 27319
rect 19334 27316 19340 27328
rect 18923 27288 19340 27316
rect 18923 27285 18935 27288
rect 18877 27279 18935 27285
rect 19334 27276 19340 27288
rect 19392 27276 19398 27328
rect 20073 27319 20131 27325
rect 20073 27285 20085 27319
rect 20119 27316 20131 27319
rect 21100 27316 21128 27356
rect 22094 27344 22100 27356
rect 22152 27344 22158 27396
rect 22186 27344 22192 27396
rect 22244 27344 22250 27396
rect 22830 27344 22836 27396
rect 22888 27344 22894 27396
rect 24857 27387 24915 27393
rect 24857 27353 24869 27387
rect 24903 27384 24915 27387
rect 25590 27384 25596 27396
rect 24903 27356 25596 27384
rect 24903 27353 24915 27356
rect 24857 27347 24915 27353
rect 25590 27344 25596 27356
rect 25648 27344 25654 27396
rect 20119 27288 21128 27316
rect 20119 27285 20131 27288
rect 20073 27279 20131 27285
rect 23106 27276 23112 27328
rect 23164 27316 23170 27328
rect 23661 27319 23719 27325
rect 23661 27316 23673 27319
rect 23164 27288 23673 27316
rect 23164 27276 23170 27288
rect 23661 27285 23673 27288
rect 23707 27285 23719 27319
rect 23661 27279 23719 27285
rect 25222 27276 25228 27328
rect 25280 27276 25286 27328
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 3191 27115 3249 27121
rect 3191 27081 3203 27115
rect 3237 27112 3249 27115
rect 3418 27112 3424 27124
rect 3237 27084 3424 27112
rect 3237 27081 3249 27084
rect 3191 27075 3249 27081
rect 3418 27072 3424 27084
rect 3476 27072 3482 27124
rect 10686 27072 10692 27124
rect 10744 27112 10750 27124
rect 11793 27115 11851 27121
rect 11793 27112 11805 27115
rect 10744 27084 11805 27112
rect 10744 27072 10750 27084
rect 11793 27081 11805 27084
rect 11839 27112 11851 27115
rect 11839 27084 12020 27112
rect 11839 27081 11851 27084
rect 11793 27075 11851 27081
rect 1578 27004 1584 27056
rect 1636 27044 1642 27056
rect 3789 27047 3847 27053
rect 3789 27044 3801 27047
rect 1636 27016 3801 27044
rect 1636 27004 1642 27016
rect 3789 27013 3801 27016
rect 3835 27013 3847 27047
rect 3789 27007 3847 27013
rect 3881 27047 3939 27053
rect 3881 27013 3893 27047
rect 3927 27044 3939 27047
rect 4338 27044 4344 27056
rect 3927 27016 4344 27044
rect 3927 27013 3939 27016
rect 3881 27007 3939 27013
rect 4338 27004 4344 27016
rect 4396 27004 4402 27056
rect 8110 27044 8116 27056
rect 8050 27016 8116 27044
rect 8110 27004 8116 27016
rect 8168 27044 8174 27056
rect 8294 27044 8300 27056
rect 8168 27016 8300 27044
rect 8168 27004 8174 27016
rect 8294 27004 8300 27016
rect 8352 27004 8358 27056
rect 10505 27047 10563 27053
rect 10505 27013 10517 27047
rect 10551 27044 10563 27047
rect 11238 27044 11244 27056
rect 10551 27016 11244 27044
rect 10551 27013 10563 27016
rect 10505 27007 10563 27013
rect 11238 27004 11244 27016
rect 11296 27004 11302 27056
rect 3120 26979 3178 26985
rect 3120 26945 3132 26979
rect 3166 26976 3178 26979
rect 3418 26976 3424 26988
rect 3166 26948 3424 26976
rect 3166 26945 3178 26948
rect 3120 26939 3178 26945
rect 3418 26936 3424 26948
rect 3476 26936 3482 26988
rect 6546 26936 6552 26988
rect 6604 26936 6610 26988
rect 9122 26936 9128 26988
rect 9180 26936 9186 26988
rect 4433 26911 4491 26917
rect 4433 26877 4445 26911
rect 4479 26908 4491 26911
rect 6825 26911 6883 26917
rect 4479 26880 4568 26908
rect 4479 26877 4491 26880
rect 4433 26871 4491 26877
rect 4540 26852 4568 26880
rect 6825 26877 6837 26911
rect 6871 26908 6883 26911
rect 7834 26908 7840 26920
rect 6871 26880 7840 26908
rect 6871 26877 6883 26880
rect 6825 26871 6883 26877
rect 7834 26868 7840 26880
rect 7892 26868 7898 26920
rect 8662 26868 8668 26920
rect 8720 26908 8726 26920
rect 9217 26911 9275 26917
rect 9217 26908 9229 26911
rect 8720 26880 9229 26908
rect 8720 26868 8726 26880
rect 9217 26877 9229 26880
rect 9263 26877 9275 26911
rect 9217 26871 9275 26877
rect 9398 26868 9404 26920
rect 9456 26868 9462 26920
rect 4522 26800 4528 26852
rect 4580 26800 4586 26852
rect 8294 26800 8300 26852
rect 8352 26840 8358 26852
rect 9674 26840 9680 26852
rect 8352 26812 9680 26840
rect 8352 26800 8358 26812
rect 9674 26800 9680 26812
rect 9732 26800 9738 26852
rect 10134 26800 10140 26852
rect 10192 26840 10198 26852
rect 10689 26843 10747 26849
rect 10689 26840 10701 26843
rect 10192 26812 10701 26840
rect 10192 26800 10198 26812
rect 10689 26809 10701 26812
rect 10735 26809 10747 26843
rect 11992 26840 12020 27084
rect 12894 27072 12900 27124
rect 12952 27112 12958 27124
rect 12952 27084 14136 27112
rect 12952 27072 12958 27084
rect 12066 27004 12072 27056
rect 12124 27044 12130 27056
rect 12124 27016 12388 27044
rect 12124 27004 12130 27016
rect 12360 26976 12388 27016
rect 12802 27004 12808 27056
rect 12860 27004 12866 27056
rect 13262 27004 13268 27056
rect 13320 27004 13326 27056
rect 14108 27044 14136 27084
rect 15102 27072 15108 27124
rect 15160 27112 15166 27124
rect 15197 27115 15255 27121
rect 15197 27112 15209 27115
rect 15160 27084 15209 27112
rect 15160 27072 15166 27084
rect 15197 27081 15209 27084
rect 15243 27081 15255 27115
rect 15197 27075 15255 27081
rect 17589 27115 17647 27121
rect 17589 27081 17601 27115
rect 17635 27112 17647 27115
rect 19981 27115 20039 27121
rect 19981 27112 19993 27115
rect 17635 27084 19993 27112
rect 17635 27081 17647 27084
rect 17589 27075 17647 27081
rect 19981 27081 19993 27084
rect 20027 27081 20039 27115
rect 19981 27075 20039 27081
rect 20162 27072 20168 27124
rect 20220 27112 20226 27124
rect 20438 27112 20444 27124
rect 20220 27084 20444 27112
rect 20220 27072 20226 27084
rect 20438 27072 20444 27084
rect 20496 27072 20502 27124
rect 24578 27112 24584 27124
rect 22848 27084 24584 27112
rect 18049 27047 18107 27053
rect 14108 27016 15332 27044
rect 12529 26979 12587 26985
rect 12529 26976 12541 26979
rect 12360 26948 12541 26976
rect 12529 26945 12541 26948
rect 12575 26945 12587 26979
rect 12529 26939 12587 26945
rect 14182 26936 14188 26988
rect 14240 26976 14246 26988
rect 15105 26979 15163 26985
rect 15105 26976 15117 26979
rect 14240 26948 15117 26976
rect 14240 26936 14246 26948
rect 15105 26945 15117 26948
rect 15151 26945 15163 26979
rect 15105 26939 15163 26945
rect 15304 26917 15332 27016
rect 18049 27013 18061 27047
rect 18095 27044 18107 27047
rect 18966 27044 18972 27056
rect 18095 27016 18972 27044
rect 18095 27013 18107 27016
rect 18049 27007 18107 27013
rect 18966 27004 18972 27016
rect 19024 27004 19030 27056
rect 17957 26979 18015 26985
rect 17957 26945 17969 26979
rect 18003 26945 18015 26979
rect 17957 26939 18015 26945
rect 19889 26979 19947 26985
rect 19889 26945 19901 26979
rect 19935 26976 19947 26979
rect 20717 26979 20775 26985
rect 20717 26976 20729 26979
rect 19935 26948 20729 26976
rect 19935 26945 19947 26948
rect 19889 26939 19947 26945
rect 20717 26945 20729 26948
rect 20763 26945 20775 26979
rect 20717 26939 20775 26945
rect 22373 26979 22431 26985
rect 22373 26945 22385 26979
rect 22419 26976 22431 26979
rect 22848 26976 22876 27084
rect 24578 27072 24584 27084
rect 24636 27072 24642 27124
rect 23106 27004 23112 27056
rect 23164 27004 23170 27056
rect 23382 27004 23388 27056
rect 23440 27044 23446 27056
rect 23440 27016 23598 27044
rect 23440 27004 23446 27016
rect 25130 27004 25136 27056
rect 25188 27004 25194 27056
rect 22419 26948 22876 26976
rect 22419 26945 22431 26948
rect 22373 26939 22431 26945
rect 15289 26911 15347 26917
rect 15289 26877 15301 26911
rect 15335 26877 15347 26911
rect 15289 26871 15347 26877
rect 12526 26840 12532 26852
rect 11992 26812 12532 26840
rect 10689 26803 10747 26809
rect 12526 26800 12532 26812
rect 12584 26800 12590 26852
rect 8757 26775 8815 26781
rect 8757 26741 8769 26775
rect 8803 26772 8815 26775
rect 10502 26772 10508 26784
rect 8803 26744 10508 26772
rect 8803 26741 8815 26744
rect 8757 26735 8815 26741
rect 10502 26732 10508 26744
rect 10560 26732 10566 26784
rect 10594 26732 10600 26784
rect 10652 26772 10658 26784
rect 12342 26772 12348 26784
rect 10652 26744 12348 26772
rect 10652 26732 10658 26744
rect 12342 26732 12348 26744
rect 12400 26732 12406 26784
rect 14277 26775 14335 26781
rect 14277 26741 14289 26775
rect 14323 26772 14335 26775
rect 14366 26772 14372 26784
rect 14323 26744 14372 26772
rect 14323 26741 14335 26744
rect 14277 26735 14335 26741
rect 14366 26732 14372 26744
rect 14424 26732 14430 26784
rect 14734 26732 14740 26784
rect 14792 26732 14798 26784
rect 17313 26775 17371 26781
rect 17313 26741 17325 26775
rect 17359 26772 17371 26775
rect 17972 26772 18000 26939
rect 18233 26911 18291 26917
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 19334 26908 19340 26920
rect 18279 26880 19340 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 19334 26868 19340 26880
rect 19392 26908 19398 26920
rect 19518 26908 19524 26920
rect 19392 26880 19524 26908
rect 19392 26868 19398 26880
rect 19518 26868 19524 26880
rect 19576 26868 19582 26920
rect 20165 26911 20223 26917
rect 20165 26877 20177 26911
rect 20211 26908 20223 26911
rect 21174 26908 21180 26920
rect 20211 26880 21180 26908
rect 20211 26877 20223 26880
rect 20165 26871 20223 26877
rect 21174 26868 21180 26880
rect 21232 26868 21238 26920
rect 22002 26868 22008 26920
rect 22060 26908 22066 26920
rect 22833 26911 22891 26917
rect 22833 26908 22845 26911
rect 22060 26880 22845 26908
rect 22060 26868 22066 26880
rect 22833 26877 22845 26880
rect 22879 26877 22891 26911
rect 23106 26908 23112 26920
rect 22833 26871 22891 26877
rect 22940 26880 23112 26908
rect 20622 26800 20628 26852
rect 20680 26840 20686 26852
rect 22940 26840 22968 26880
rect 23106 26868 23112 26880
rect 23164 26868 23170 26920
rect 23474 26868 23480 26920
rect 23532 26908 23538 26920
rect 24581 26911 24639 26917
rect 24581 26908 24593 26911
rect 23532 26880 24593 26908
rect 23532 26868 23538 26880
rect 24581 26877 24593 26880
rect 24627 26877 24639 26911
rect 24581 26871 24639 26877
rect 20680 26812 22968 26840
rect 25317 26843 25375 26849
rect 20680 26800 20686 26812
rect 25317 26809 25329 26843
rect 25363 26840 25375 26843
rect 25406 26840 25412 26852
rect 25363 26812 25412 26840
rect 25363 26809 25375 26812
rect 25317 26803 25375 26809
rect 25406 26800 25412 26812
rect 25464 26800 25470 26852
rect 18322 26772 18328 26784
rect 17359 26744 18328 26772
rect 17359 26741 17371 26744
rect 17313 26735 17371 26741
rect 18322 26732 18328 26744
rect 18380 26732 18386 26784
rect 19518 26732 19524 26784
rect 19576 26732 19582 26784
rect 22189 26775 22247 26781
rect 22189 26741 22201 26775
rect 22235 26772 22247 26775
rect 23842 26772 23848 26784
rect 22235 26744 23848 26772
rect 22235 26741 22247 26744
rect 22189 26735 22247 26741
rect 23842 26732 23848 26744
rect 23900 26732 23906 26784
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 4062 26528 4068 26580
rect 4120 26528 4126 26580
rect 7098 26528 7104 26580
rect 7156 26568 7162 26580
rect 7742 26568 7748 26580
rect 7156 26540 7748 26568
rect 7156 26528 7162 26540
rect 7742 26528 7748 26540
rect 7800 26568 7806 26580
rect 8205 26571 8263 26577
rect 8205 26568 8217 26571
rect 7800 26540 8217 26568
rect 7800 26528 7806 26540
rect 8205 26537 8217 26540
rect 8251 26537 8263 26571
rect 8205 26531 8263 26537
rect 9214 26528 9220 26580
rect 9272 26568 9278 26580
rect 9272 26540 11468 26568
rect 9272 26528 9278 26540
rect 6454 26392 6460 26444
rect 6512 26392 6518 26444
rect 6733 26435 6791 26441
rect 6733 26401 6745 26435
rect 6779 26432 6791 26435
rect 8294 26432 8300 26444
rect 6779 26404 8300 26432
rect 6779 26401 6791 26404
rect 6733 26395 6791 26401
rect 8294 26392 8300 26404
rect 8352 26392 8358 26444
rect 9122 26392 9128 26444
rect 9180 26392 9186 26444
rect 10226 26392 10232 26444
rect 10284 26392 10290 26444
rect 1765 26367 1823 26373
rect 1765 26333 1777 26367
rect 1811 26364 1823 26367
rect 2038 26364 2044 26376
rect 1811 26336 2044 26364
rect 1811 26333 1823 26336
rect 1765 26327 1823 26333
rect 2038 26324 2044 26336
rect 2096 26324 2102 26376
rect 9950 26324 9956 26376
rect 10008 26324 10014 26376
rect 11440 26364 11468 26540
rect 12526 26528 12532 26580
rect 12584 26568 12590 26580
rect 14369 26571 14427 26577
rect 14369 26568 14381 26571
rect 12584 26540 14381 26568
rect 12584 26528 12590 26540
rect 14369 26537 14381 26540
rect 14415 26568 14427 26571
rect 14642 26568 14648 26580
rect 14415 26540 14648 26568
rect 14415 26537 14427 26540
rect 14369 26531 14427 26537
rect 14642 26528 14648 26540
rect 14700 26528 14706 26580
rect 16666 26528 16672 26580
rect 16724 26568 16730 26580
rect 17129 26571 17187 26577
rect 17129 26568 17141 26571
rect 16724 26540 17141 26568
rect 16724 26528 16730 26540
rect 17129 26537 17141 26540
rect 17175 26568 17187 26571
rect 17770 26568 17776 26580
rect 17175 26540 17776 26568
rect 17175 26537 17187 26540
rect 17129 26531 17187 26537
rect 17770 26528 17776 26540
rect 17828 26528 17834 26580
rect 21910 26528 21916 26580
rect 21968 26568 21974 26580
rect 21968 26540 23244 26568
rect 21968 26528 21974 26540
rect 12161 26503 12219 26509
rect 12161 26469 12173 26503
rect 12207 26500 12219 26503
rect 12250 26500 12256 26512
rect 12207 26472 12256 26500
rect 12207 26469 12219 26472
rect 12161 26463 12219 26469
rect 12250 26460 12256 26472
rect 12308 26460 12314 26512
rect 12342 26460 12348 26512
rect 12400 26500 12406 26512
rect 19429 26503 19487 26509
rect 12400 26460 12434 26500
rect 19429 26469 19441 26503
rect 19475 26500 19487 26503
rect 19702 26500 19708 26512
rect 19475 26472 19708 26500
rect 19475 26469 19487 26472
rect 19429 26463 19487 26469
rect 19702 26460 19708 26472
rect 19760 26460 19766 26512
rect 22002 26460 22008 26512
rect 22060 26460 22066 26512
rect 22186 26460 22192 26512
rect 22244 26500 22250 26512
rect 22373 26503 22431 26509
rect 22373 26500 22385 26503
rect 22244 26472 22385 26500
rect 22244 26460 22250 26472
rect 22373 26469 22385 26472
rect 22419 26469 22431 26503
rect 22373 26463 22431 26469
rect 22554 26460 22560 26512
rect 22612 26500 22618 26512
rect 22833 26503 22891 26509
rect 22833 26500 22845 26503
rect 22612 26472 22845 26500
rect 22612 26460 22618 26472
rect 22833 26469 22845 26472
rect 22879 26469 22891 26503
rect 22833 26463 22891 26469
rect 12406 26432 12434 26460
rect 12713 26435 12771 26441
rect 12713 26432 12725 26435
rect 12406 26404 12725 26432
rect 12713 26401 12725 26404
rect 12759 26401 12771 26435
rect 12713 26395 12771 26401
rect 15657 26435 15715 26441
rect 15657 26401 15669 26435
rect 15703 26432 15715 26435
rect 17034 26432 17040 26444
rect 15703 26404 17040 26432
rect 15703 26401 15715 26404
rect 15657 26395 15715 26401
rect 17034 26392 17040 26404
rect 17092 26432 17098 26444
rect 17092 26404 17540 26432
rect 17092 26392 17098 26404
rect 12529 26367 12587 26373
rect 12529 26364 12541 26367
rect 11440 26336 12541 26364
rect 12529 26333 12541 26336
rect 12575 26333 12587 26367
rect 12529 26327 12587 26333
rect 12621 26367 12679 26373
rect 12621 26333 12633 26367
rect 12667 26364 12679 26367
rect 14274 26364 14280 26376
rect 12667 26336 14280 26364
rect 12667 26333 12679 26336
rect 12621 26327 12679 26333
rect 14274 26324 14280 26336
rect 14332 26324 14338 26376
rect 15378 26324 15384 26376
rect 15436 26324 15442 26376
rect 2774 26256 2780 26308
rect 2832 26256 2838 26308
rect 8110 26296 8116 26308
rect 7958 26268 8116 26296
rect 8110 26256 8116 26268
rect 8168 26296 8174 26308
rect 8478 26296 8484 26308
rect 8168 26268 8484 26296
rect 8168 26256 8174 26268
rect 8478 26256 8484 26268
rect 8536 26256 8542 26308
rect 8662 26256 8668 26308
rect 8720 26256 8726 26308
rect 9582 26256 9588 26308
rect 9640 26296 9646 26308
rect 9640 26268 10640 26296
rect 9640 26256 9646 26268
rect 10612 26228 10640 26268
rect 10686 26256 10692 26308
rect 10744 26256 10750 26308
rect 14826 26296 14832 26308
rect 11716 26268 14832 26296
rect 11716 26237 11744 26268
rect 14826 26256 14832 26268
rect 14884 26256 14890 26308
rect 17512 26305 17540 26404
rect 17862 26392 17868 26444
rect 17920 26432 17926 26444
rect 19889 26435 19947 26441
rect 19889 26432 19901 26435
rect 17920 26404 19901 26432
rect 17920 26392 17926 26404
rect 19889 26401 19901 26404
rect 19935 26401 19947 26435
rect 19889 26395 19947 26401
rect 20073 26435 20131 26441
rect 20073 26401 20085 26435
rect 20119 26432 20131 26435
rect 20162 26432 20168 26444
rect 20119 26404 20168 26432
rect 20119 26401 20131 26404
rect 20073 26395 20131 26401
rect 20162 26392 20168 26404
rect 20220 26392 20226 26444
rect 20625 26435 20683 26441
rect 20625 26401 20637 26435
rect 20671 26432 20683 26435
rect 22020 26432 22048 26460
rect 20671 26404 22048 26432
rect 20671 26401 20683 26404
rect 20625 26395 20683 26401
rect 19797 26367 19855 26373
rect 19797 26333 19809 26367
rect 19843 26364 19855 26367
rect 20254 26364 20260 26376
rect 19843 26336 20260 26364
rect 19843 26333 19855 26336
rect 19797 26327 19855 26333
rect 20254 26324 20260 26336
rect 20312 26324 20318 26376
rect 23216 26373 23244 26540
rect 23566 26528 23572 26580
rect 23624 26568 23630 26580
rect 23845 26571 23903 26577
rect 23845 26568 23857 26571
rect 23624 26540 23857 26568
rect 23624 26528 23630 26540
rect 23845 26537 23857 26540
rect 23891 26568 23903 26571
rect 25038 26568 25044 26580
rect 23891 26540 25044 26568
rect 23891 26537 23903 26540
rect 23845 26531 23903 26537
rect 25038 26528 25044 26540
rect 25096 26568 25102 26580
rect 25133 26571 25191 26577
rect 25133 26568 25145 26571
rect 25096 26540 25145 26568
rect 25096 26528 25102 26540
rect 25133 26537 25145 26540
rect 25179 26568 25191 26571
rect 25222 26568 25228 26580
rect 25179 26540 25228 26568
rect 25179 26537 25191 26540
rect 25133 26531 25191 26537
rect 25222 26528 25228 26540
rect 25280 26528 25286 26580
rect 23477 26435 23535 26441
rect 23477 26401 23489 26435
rect 23523 26432 23535 26435
rect 24486 26432 24492 26444
rect 23523 26404 24492 26432
rect 23523 26401 23535 26404
rect 23477 26395 23535 26401
rect 24486 26392 24492 26404
rect 24544 26392 24550 26444
rect 23201 26367 23259 26373
rect 23201 26333 23213 26367
rect 23247 26333 23259 26367
rect 23201 26327 23259 26333
rect 24394 26324 24400 26376
rect 24452 26364 24458 26376
rect 24673 26367 24731 26373
rect 24673 26364 24685 26367
rect 24452 26336 24685 26364
rect 24452 26324 24458 26336
rect 24673 26333 24685 26336
rect 24719 26333 24731 26367
rect 24673 26327 24731 26333
rect 17497 26299 17555 26305
rect 16040 26268 16146 26296
rect 11701 26231 11759 26237
rect 11701 26228 11713 26231
rect 10612 26200 11713 26228
rect 11701 26197 11713 26200
rect 11747 26197 11759 26231
rect 11701 26191 11759 26197
rect 14642 26188 14648 26240
rect 14700 26228 14706 26240
rect 16040 26228 16068 26268
rect 17497 26265 17509 26299
rect 17543 26296 17555 26299
rect 17678 26296 17684 26308
rect 17543 26268 17684 26296
rect 17543 26265 17555 26268
rect 17497 26259 17555 26265
rect 17678 26256 17684 26268
rect 17736 26256 17742 26308
rect 20901 26299 20959 26305
rect 20901 26265 20913 26299
rect 20947 26296 20959 26299
rect 21174 26296 21180 26308
rect 20947 26268 21180 26296
rect 20947 26265 20959 26268
rect 20901 26259 20959 26265
rect 21174 26256 21180 26268
rect 21232 26256 21238 26308
rect 21634 26256 21640 26308
rect 21692 26256 21698 26308
rect 22462 26256 22468 26308
rect 22520 26296 22526 26308
rect 23293 26299 23351 26305
rect 23293 26296 23305 26299
rect 22520 26268 23305 26296
rect 22520 26256 22526 26268
rect 23293 26265 23305 26268
rect 23339 26265 23351 26299
rect 23293 26259 23351 26265
rect 24857 26299 24915 26305
rect 24857 26265 24869 26299
rect 24903 26296 24915 26299
rect 25222 26296 25228 26308
rect 24903 26268 25228 26296
rect 24903 26265 24915 26268
rect 24857 26259 24915 26265
rect 25222 26256 25228 26268
rect 25280 26256 25286 26308
rect 17586 26228 17592 26240
rect 14700 26200 17592 26228
rect 14700 26188 14706 26200
rect 17586 26188 17592 26200
rect 17644 26188 17650 26240
rect 22646 26188 22652 26240
rect 22704 26228 22710 26240
rect 23382 26228 23388 26240
rect 22704 26200 23388 26228
rect 22704 26188 22710 26200
rect 23382 26188 23388 26200
rect 23440 26188 23446 26240
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 1762 25984 1768 26036
rect 1820 26024 1826 26036
rect 2133 26027 2191 26033
rect 2133 26024 2145 26027
rect 1820 25996 2145 26024
rect 1820 25984 1826 25996
rect 2133 25993 2145 25996
rect 2179 25993 2191 26027
rect 2133 25987 2191 25993
rect 6730 25984 6736 26036
rect 6788 26024 6794 26036
rect 8846 26024 8852 26036
rect 6788 25996 8852 26024
rect 6788 25984 6794 25996
rect 8846 25984 8852 25996
rect 8904 25984 8910 26036
rect 9214 25984 9220 26036
rect 9272 25984 9278 26036
rect 10502 25984 10508 26036
rect 10560 26024 10566 26036
rect 10781 26027 10839 26033
rect 10781 26024 10793 26027
rect 10560 25996 10793 26024
rect 10560 25984 10566 25996
rect 10781 25993 10793 25996
rect 10827 25993 10839 26027
rect 10781 25987 10839 25993
rect 10870 25984 10876 26036
rect 10928 25984 10934 26036
rect 15378 26024 15384 26036
rect 12728 25996 15384 26024
rect 3510 25916 3516 25968
rect 3568 25956 3574 25968
rect 4062 25956 4068 25968
rect 3568 25928 4068 25956
rect 3568 25916 3574 25928
rect 4062 25916 4068 25928
rect 4120 25956 4126 25968
rect 4120 25928 4200 25956
rect 4120 25916 4126 25928
rect 2317 25891 2375 25897
rect 2317 25857 2329 25891
rect 2363 25888 2375 25891
rect 2866 25888 2872 25900
rect 2363 25860 2872 25888
rect 2363 25857 2375 25860
rect 2317 25851 2375 25857
rect 2866 25848 2872 25860
rect 2924 25848 2930 25900
rect 4172 25897 4200 25928
rect 8478 25916 8484 25968
rect 8536 25916 8542 25968
rect 9766 25916 9772 25968
rect 9824 25956 9830 25968
rect 10686 25956 10692 25968
rect 9824 25928 10692 25956
rect 9824 25916 9830 25928
rect 10686 25916 10692 25928
rect 10744 25916 10750 25968
rect 3053 25891 3111 25897
rect 3053 25857 3065 25891
rect 3099 25888 3111 25891
rect 4157 25891 4215 25897
rect 3099 25860 4108 25888
rect 3099 25857 3111 25860
rect 3053 25851 3111 25857
rect 2774 25780 2780 25832
rect 2832 25820 2838 25832
rect 3237 25823 3295 25829
rect 3237 25820 3249 25823
rect 2832 25792 3249 25820
rect 2832 25780 2838 25792
rect 3237 25789 3249 25792
rect 3283 25820 3295 25823
rect 3602 25820 3608 25832
rect 3283 25792 3608 25820
rect 3283 25789 3295 25792
rect 3237 25783 3295 25789
rect 3602 25780 3608 25792
rect 3660 25780 3666 25832
rect 4080 25820 4108 25860
rect 4157 25857 4169 25891
rect 4203 25857 4215 25891
rect 4157 25851 4215 25857
rect 9398 25848 9404 25900
rect 9456 25888 9462 25900
rect 12728 25897 12756 25996
rect 15378 25984 15384 25996
rect 15436 25984 15442 26036
rect 15562 25984 15568 26036
rect 15620 26024 15626 26036
rect 15841 26027 15899 26033
rect 15841 26024 15853 26027
rect 15620 25996 15853 26024
rect 15620 25984 15626 25996
rect 15841 25993 15853 25996
rect 15887 25993 15899 26027
rect 15841 25987 15899 25993
rect 17586 25984 17592 26036
rect 17644 26024 17650 26036
rect 17644 25996 17724 26024
rect 17644 25984 17650 25996
rect 14642 25956 14648 25968
rect 14214 25928 14648 25956
rect 14642 25916 14648 25928
rect 14700 25956 14706 25968
rect 14737 25959 14795 25965
rect 14737 25956 14749 25959
rect 14700 25928 14749 25956
rect 14700 25916 14706 25928
rect 14737 25925 14749 25928
rect 14783 25925 14795 25959
rect 15396 25956 15424 25984
rect 17696 25956 17724 25996
rect 18248 25996 19196 26024
rect 18248 25956 18276 25996
rect 19168 25956 19196 25996
rect 19334 25984 19340 26036
rect 19392 25984 19398 26036
rect 19518 25984 19524 26036
rect 19576 26024 19582 26036
rect 20257 26027 20315 26033
rect 20257 26024 20269 26027
rect 19576 25996 20269 26024
rect 19576 25984 19582 25996
rect 20257 25993 20269 25996
rect 20303 25993 20315 26027
rect 20257 25987 20315 25993
rect 20346 25984 20352 26036
rect 20404 25984 20410 26036
rect 22370 25984 22376 26036
rect 22428 26024 22434 26036
rect 22465 26027 22523 26033
rect 22465 26024 22477 26027
rect 22428 25996 22477 26024
rect 22428 25984 22434 25996
rect 22465 25993 22477 25996
rect 22511 25993 22523 26027
rect 22465 25987 22523 25993
rect 20901 25959 20959 25965
rect 20901 25956 20913 25959
rect 15396 25928 17632 25956
rect 17696 25928 18354 25956
rect 19168 25928 20913 25956
rect 14737 25919 14795 25925
rect 17604 25897 17632 25928
rect 20901 25925 20913 25928
rect 20947 25925 20959 25959
rect 20901 25919 20959 25925
rect 21358 25916 21364 25968
rect 21416 25956 21422 25968
rect 23293 25959 23351 25965
rect 23293 25956 23305 25959
rect 21416 25928 23305 25956
rect 21416 25916 21422 25928
rect 23293 25925 23305 25928
rect 23339 25925 23351 25959
rect 23293 25919 23351 25925
rect 9585 25891 9643 25897
rect 9585 25888 9597 25891
rect 9456 25860 9597 25888
rect 9456 25848 9462 25860
rect 9585 25857 9597 25860
rect 9631 25857 9643 25891
rect 9585 25851 9643 25857
rect 12713 25891 12771 25897
rect 12713 25857 12725 25891
rect 12759 25857 12771 25891
rect 12713 25851 12771 25857
rect 15749 25891 15807 25897
rect 15749 25857 15761 25891
rect 15795 25857 15807 25891
rect 15749 25851 15807 25857
rect 17589 25891 17647 25897
rect 17589 25857 17601 25891
rect 17635 25857 17647 25891
rect 22186 25888 22192 25900
rect 17589 25851 17647 25857
rect 20548 25860 22192 25888
rect 6178 25820 6184 25832
rect 4080 25792 6184 25820
rect 6178 25780 6184 25792
rect 6236 25780 6242 25832
rect 7834 25780 7840 25832
rect 7892 25820 7898 25832
rect 8021 25823 8079 25829
rect 8021 25820 8033 25823
rect 7892 25792 8033 25820
rect 7892 25780 7898 25792
rect 8021 25789 8033 25792
rect 8067 25789 8079 25823
rect 8754 25820 8760 25832
rect 8021 25783 8079 25789
rect 8496 25792 8760 25820
rect 3326 25712 3332 25764
rect 3384 25752 3390 25764
rect 3421 25755 3479 25761
rect 3421 25752 3433 25755
rect 3384 25724 3433 25752
rect 3384 25712 3390 25724
rect 3421 25721 3433 25724
rect 3467 25721 3479 25755
rect 3620 25752 3648 25780
rect 4617 25755 4675 25761
rect 4617 25752 4629 25755
rect 3620 25724 4629 25752
rect 3421 25715 3479 25721
rect 4617 25721 4629 25724
rect 4663 25721 4675 25755
rect 4617 25715 4675 25721
rect 4246 25644 4252 25696
rect 4304 25644 4310 25696
rect 5442 25644 5448 25696
rect 5500 25684 5506 25696
rect 8496 25684 8524 25792
rect 8754 25780 8760 25792
rect 8812 25820 8818 25832
rect 9677 25823 9735 25829
rect 9677 25820 9689 25823
rect 8812 25792 9689 25820
rect 8812 25780 8818 25792
rect 9677 25789 9689 25792
rect 9723 25789 9735 25823
rect 9677 25783 9735 25789
rect 9769 25823 9827 25829
rect 9769 25789 9781 25823
rect 9815 25789 9827 25823
rect 9769 25783 9827 25789
rect 8570 25712 8576 25764
rect 8628 25752 8634 25764
rect 9582 25752 9588 25764
rect 8628 25724 9588 25752
rect 8628 25712 8634 25724
rect 9582 25712 9588 25724
rect 9640 25752 9646 25764
rect 9784 25752 9812 25783
rect 9858 25780 9864 25832
rect 9916 25820 9922 25832
rect 10965 25823 11023 25829
rect 10965 25820 10977 25823
rect 9916 25792 10977 25820
rect 9916 25780 9922 25792
rect 10965 25789 10977 25792
rect 11011 25789 11023 25823
rect 10965 25783 11023 25789
rect 11790 25780 11796 25832
rect 11848 25820 11854 25832
rect 11977 25823 12035 25829
rect 11977 25820 11989 25823
rect 11848 25792 11989 25820
rect 11848 25780 11854 25792
rect 11977 25789 11989 25792
rect 12023 25789 12035 25823
rect 11977 25783 12035 25789
rect 12989 25823 13047 25829
rect 12989 25789 13001 25823
rect 13035 25820 13047 25823
rect 14366 25820 14372 25832
rect 13035 25792 14372 25820
rect 13035 25789 13047 25792
rect 12989 25783 13047 25789
rect 14366 25780 14372 25792
rect 14424 25780 14430 25832
rect 14458 25780 14464 25832
rect 14516 25780 14522 25832
rect 9640 25724 9812 25752
rect 9640 25712 9646 25724
rect 8849 25687 8907 25693
rect 8849 25684 8861 25687
rect 5500 25656 8861 25684
rect 5500 25644 5506 25656
rect 8849 25653 8861 25656
rect 8895 25653 8907 25687
rect 8849 25647 8907 25653
rect 10413 25687 10471 25693
rect 10413 25653 10425 25687
rect 10459 25684 10471 25687
rect 12342 25684 12348 25696
rect 10459 25656 12348 25684
rect 10459 25653 10471 25656
rect 10413 25647 10471 25653
rect 12342 25644 12348 25656
rect 12400 25644 12406 25696
rect 15102 25644 15108 25696
rect 15160 25684 15166 25696
rect 15381 25687 15439 25693
rect 15381 25684 15393 25687
rect 15160 25656 15393 25684
rect 15160 25644 15166 25656
rect 15381 25653 15393 25656
rect 15427 25653 15439 25687
rect 15764 25684 15792 25851
rect 16022 25780 16028 25832
rect 16080 25780 16086 25832
rect 17862 25780 17868 25832
rect 17920 25780 17926 25832
rect 20548 25829 20576 25860
rect 22186 25848 22192 25860
rect 22244 25848 22250 25900
rect 22278 25848 22284 25900
rect 22336 25888 22342 25900
rect 22373 25891 22431 25897
rect 22373 25888 22385 25891
rect 22336 25860 22385 25888
rect 22336 25848 22342 25860
rect 22373 25857 22385 25860
rect 22419 25888 22431 25891
rect 23382 25888 23388 25900
rect 22419 25860 23388 25888
rect 22419 25857 22431 25860
rect 22373 25851 22431 25857
rect 23382 25848 23388 25860
rect 23440 25848 23446 25900
rect 23842 25848 23848 25900
rect 23900 25888 23906 25900
rect 23937 25891 23995 25897
rect 23937 25888 23949 25891
rect 23900 25860 23949 25888
rect 23900 25848 23906 25860
rect 23937 25857 23949 25860
rect 23983 25857 23995 25891
rect 23937 25851 23995 25857
rect 20533 25823 20591 25829
rect 20533 25789 20545 25823
rect 20579 25789 20591 25823
rect 20533 25783 20591 25789
rect 21266 25780 21272 25832
rect 21324 25780 21330 25832
rect 22557 25823 22615 25829
rect 22557 25789 22569 25823
rect 22603 25789 22615 25823
rect 22557 25783 22615 25789
rect 19889 25755 19947 25761
rect 19889 25752 19901 25755
rect 18892 25724 19901 25752
rect 18892 25696 18920 25724
rect 19889 25721 19901 25724
rect 19935 25721 19947 25755
rect 19889 25715 19947 25721
rect 22278 25712 22284 25764
rect 22336 25752 22342 25764
rect 22572 25752 22600 25783
rect 25130 25780 25136 25832
rect 25188 25780 25194 25832
rect 22336 25724 22600 25752
rect 23477 25755 23535 25761
rect 22336 25712 22342 25724
rect 23477 25721 23489 25755
rect 23523 25752 23535 25755
rect 24394 25752 24400 25764
rect 23523 25724 24400 25752
rect 23523 25721 23535 25724
rect 23477 25715 23535 25721
rect 24394 25712 24400 25724
rect 24452 25712 24458 25764
rect 18414 25684 18420 25696
rect 15764 25656 18420 25684
rect 15381 25647 15439 25653
rect 18414 25644 18420 25656
rect 18472 25644 18478 25696
rect 18874 25644 18880 25696
rect 18932 25644 18938 25696
rect 21358 25644 21364 25696
rect 21416 25684 21422 25696
rect 22005 25687 22063 25693
rect 22005 25684 22017 25687
rect 21416 25656 22017 25684
rect 21416 25644 21422 25656
rect 22005 25653 22017 25656
rect 22051 25653 22063 25687
rect 22005 25647 22063 25653
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 11425 25483 11483 25489
rect 11425 25449 11437 25483
rect 11471 25480 11483 25483
rect 14182 25480 14188 25492
rect 11471 25452 14188 25480
rect 11471 25449 11483 25452
rect 11425 25443 11483 25449
rect 14182 25440 14188 25452
rect 14240 25440 14246 25492
rect 14737 25483 14795 25489
rect 14737 25449 14749 25483
rect 14783 25480 14795 25483
rect 16758 25480 16764 25492
rect 14783 25452 16764 25480
rect 14783 25449 14795 25452
rect 14737 25443 14795 25449
rect 16758 25440 16764 25452
rect 16816 25440 16822 25492
rect 17586 25440 17592 25492
rect 17644 25480 17650 25492
rect 17770 25480 17776 25492
rect 17644 25452 17776 25480
rect 17644 25440 17650 25452
rect 17770 25440 17776 25452
rect 17828 25480 17834 25492
rect 17957 25483 18015 25489
rect 17957 25480 17969 25483
rect 17828 25452 17969 25480
rect 17828 25440 17834 25452
rect 17957 25449 17969 25452
rect 18003 25449 18015 25483
rect 17957 25443 18015 25449
rect 22370 25440 22376 25492
rect 22428 25480 22434 25492
rect 23109 25483 23167 25489
rect 23109 25480 23121 25483
rect 22428 25452 23121 25480
rect 22428 25440 22434 25452
rect 23109 25449 23121 25452
rect 23155 25449 23167 25483
rect 23109 25443 23167 25449
rect 23382 25440 23388 25492
rect 23440 25440 23446 25492
rect 24854 25440 24860 25492
rect 24912 25480 24918 25492
rect 25038 25480 25044 25492
rect 24912 25452 25044 25480
rect 24912 25440 24918 25452
rect 25038 25440 25044 25452
rect 25096 25480 25102 25492
rect 25133 25483 25191 25489
rect 25133 25480 25145 25483
rect 25096 25452 25145 25480
rect 25096 25440 25102 25452
rect 25133 25449 25145 25452
rect 25179 25449 25191 25483
rect 25133 25443 25191 25449
rect 25498 25440 25504 25492
rect 25556 25440 25562 25492
rect 14458 25412 14464 25424
rect 12406 25384 14464 25412
rect 6825 25347 6883 25353
rect 6825 25313 6837 25347
rect 6871 25344 6883 25347
rect 7650 25344 7656 25356
rect 6871 25316 7656 25344
rect 6871 25313 6883 25316
rect 6825 25307 6883 25313
rect 7650 25304 7656 25316
rect 7708 25304 7714 25356
rect 9398 25304 9404 25356
rect 9456 25304 9462 25356
rect 9674 25304 9680 25356
rect 9732 25344 9738 25356
rect 10597 25347 10655 25353
rect 10597 25344 10609 25347
rect 9732 25316 10609 25344
rect 9732 25304 9738 25316
rect 10597 25313 10609 25316
rect 10643 25313 10655 25347
rect 10597 25307 10655 25313
rect 11422 25304 11428 25356
rect 11480 25344 11486 25356
rect 11977 25347 12035 25353
rect 11977 25344 11989 25347
rect 11480 25316 11989 25344
rect 11480 25304 11486 25316
rect 11977 25313 11989 25316
rect 12023 25344 12035 25347
rect 12406 25344 12434 25384
rect 14458 25372 14464 25384
rect 14516 25372 14522 25424
rect 22097 25415 22155 25421
rect 15304 25384 16068 25412
rect 12023 25316 12434 25344
rect 12023 25313 12035 25316
rect 11977 25307 12035 25313
rect 12802 25304 12808 25356
rect 12860 25344 12866 25356
rect 13173 25347 13231 25353
rect 13173 25344 13185 25347
rect 12860 25316 13185 25344
rect 12860 25304 12866 25316
rect 13173 25313 13185 25316
rect 13219 25313 13231 25347
rect 13173 25307 13231 25313
rect 13814 25304 13820 25356
rect 13872 25344 13878 25356
rect 14182 25344 14188 25356
rect 13872 25316 14188 25344
rect 13872 25304 13878 25316
rect 14182 25304 14188 25316
rect 14240 25304 14246 25356
rect 15304 25353 15332 25384
rect 15289 25347 15347 25353
rect 15289 25313 15301 25347
rect 15335 25313 15347 25347
rect 15289 25307 15347 25313
rect 15378 25304 15384 25356
rect 15436 25344 15442 25356
rect 15933 25347 15991 25353
rect 15933 25344 15945 25347
rect 15436 25316 15945 25344
rect 15436 25304 15442 25316
rect 15933 25313 15945 25316
rect 15979 25313 15991 25347
rect 16040 25344 16068 25384
rect 22097 25381 22109 25415
rect 22143 25412 22155 25415
rect 24946 25412 24952 25424
rect 22143 25384 24952 25412
rect 22143 25381 22155 25384
rect 22097 25375 22155 25381
rect 24946 25372 24952 25384
rect 25004 25372 25010 25424
rect 16209 25347 16267 25353
rect 16209 25344 16221 25347
rect 16040 25316 16221 25344
rect 15933 25307 15991 25313
rect 16209 25313 16221 25316
rect 16255 25344 16267 25347
rect 16666 25344 16672 25356
rect 16255 25316 16672 25344
rect 16255 25313 16267 25316
rect 16209 25307 16267 25313
rect 16666 25304 16672 25316
rect 16724 25304 16730 25356
rect 19058 25304 19064 25356
rect 19116 25344 19122 25356
rect 19889 25347 19947 25353
rect 19889 25344 19901 25347
rect 19116 25316 19901 25344
rect 19116 25304 19122 25316
rect 19889 25313 19901 25316
rect 19935 25313 19947 25347
rect 19889 25307 19947 25313
rect 20070 25304 20076 25356
rect 20128 25304 20134 25356
rect 22646 25304 22652 25356
rect 22704 25304 22710 25356
rect 4062 25285 4068 25288
rect 4040 25279 4068 25285
rect 4040 25245 4052 25279
rect 4040 25239 4068 25245
rect 4062 25236 4068 25239
rect 4120 25236 4126 25288
rect 8386 25236 8392 25288
rect 8444 25276 8450 25288
rect 10413 25279 10471 25285
rect 10413 25276 10425 25279
rect 8444 25248 10425 25276
rect 8444 25236 8450 25248
rect 10413 25245 10425 25248
rect 10459 25245 10471 25279
rect 10413 25239 10471 25245
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25276 10563 25279
rect 10778 25276 10784 25288
rect 10551 25248 10784 25276
rect 10551 25245 10563 25248
rect 10505 25239 10563 25245
rect 10778 25236 10784 25248
rect 10836 25236 10842 25288
rect 11790 25236 11796 25288
rect 11848 25236 11854 25288
rect 12618 25236 12624 25288
rect 12676 25276 12682 25288
rect 13081 25279 13139 25285
rect 13081 25276 13093 25279
rect 12676 25248 13093 25276
rect 12676 25236 12682 25248
rect 13081 25245 13093 25248
rect 13127 25245 13139 25279
rect 13081 25239 13139 25245
rect 19426 25236 19432 25288
rect 19484 25276 19490 25288
rect 19797 25279 19855 25285
rect 19797 25276 19809 25279
rect 19484 25248 19809 25276
rect 19484 25236 19490 25248
rect 19797 25245 19809 25248
rect 19843 25245 19855 25279
rect 19797 25239 19855 25245
rect 21266 25236 21272 25288
rect 21324 25276 21330 25288
rect 22465 25279 22523 25285
rect 22465 25276 22477 25279
rect 21324 25248 22477 25276
rect 21324 25236 21330 25248
rect 22465 25245 22477 25248
rect 22511 25245 22523 25279
rect 22465 25239 22523 25245
rect 23845 25279 23903 25285
rect 23845 25245 23857 25279
rect 23891 25276 23903 25279
rect 24026 25276 24032 25288
rect 23891 25248 24032 25276
rect 23891 25245 23903 25248
rect 23845 25239 23903 25245
rect 24026 25236 24032 25248
rect 24084 25236 24090 25288
rect 24302 25236 24308 25288
rect 24360 25276 24366 25288
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 24360 25248 24685 25276
rect 24360 25236 24366 25248
rect 24673 25245 24685 25248
rect 24719 25245 24731 25279
rect 24673 25239 24731 25245
rect 7098 25168 7104 25220
rect 7156 25168 7162 25220
rect 8941 25211 8999 25217
rect 8941 25208 8953 25211
rect 8326 25180 8953 25208
rect 8941 25177 8953 25180
rect 8987 25208 8999 25211
rect 9766 25208 9772 25220
rect 8987 25180 9772 25208
rect 8987 25177 8999 25180
rect 8941 25171 8999 25177
rect 9766 25168 9772 25180
rect 9824 25168 9830 25220
rect 13446 25208 13452 25220
rect 10060 25180 13452 25208
rect 3970 25100 3976 25152
rect 4028 25140 4034 25152
rect 4111 25143 4169 25149
rect 4111 25140 4123 25143
rect 4028 25112 4123 25140
rect 4028 25100 4034 25112
rect 4111 25109 4123 25112
rect 4157 25109 4169 25143
rect 4111 25103 4169 25109
rect 8570 25100 8576 25152
rect 8628 25100 8634 25152
rect 10060 25149 10088 25180
rect 13446 25168 13452 25180
rect 13504 25168 13510 25220
rect 14642 25168 14648 25220
rect 14700 25208 14706 25220
rect 14700 25180 16698 25208
rect 14700 25168 14706 25180
rect 22094 25168 22100 25220
rect 22152 25208 22158 25220
rect 22557 25211 22615 25217
rect 22557 25208 22569 25211
rect 22152 25180 22569 25208
rect 22152 25168 22158 25180
rect 22557 25177 22569 25180
rect 22603 25177 22615 25211
rect 22557 25171 22615 25177
rect 24857 25211 24915 25217
rect 24857 25177 24869 25211
rect 24903 25208 24915 25211
rect 25038 25208 25044 25220
rect 24903 25180 25044 25208
rect 24903 25177 24915 25180
rect 24857 25171 24915 25177
rect 25038 25168 25044 25180
rect 25096 25168 25102 25220
rect 10045 25143 10103 25149
rect 10045 25109 10057 25143
rect 10091 25109 10103 25143
rect 10045 25103 10103 25109
rect 11146 25100 11152 25152
rect 11204 25140 11210 25152
rect 11885 25143 11943 25149
rect 11885 25140 11897 25143
rect 11204 25112 11897 25140
rect 11204 25100 11210 25112
rect 11885 25109 11897 25112
rect 11931 25140 11943 25143
rect 11974 25140 11980 25152
rect 11931 25112 11980 25140
rect 11931 25109 11943 25112
rect 11885 25103 11943 25109
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 12618 25100 12624 25152
rect 12676 25100 12682 25152
rect 12802 25100 12808 25152
rect 12860 25140 12866 25152
rect 12989 25143 13047 25149
rect 12989 25140 13001 25143
rect 12860 25112 13001 25140
rect 12860 25100 12866 25112
rect 12989 25109 13001 25112
rect 13035 25109 13047 25143
rect 12989 25103 13047 25109
rect 14918 25100 14924 25152
rect 14976 25140 14982 25152
rect 15105 25143 15163 25149
rect 15105 25140 15117 25143
rect 14976 25112 15117 25140
rect 14976 25100 14982 25112
rect 15105 25109 15117 25112
rect 15151 25109 15163 25143
rect 15105 25103 15163 25109
rect 15197 25143 15255 25149
rect 15197 25109 15209 25143
rect 15243 25140 15255 25143
rect 16850 25140 16856 25152
rect 15243 25112 16856 25140
rect 15243 25109 15255 25112
rect 15197 25103 15255 25109
rect 16850 25100 16856 25112
rect 16908 25100 16914 25152
rect 17034 25100 17040 25152
rect 17092 25140 17098 25152
rect 17681 25143 17739 25149
rect 17681 25140 17693 25143
rect 17092 25112 17693 25140
rect 17092 25100 17098 25112
rect 17681 25109 17693 25112
rect 17727 25140 17739 25143
rect 17862 25140 17868 25152
rect 17727 25112 17868 25140
rect 17727 25109 17739 25112
rect 17681 25103 17739 25109
rect 17862 25100 17868 25112
rect 17920 25100 17926 25152
rect 18233 25143 18291 25149
rect 18233 25109 18245 25143
rect 18279 25140 18291 25143
rect 18322 25140 18328 25152
rect 18279 25112 18328 25140
rect 18279 25109 18291 25112
rect 18233 25103 18291 25109
rect 18322 25100 18328 25112
rect 18380 25100 18386 25152
rect 19429 25143 19487 25149
rect 19429 25109 19441 25143
rect 19475 25140 19487 25143
rect 19518 25140 19524 25152
rect 19475 25112 19524 25140
rect 19475 25109 19487 25112
rect 19429 25103 19487 25109
rect 19518 25100 19524 25112
rect 19576 25100 19582 25152
rect 23934 25100 23940 25152
rect 23992 25100 23998 25152
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 4246 24896 4252 24948
rect 4304 24936 4310 24948
rect 5445 24939 5503 24945
rect 5445 24936 5457 24939
rect 4304 24908 5457 24936
rect 4304 24896 4310 24908
rect 5445 24905 5457 24908
rect 5491 24905 5503 24939
rect 5445 24899 5503 24905
rect 7834 24896 7840 24948
rect 7892 24936 7898 24948
rect 8021 24939 8079 24945
rect 8021 24936 8033 24939
rect 7892 24908 8033 24936
rect 7892 24896 7898 24908
rect 8021 24905 8033 24908
rect 8067 24905 8079 24939
rect 8021 24899 8079 24905
rect 9490 24896 9496 24948
rect 9548 24936 9554 24948
rect 11146 24936 11152 24948
rect 9548 24908 11152 24936
rect 9548 24896 9554 24908
rect 11146 24896 11152 24908
rect 11204 24896 11210 24948
rect 12618 24896 12624 24948
rect 12676 24936 12682 24948
rect 15197 24939 15255 24945
rect 15197 24936 15209 24939
rect 12676 24908 15209 24936
rect 12676 24896 12682 24908
rect 15197 24905 15209 24908
rect 15243 24905 15255 24939
rect 15197 24899 15255 24905
rect 16850 24896 16856 24948
rect 16908 24896 16914 24948
rect 7098 24828 7104 24880
rect 7156 24868 7162 24880
rect 9217 24871 9275 24877
rect 7156 24840 8340 24868
rect 7156 24828 7162 24840
rect 7377 24803 7435 24809
rect 5106 24772 6132 24800
rect 3697 24735 3755 24741
rect 3697 24701 3709 24735
rect 3743 24701 3755 24735
rect 3697 24695 3755 24701
rect 3973 24735 4031 24741
rect 3973 24701 3985 24735
rect 4019 24732 4031 24735
rect 5994 24732 6000 24744
rect 4019 24704 6000 24732
rect 4019 24701 4031 24704
rect 3973 24695 4031 24701
rect 3712 24596 3740 24695
rect 5994 24692 6000 24704
rect 6052 24692 6058 24744
rect 3970 24596 3976 24608
rect 3712 24568 3976 24596
rect 3970 24556 3976 24568
rect 4028 24556 4034 24608
rect 5813 24599 5871 24605
rect 5813 24565 5825 24599
rect 5859 24596 5871 24599
rect 6104 24596 6132 24772
rect 7377 24769 7389 24803
rect 7423 24800 7435 24803
rect 7558 24800 7564 24812
rect 7423 24772 7564 24800
rect 7423 24769 7435 24772
rect 7377 24763 7435 24769
rect 7558 24760 7564 24772
rect 7616 24760 7622 24812
rect 7742 24760 7748 24812
rect 7800 24800 7806 24812
rect 8312 24800 8340 24840
rect 9217 24837 9229 24871
rect 9263 24868 9275 24871
rect 12069 24871 12127 24877
rect 9263 24840 10088 24868
rect 9263 24837 9275 24840
rect 9217 24831 9275 24837
rect 10060 24809 10088 24840
rect 12069 24837 12081 24871
rect 12115 24868 12127 24871
rect 12986 24868 12992 24880
rect 12115 24840 12992 24868
rect 12115 24837 12127 24840
rect 12069 24831 12127 24837
rect 12986 24828 12992 24840
rect 13044 24828 13050 24880
rect 17218 24828 17224 24880
rect 17276 24828 17282 24880
rect 18322 24868 18328 24880
rect 17880 24840 18328 24868
rect 10045 24803 10103 24809
rect 7800 24772 8248 24800
rect 8312 24772 9444 24800
rect 7800 24760 7806 24772
rect 7576 24732 7604 24760
rect 8110 24732 8116 24744
rect 7576 24704 8116 24732
rect 8110 24692 8116 24704
rect 8168 24692 8174 24744
rect 8220 24741 8248 24772
rect 8205 24735 8263 24741
rect 8205 24701 8217 24735
rect 8251 24701 8263 24735
rect 8205 24695 8263 24701
rect 9306 24692 9312 24744
rect 9364 24692 9370 24744
rect 9416 24741 9444 24772
rect 10045 24769 10057 24803
rect 10091 24769 10103 24803
rect 10045 24763 10103 24769
rect 12161 24803 12219 24809
rect 12161 24769 12173 24803
rect 12207 24800 12219 24803
rect 12434 24800 12440 24812
rect 12207 24772 12440 24800
rect 12207 24769 12219 24772
rect 12161 24763 12219 24769
rect 12434 24760 12440 24772
rect 12492 24760 12498 24812
rect 12618 24760 12624 24812
rect 12676 24800 12682 24812
rect 13173 24803 13231 24809
rect 13173 24800 13185 24803
rect 12676 24772 13185 24800
rect 12676 24760 12682 24772
rect 13173 24769 13185 24772
rect 13219 24800 13231 24803
rect 13262 24800 13268 24812
rect 13219 24772 13268 24800
rect 13219 24769 13231 24772
rect 13173 24763 13231 24769
rect 13262 24760 13268 24772
rect 13320 24760 13326 24812
rect 13814 24760 13820 24812
rect 13872 24760 13878 24812
rect 14642 24800 14648 24812
rect 14108 24772 14648 24800
rect 9401 24735 9459 24741
rect 9401 24701 9413 24735
rect 9447 24701 9459 24735
rect 9401 24695 9459 24701
rect 9674 24692 9680 24744
rect 9732 24732 9738 24744
rect 12253 24735 12311 24741
rect 12253 24732 12265 24735
rect 9732 24704 12265 24732
rect 9732 24692 9738 24704
rect 12253 24701 12265 24704
rect 12299 24701 12311 24735
rect 12526 24732 12532 24744
rect 12253 24695 12311 24701
rect 12406 24704 12532 24732
rect 7653 24667 7711 24673
rect 7653 24633 7665 24667
rect 7699 24664 7711 24667
rect 8386 24664 8392 24676
rect 7699 24636 8392 24664
rect 7699 24633 7711 24636
rect 7653 24627 7711 24633
rect 8386 24624 8392 24636
rect 8444 24624 8450 24676
rect 11701 24667 11759 24673
rect 11701 24664 11713 24667
rect 8496 24636 11713 24664
rect 6914 24596 6920 24608
rect 5859 24568 6920 24596
rect 5859 24565 5871 24568
rect 5813 24559 5871 24565
rect 6914 24556 6920 24568
rect 6972 24556 6978 24608
rect 7466 24556 7472 24608
rect 7524 24596 7530 24608
rect 8496 24596 8524 24636
rect 11701 24633 11713 24636
rect 11747 24633 11759 24667
rect 11701 24627 11759 24633
rect 7524 24568 8524 24596
rect 8849 24599 8907 24605
rect 7524 24556 7530 24568
rect 8849 24565 8861 24599
rect 8895 24596 8907 24599
rect 11146 24596 11152 24608
rect 8895 24568 11152 24596
rect 8895 24565 8907 24568
rect 8849 24559 8907 24565
rect 11146 24556 11152 24568
rect 11204 24556 11210 24608
rect 12066 24556 12072 24608
rect 12124 24596 12130 24608
rect 12406 24596 12434 24704
rect 12526 24692 12532 24704
rect 12584 24692 12590 24744
rect 13280 24732 13308 24760
rect 14108 24741 14136 24772
rect 14642 24760 14648 24772
rect 14700 24760 14706 24812
rect 15010 24760 15016 24812
rect 15068 24800 15074 24812
rect 15289 24803 15347 24809
rect 15289 24800 15301 24803
rect 15068 24772 15301 24800
rect 15068 24760 15074 24772
rect 15289 24769 15301 24772
rect 15335 24769 15347 24803
rect 15289 24763 15347 24769
rect 16850 24760 16856 24812
rect 16908 24800 16914 24812
rect 17236 24800 17264 24828
rect 17880 24812 17908 24840
rect 18322 24828 18328 24840
rect 18380 24868 18386 24880
rect 18417 24871 18475 24877
rect 18417 24868 18429 24871
rect 18380 24840 18429 24868
rect 18380 24828 18386 24840
rect 18417 24837 18429 24840
rect 18463 24837 18475 24871
rect 18417 24831 18475 24837
rect 18506 24828 18512 24880
rect 18564 24868 18570 24880
rect 18564 24840 19932 24868
rect 18564 24828 18570 24840
rect 19904 24812 19932 24840
rect 22646 24828 22652 24880
rect 22704 24868 22710 24880
rect 23201 24871 23259 24877
rect 23201 24868 23213 24871
rect 22704 24840 23213 24868
rect 22704 24828 22710 24840
rect 23201 24837 23213 24840
rect 23247 24837 23259 24871
rect 23201 24831 23259 24837
rect 16908 24772 17264 24800
rect 17313 24803 17371 24809
rect 16908 24760 16914 24772
rect 17313 24769 17325 24803
rect 17359 24800 17371 24803
rect 17678 24800 17684 24812
rect 17359 24772 17448 24800
rect 17359 24769 17371 24772
rect 17313 24763 17371 24769
rect 13909 24735 13967 24741
rect 13909 24732 13921 24735
rect 13280 24704 13921 24732
rect 13909 24701 13921 24704
rect 13955 24701 13967 24735
rect 13909 24695 13967 24701
rect 14093 24735 14151 24741
rect 14093 24701 14105 24735
rect 14139 24701 14151 24735
rect 14093 24695 14151 24701
rect 14366 24692 14372 24744
rect 14424 24732 14430 24744
rect 15381 24735 15439 24741
rect 15381 24732 15393 24735
rect 14424 24704 15393 24732
rect 14424 24692 14430 24704
rect 15381 24701 15393 24704
rect 15427 24701 15439 24735
rect 15381 24695 15439 24701
rect 13449 24667 13507 24673
rect 13449 24633 13461 24667
rect 13495 24664 13507 24667
rect 14918 24664 14924 24676
rect 13495 24636 14924 24664
rect 13495 24633 13507 24636
rect 13449 24627 13507 24633
rect 14918 24624 14924 24636
rect 14976 24624 14982 24676
rect 17420 24664 17448 24772
rect 17512 24772 17684 24800
rect 17512 24741 17540 24772
rect 17678 24760 17684 24772
rect 17736 24760 17742 24812
rect 17862 24760 17868 24812
rect 17920 24760 17926 24812
rect 19886 24760 19892 24812
rect 19944 24800 19950 24812
rect 20625 24803 20683 24809
rect 20625 24800 20637 24803
rect 19944 24772 20637 24800
rect 19944 24760 19950 24772
rect 20625 24769 20637 24772
rect 20671 24769 20683 24803
rect 20625 24763 20683 24769
rect 20732 24772 20944 24800
rect 17497 24735 17555 24741
rect 17497 24701 17509 24735
rect 17543 24701 17555 24735
rect 17497 24695 17555 24701
rect 17586 24692 17592 24744
rect 17644 24732 17650 24744
rect 18509 24735 18567 24741
rect 18509 24732 18521 24735
rect 17644 24704 18521 24732
rect 17644 24692 17650 24704
rect 18509 24701 18521 24704
rect 18555 24701 18567 24735
rect 18509 24695 18567 24701
rect 18601 24735 18659 24741
rect 18601 24701 18613 24735
rect 18647 24732 18659 24735
rect 18782 24732 18788 24744
rect 18647 24704 18788 24732
rect 18647 24701 18659 24704
rect 18601 24695 18659 24701
rect 18782 24692 18788 24704
rect 18840 24692 18846 24744
rect 19242 24692 19248 24744
rect 19300 24732 19306 24744
rect 20732 24741 20760 24772
rect 20717 24735 20775 24741
rect 20717 24732 20729 24735
rect 19300 24704 20729 24732
rect 19300 24692 19306 24704
rect 20717 24701 20729 24704
rect 20763 24701 20775 24735
rect 20717 24695 20775 24701
rect 20809 24735 20867 24741
rect 20809 24701 20821 24735
rect 20855 24701 20867 24735
rect 20916 24732 20944 24772
rect 22002 24760 22008 24812
rect 22060 24800 22066 24812
rect 22094 24800 22100 24812
rect 22060 24772 22100 24800
rect 22060 24760 22066 24772
rect 22094 24760 22100 24772
rect 22152 24760 22158 24812
rect 24302 24760 24308 24812
rect 24360 24800 24366 24812
rect 24854 24800 24860 24812
rect 24360 24772 24860 24800
rect 24360 24760 24366 24772
rect 24854 24760 24860 24772
rect 24912 24760 24918 24812
rect 25317 24803 25375 24809
rect 25317 24769 25329 24803
rect 25363 24800 25375 24803
rect 25498 24800 25504 24812
rect 25363 24772 25504 24800
rect 25363 24769 25375 24772
rect 25317 24763 25375 24769
rect 25498 24760 25504 24772
rect 25556 24760 25562 24812
rect 22830 24732 22836 24744
rect 20916 24704 22836 24732
rect 20809 24695 20867 24701
rect 18690 24664 18696 24676
rect 16316 24636 17356 24664
rect 17420 24636 18696 24664
rect 12713 24599 12771 24605
rect 12713 24596 12725 24599
rect 12124 24568 12725 24596
rect 12124 24556 12130 24568
rect 12713 24565 12725 24568
rect 12759 24565 12771 24599
rect 12713 24559 12771 24565
rect 12986 24556 12992 24608
rect 13044 24596 13050 24608
rect 13722 24596 13728 24608
rect 13044 24568 13728 24596
rect 13044 24556 13050 24568
rect 13722 24556 13728 24568
rect 13780 24556 13786 24608
rect 14553 24599 14611 24605
rect 14553 24565 14565 24599
rect 14599 24596 14611 24599
rect 14642 24596 14648 24608
rect 14599 24568 14648 24596
rect 14599 24565 14611 24568
rect 14553 24559 14611 24565
rect 14642 24556 14648 24568
rect 14700 24556 14706 24608
rect 14829 24599 14887 24605
rect 14829 24565 14841 24599
rect 14875 24596 14887 24599
rect 16316 24596 16344 24636
rect 17328 24608 17356 24636
rect 18690 24624 18696 24636
rect 18748 24624 18754 24676
rect 20530 24624 20536 24676
rect 20588 24664 20594 24676
rect 20824 24664 20852 24695
rect 22830 24692 22836 24704
rect 22888 24692 22894 24744
rect 22925 24735 22983 24741
rect 22925 24701 22937 24735
rect 22971 24701 22983 24735
rect 22925 24695 22983 24701
rect 20588 24636 20852 24664
rect 20588 24624 20594 24636
rect 22094 24624 22100 24676
rect 22152 24664 22158 24676
rect 22940 24664 22968 24695
rect 24670 24692 24676 24744
rect 24728 24692 24734 24744
rect 22152 24636 22968 24664
rect 22152 24624 22158 24636
rect 14875 24568 16344 24596
rect 16485 24599 16543 24605
rect 14875 24565 14887 24568
rect 14829 24559 14887 24565
rect 16485 24565 16497 24599
rect 16531 24596 16543 24599
rect 16850 24596 16856 24608
rect 16531 24568 16856 24596
rect 16531 24565 16543 24568
rect 16485 24559 16543 24565
rect 16850 24556 16856 24568
rect 16908 24556 16914 24608
rect 17310 24556 17316 24608
rect 17368 24556 17374 24608
rect 18049 24599 18107 24605
rect 18049 24565 18061 24599
rect 18095 24596 18107 24599
rect 18506 24596 18512 24608
rect 18095 24568 18512 24596
rect 18095 24565 18107 24568
rect 18049 24559 18107 24565
rect 18506 24556 18512 24568
rect 18564 24556 18570 24608
rect 19886 24556 19892 24608
rect 19944 24556 19950 24608
rect 20257 24599 20315 24605
rect 20257 24565 20269 24599
rect 20303 24596 20315 24599
rect 24578 24596 24584 24608
rect 20303 24568 24584 24596
rect 20303 24565 20315 24568
rect 20257 24559 20315 24565
rect 24578 24556 24584 24568
rect 24636 24556 24642 24608
rect 24762 24556 24768 24608
rect 24820 24596 24826 24608
rect 25133 24599 25191 24605
rect 25133 24596 25145 24599
rect 24820 24568 25145 24596
rect 24820 24556 24826 24568
rect 25133 24565 25145 24568
rect 25179 24565 25191 24599
rect 25133 24559 25191 24565
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 3237 24395 3295 24401
rect 3237 24361 3249 24395
rect 3283 24361 3295 24395
rect 3237 24355 3295 24361
rect 3252 24324 3280 24355
rect 3418 24352 3424 24404
rect 3476 24352 3482 24404
rect 4430 24392 4436 24404
rect 3620 24364 4436 24392
rect 3620 24324 3648 24364
rect 4430 24352 4436 24364
rect 4488 24392 4494 24404
rect 5721 24395 5779 24401
rect 5721 24392 5733 24395
rect 4488 24364 5733 24392
rect 4488 24352 4494 24364
rect 5721 24361 5733 24364
rect 5767 24361 5779 24395
rect 5721 24355 5779 24361
rect 6178 24352 6184 24404
rect 6236 24352 6242 24404
rect 8754 24352 8760 24404
rect 8812 24392 8818 24404
rect 9306 24392 9312 24404
rect 8812 24364 9312 24392
rect 8812 24352 8818 24364
rect 9306 24352 9312 24364
rect 9364 24352 9370 24404
rect 10318 24352 10324 24404
rect 10376 24392 10382 24404
rect 10376 24364 12434 24392
rect 10376 24352 10382 24364
rect 3252 24296 3648 24324
rect 6362 24284 6368 24336
rect 6420 24284 6426 24336
rect 8570 24284 8576 24336
rect 8628 24324 8634 24336
rect 8628 24296 11376 24324
rect 8628 24284 8634 24296
rect 4246 24216 4252 24268
rect 4304 24216 4310 24268
rect 6380 24256 6408 24284
rect 9858 24256 9864 24268
rect 6380 24228 9864 24256
rect 9858 24216 9864 24228
rect 9916 24216 9922 24268
rect 10045 24259 10103 24265
rect 10045 24225 10057 24259
rect 10091 24256 10103 24259
rect 10410 24256 10416 24268
rect 10091 24228 10416 24256
rect 10091 24225 10103 24228
rect 10045 24219 10103 24225
rect 10410 24216 10416 24228
rect 10468 24216 10474 24268
rect 10505 24259 10563 24265
rect 10505 24225 10517 24259
rect 10551 24256 10563 24259
rect 11054 24256 11060 24268
rect 10551 24228 11060 24256
rect 10551 24225 10563 24228
rect 10505 24219 10563 24225
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2774 24188 2780 24200
rect 2271 24160 2780 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2774 24148 2780 24160
rect 2832 24148 2838 24200
rect 2961 24191 3019 24197
rect 2961 24157 2973 24191
rect 3007 24188 3019 24191
rect 3510 24188 3516 24200
rect 3007 24160 3516 24188
rect 3007 24157 3019 24160
rect 2961 24151 3019 24157
rect 2685 24123 2743 24129
rect 2685 24089 2697 24123
rect 2731 24120 2743 24123
rect 2976 24120 3004 24151
rect 3510 24148 3516 24160
rect 3568 24148 3574 24200
rect 3970 24148 3976 24200
rect 4028 24148 4034 24200
rect 6365 24191 6423 24197
rect 6365 24157 6377 24191
rect 6411 24188 6423 24191
rect 7098 24188 7104 24200
rect 6411 24160 7104 24188
rect 6411 24157 6423 24160
rect 6365 24151 6423 24157
rect 7098 24148 7104 24160
rect 7156 24148 7162 24200
rect 9876 24160 10088 24188
rect 2731 24092 3004 24120
rect 3528 24120 3556 24148
rect 4246 24120 4252 24132
rect 3528 24092 4252 24120
rect 2731 24089 2743 24092
rect 2685 24083 2743 24089
rect 4246 24080 4252 24092
rect 4304 24080 4310 24132
rect 9876 24129 9904 24160
rect 9861 24123 9919 24129
rect 5474 24092 6776 24120
rect 1854 24012 1860 24064
rect 1912 24052 1918 24064
rect 6748 24061 6776 24092
rect 9861 24089 9873 24123
rect 9907 24089 9919 24123
rect 10060 24120 10088 24160
rect 10612 24120 10640 24228
rect 11054 24216 11060 24228
rect 11112 24216 11118 24268
rect 11348 24265 11376 24296
rect 11333 24259 11391 24265
rect 11333 24225 11345 24259
rect 11379 24225 11391 24259
rect 12406 24256 12434 24364
rect 12526 24352 12532 24404
rect 12584 24392 12590 24404
rect 13354 24392 13360 24404
rect 12584 24364 13360 24392
rect 12584 24352 12590 24364
rect 13354 24352 13360 24364
rect 13412 24352 13418 24404
rect 13725 24395 13783 24401
rect 13725 24361 13737 24395
rect 13771 24392 13783 24395
rect 15194 24392 15200 24404
rect 13771 24364 15200 24392
rect 13771 24361 13783 24364
rect 13725 24355 13783 24361
rect 12529 24259 12587 24265
rect 12529 24256 12541 24259
rect 12406 24228 12541 24256
rect 11333 24219 11391 24225
rect 12529 24225 12541 24228
rect 12575 24225 12587 24259
rect 12529 24219 12587 24225
rect 12802 24216 12808 24268
rect 12860 24256 12866 24268
rect 13173 24259 13231 24265
rect 13173 24256 13185 24259
rect 12860 24228 13185 24256
rect 12860 24216 12866 24228
rect 13173 24225 13185 24228
rect 13219 24225 13231 24259
rect 13173 24219 13231 24225
rect 11146 24148 11152 24200
rect 11204 24148 11210 24200
rect 11241 24191 11299 24197
rect 11241 24157 11253 24191
rect 11287 24188 11299 24191
rect 13538 24188 13544 24200
rect 11287 24160 13544 24188
rect 11287 24157 11299 24160
rect 11241 24151 11299 24157
rect 13538 24148 13544 24160
rect 13596 24148 13602 24200
rect 10060 24092 10640 24120
rect 9861 24083 9919 24089
rect 11514 24080 11520 24132
rect 11572 24120 11578 24132
rect 11790 24120 11796 24132
rect 11572 24092 11796 24120
rect 11572 24080 11578 24092
rect 11790 24080 11796 24092
rect 11848 24120 11854 24132
rect 12437 24123 12495 24129
rect 12437 24120 12449 24123
rect 11848 24092 12449 24120
rect 11848 24080 11854 24092
rect 12437 24089 12449 24092
rect 12483 24089 12495 24123
rect 12437 24083 12495 24089
rect 2041 24055 2099 24061
rect 2041 24052 2053 24055
rect 1912 24024 2053 24052
rect 1912 24012 1918 24024
rect 2041 24021 2053 24024
rect 2087 24021 2099 24055
rect 2041 24015 2099 24021
rect 6733 24055 6791 24061
rect 6733 24021 6745 24055
rect 6779 24052 6791 24055
rect 6914 24052 6920 24064
rect 6779 24024 6920 24052
rect 6779 24021 6791 24024
rect 6733 24015 6791 24021
rect 6914 24012 6920 24024
rect 6972 24052 6978 24064
rect 7834 24052 7840 24064
rect 6972 24024 7840 24052
rect 6972 24012 6978 24024
rect 7834 24012 7840 24024
rect 7892 24052 7898 24064
rect 8478 24052 8484 24064
rect 7892 24024 8484 24052
rect 7892 24012 7898 24024
rect 8478 24012 8484 24024
rect 8536 24052 8542 24064
rect 9306 24052 9312 24064
rect 8536 24024 9312 24052
rect 8536 24012 8542 24024
rect 9306 24012 9312 24024
rect 9364 24012 9370 24064
rect 9398 24012 9404 24064
rect 9456 24012 9462 24064
rect 9766 24012 9772 24064
rect 9824 24012 9830 24064
rect 10778 24012 10784 24064
rect 10836 24012 10842 24064
rect 11974 24012 11980 24064
rect 12032 24012 12038 24064
rect 12345 24055 12403 24061
rect 12345 24021 12357 24055
rect 12391 24052 12403 24055
rect 13740 24052 13768 24355
rect 15194 24352 15200 24364
rect 15252 24392 15258 24404
rect 15654 24392 15660 24404
rect 15252 24364 15660 24392
rect 15252 24352 15258 24364
rect 15654 24352 15660 24364
rect 15712 24352 15718 24404
rect 17586 24352 17592 24404
rect 17644 24392 17650 24404
rect 21818 24392 21824 24404
rect 17644 24364 21824 24392
rect 17644 24352 17650 24364
rect 21818 24352 21824 24364
rect 21876 24352 21882 24404
rect 24670 24352 24676 24404
rect 24728 24392 24734 24404
rect 24728 24364 25176 24392
rect 24728 24352 24734 24364
rect 14642 24284 14648 24336
rect 14700 24324 14706 24336
rect 17678 24324 17684 24336
rect 14700 24296 17684 24324
rect 14700 24284 14706 24296
rect 17678 24284 17684 24296
rect 17736 24284 17742 24336
rect 18233 24327 18291 24333
rect 18233 24293 18245 24327
rect 18279 24324 18291 24327
rect 18690 24324 18696 24336
rect 18279 24296 18696 24324
rect 18279 24293 18291 24296
rect 18233 24287 18291 24293
rect 18690 24284 18696 24296
rect 18748 24284 18754 24336
rect 24762 24324 24768 24336
rect 22204 24296 24768 24324
rect 13814 24216 13820 24268
rect 13872 24256 13878 24268
rect 14277 24259 14335 24265
rect 14277 24256 14289 24259
rect 13872 24228 14289 24256
rect 13872 24216 13878 24228
rect 14277 24225 14289 24228
rect 14323 24225 14335 24259
rect 14277 24219 14335 24225
rect 16853 24259 16911 24265
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 16942 24256 16948 24268
rect 16899 24228 16948 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 17034 24216 17040 24268
rect 17092 24216 17098 24268
rect 19705 24259 19763 24265
rect 19705 24225 19717 24259
rect 19751 24256 19763 24259
rect 22094 24256 22100 24268
rect 19751 24228 22100 24256
rect 19751 24225 19763 24228
rect 19705 24219 19763 24225
rect 22094 24216 22100 24228
rect 22152 24216 22158 24268
rect 16758 24148 16764 24200
rect 16816 24148 16822 24200
rect 17773 24191 17831 24197
rect 17773 24157 17785 24191
rect 17819 24157 17831 24191
rect 17773 24151 17831 24157
rect 14550 24080 14556 24132
rect 14608 24120 14614 24132
rect 17788 24120 17816 24151
rect 21726 24148 21732 24200
rect 21784 24188 21790 24200
rect 22005 24191 22063 24197
rect 22005 24188 22017 24191
rect 21784 24160 22017 24188
rect 21784 24148 21790 24160
rect 22005 24157 22017 24160
rect 22051 24157 22063 24191
rect 22204 24188 22232 24296
rect 24762 24284 24768 24296
rect 24820 24284 24826 24336
rect 23845 24259 23903 24265
rect 23845 24225 23857 24259
rect 23891 24256 23903 24259
rect 24854 24256 24860 24268
rect 23891 24228 24860 24256
rect 23891 24225 23903 24228
rect 23845 24219 23903 24225
rect 24854 24216 24860 24228
rect 24912 24216 24918 24268
rect 25148 24265 25176 24364
rect 25133 24259 25191 24265
rect 25133 24225 25145 24259
rect 25179 24225 25191 24259
rect 25133 24219 25191 24225
rect 22005 24151 22063 24157
rect 22112 24160 22232 24188
rect 22833 24191 22891 24197
rect 14608 24092 17816 24120
rect 14608 24080 14614 24092
rect 18782 24080 18788 24132
rect 18840 24120 18846 24132
rect 19242 24120 19248 24132
rect 18840 24092 19248 24120
rect 18840 24080 18846 24092
rect 19242 24080 19248 24092
rect 19300 24120 19306 24132
rect 19981 24123 20039 24129
rect 19981 24120 19993 24123
rect 19300 24092 19993 24120
rect 19300 24080 19306 24092
rect 19981 24089 19993 24092
rect 20027 24089 20039 24123
rect 21634 24120 21640 24132
rect 21206 24092 21640 24120
rect 19981 24083 20039 24089
rect 21634 24080 21640 24092
rect 21692 24080 21698 24132
rect 21818 24080 21824 24132
rect 21876 24120 21882 24132
rect 22112 24120 22140 24160
rect 22833 24157 22845 24191
rect 22879 24188 22891 24191
rect 23290 24188 23296 24200
rect 22879 24160 23296 24188
rect 22879 24157 22891 24160
rect 22833 24151 22891 24157
rect 23290 24148 23296 24160
rect 23348 24148 23354 24200
rect 24946 24148 24952 24200
rect 25004 24148 25010 24200
rect 25041 24191 25099 24197
rect 25041 24157 25053 24191
rect 25087 24188 25099 24191
rect 25682 24188 25688 24200
rect 25087 24160 25688 24188
rect 25087 24157 25099 24160
rect 25041 24151 25099 24157
rect 25682 24148 25688 24160
rect 25740 24148 25746 24200
rect 21876 24092 22140 24120
rect 21876 24080 21882 24092
rect 22186 24080 22192 24132
rect 22244 24080 22250 24132
rect 12391 24024 13768 24052
rect 16393 24055 16451 24061
rect 12391 24021 12403 24024
rect 12345 24015 12403 24021
rect 16393 24021 16405 24055
rect 16439 24052 16451 24055
rect 17126 24052 17132 24064
rect 16439 24024 17132 24052
rect 16439 24021 16451 24024
rect 16393 24015 16451 24021
rect 17126 24012 17132 24024
rect 17184 24012 17190 24064
rect 17402 24012 17408 24064
rect 17460 24052 17466 24064
rect 17589 24055 17647 24061
rect 17589 24052 17601 24055
rect 17460 24024 17601 24052
rect 17460 24012 17466 24024
rect 17589 24021 17601 24024
rect 17635 24021 17647 24055
rect 17589 24015 17647 24021
rect 17678 24012 17684 24064
rect 17736 24052 17742 24064
rect 18141 24055 18199 24061
rect 18141 24052 18153 24055
rect 17736 24024 18153 24052
rect 17736 24012 17742 24024
rect 18141 24021 18153 24024
rect 18187 24052 18199 24055
rect 19426 24052 19432 24064
rect 18187 24024 19432 24052
rect 18187 24021 18199 24024
rect 18141 24015 18199 24021
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 20254 24012 20260 24064
rect 20312 24052 20318 24064
rect 21453 24055 21511 24061
rect 21453 24052 21465 24055
rect 20312 24024 21465 24052
rect 20312 24012 20318 24024
rect 21453 24021 21465 24024
rect 21499 24021 21511 24055
rect 21453 24015 21511 24021
rect 23566 24012 23572 24064
rect 23624 24052 23630 24064
rect 24581 24055 24639 24061
rect 24581 24052 24593 24055
rect 23624 24024 24593 24052
rect 23624 24012 23630 24024
rect 24581 24021 24593 24024
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 5994 23808 6000 23860
rect 6052 23808 6058 23860
rect 6822 23808 6828 23860
rect 6880 23848 6886 23860
rect 9401 23851 9459 23857
rect 9401 23848 9413 23851
rect 6880 23820 9413 23848
rect 6880 23808 6886 23820
rect 9401 23817 9413 23820
rect 9447 23848 9459 23851
rect 9674 23848 9680 23860
rect 9447 23820 9680 23848
rect 9447 23817 9459 23820
rect 9401 23811 9459 23817
rect 9674 23808 9680 23820
rect 9732 23808 9738 23860
rect 9766 23808 9772 23860
rect 9824 23848 9830 23860
rect 9861 23851 9919 23857
rect 9861 23848 9873 23851
rect 9824 23820 9873 23848
rect 9824 23808 9830 23820
rect 9861 23817 9873 23820
rect 9907 23817 9919 23851
rect 9861 23811 9919 23817
rect 10778 23808 10784 23860
rect 10836 23848 10842 23860
rect 14826 23848 14832 23860
rect 10836 23820 14832 23848
rect 10836 23808 10842 23820
rect 14826 23808 14832 23820
rect 14884 23808 14890 23860
rect 19242 23808 19248 23860
rect 19300 23848 19306 23860
rect 19300 23820 20484 23848
rect 19300 23808 19306 23820
rect 4154 23740 4160 23792
rect 4212 23780 4218 23792
rect 4430 23780 4436 23792
rect 4212 23752 4436 23780
rect 4212 23740 4218 23752
rect 4430 23740 4436 23752
rect 4488 23740 4494 23792
rect 6457 23783 6515 23789
rect 6457 23780 6469 23783
rect 5750 23752 6469 23780
rect 6457 23749 6469 23752
rect 6503 23780 6515 23783
rect 6914 23780 6920 23792
rect 6503 23752 6920 23780
rect 6503 23749 6515 23752
rect 6457 23743 6515 23749
rect 6914 23740 6920 23752
rect 6972 23740 6978 23792
rect 8478 23740 8484 23792
rect 8536 23740 8542 23792
rect 9306 23740 9312 23792
rect 9364 23780 9370 23792
rect 10321 23783 10379 23789
rect 10321 23780 10333 23783
rect 9364 23752 10333 23780
rect 9364 23740 9370 23752
rect 10321 23749 10333 23752
rect 10367 23749 10379 23783
rect 10321 23743 10379 23749
rect 11790 23740 11796 23792
rect 11848 23740 11854 23792
rect 11882 23740 11888 23792
rect 11940 23780 11946 23792
rect 17862 23780 17868 23792
rect 11940 23752 17868 23780
rect 11940 23740 11946 23752
rect 17862 23740 17868 23752
rect 17920 23740 17926 23792
rect 18966 23780 18972 23792
rect 17972 23752 18972 23780
rect 1762 23672 1768 23724
rect 1820 23672 1826 23724
rect 9858 23672 9864 23724
rect 9916 23712 9922 23724
rect 11808 23712 11836 23740
rect 9916 23684 11836 23712
rect 9916 23672 9922 23684
rect 12158 23672 12164 23724
rect 12216 23712 12222 23724
rect 12216 23684 13676 23712
rect 12216 23672 12222 23684
rect 1302 23604 1308 23656
rect 1360 23644 1366 23656
rect 2041 23647 2099 23653
rect 2041 23644 2053 23647
rect 1360 23616 2053 23644
rect 1360 23604 1366 23616
rect 2041 23613 2053 23616
rect 2087 23613 2099 23647
rect 2041 23607 2099 23613
rect 3970 23604 3976 23656
rect 4028 23644 4034 23656
rect 4249 23647 4307 23653
rect 4249 23644 4261 23647
rect 4028 23616 4261 23644
rect 4028 23604 4034 23616
rect 4249 23613 4261 23616
rect 4295 23613 4307 23647
rect 4249 23607 4307 23613
rect 4525 23647 4583 23653
rect 4525 23613 4537 23647
rect 4571 23644 4583 23647
rect 7558 23644 7564 23656
rect 4571 23616 7564 23644
rect 4571 23613 4583 23616
rect 4525 23607 4583 23613
rect 4264 23508 4292 23607
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 7650 23604 7656 23656
rect 7708 23604 7714 23656
rect 7929 23647 7987 23653
rect 7929 23613 7941 23647
rect 7975 23644 7987 23647
rect 8570 23644 8576 23656
rect 7975 23616 8576 23644
rect 7975 23613 7987 23616
rect 7929 23607 7987 23613
rect 8570 23604 8576 23616
rect 8628 23604 8634 23656
rect 10873 23647 10931 23653
rect 10873 23613 10885 23647
rect 10919 23644 10931 23647
rect 11698 23644 11704 23656
rect 10919 23616 11704 23644
rect 10919 23613 10931 23616
rect 10873 23607 10931 23613
rect 11698 23604 11704 23616
rect 11756 23604 11762 23656
rect 12437 23647 12495 23653
rect 12437 23613 12449 23647
rect 12483 23644 12495 23647
rect 12618 23644 12624 23656
rect 12483 23616 12624 23644
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 12618 23604 12624 23616
rect 12676 23604 12682 23656
rect 13648 23644 13676 23684
rect 13722 23672 13728 23724
rect 13780 23712 13786 23724
rect 17218 23712 17224 23724
rect 13780 23684 17224 23712
rect 13780 23672 13786 23684
rect 17218 23672 17224 23684
rect 17276 23672 17282 23724
rect 14366 23644 14372 23656
rect 13648 23616 14372 23644
rect 14366 23604 14372 23616
rect 14424 23644 14430 23656
rect 14918 23644 14924 23656
rect 14424 23616 14924 23644
rect 14424 23604 14430 23616
rect 14918 23604 14924 23616
rect 14976 23604 14982 23656
rect 17034 23604 17040 23656
rect 17092 23604 17098 23656
rect 5718 23508 5724 23520
rect 4264 23480 5724 23508
rect 5718 23468 5724 23480
rect 5776 23468 5782 23520
rect 7668 23508 7696 23604
rect 16482 23576 16488 23588
rect 11532 23548 16488 23576
rect 9950 23508 9956 23520
rect 7668 23480 9956 23508
rect 9950 23468 9956 23480
rect 10008 23468 10014 23520
rect 10962 23468 10968 23520
rect 11020 23508 11026 23520
rect 11532 23517 11560 23548
rect 16482 23536 16488 23548
rect 16540 23536 16546 23588
rect 11517 23511 11575 23517
rect 11517 23508 11529 23511
rect 11020 23480 11529 23508
rect 11020 23468 11026 23480
rect 11517 23477 11529 23480
rect 11563 23477 11575 23511
rect 11517 23471 11575 23477
rect 12158 23468 12164 23520
rect 12216 23468 12222 23520
rect 12434 23468 12440 23520
rect 12492 23508 12498 23520
rect 12529 23511 12587 23517
rect 12529 23508 12541 23511
rect 12492 23480 12541 23508
rect 12492 23468 12498 23480
rect 12529 23477 12541 23480
rect 12575 23508 12587 23511
rect 13722 23508 13728 23520
rect 12575 23480 13728 23508
rect 12575 23477 12587 23480
rect 12529 23471 12587 23477
rect 13722 23468 13728 23480
rect 13780 23468 13786 23520
rect 13906 23468 13912 23520
rect 13964 23508 13970 23520
rect 17972 23508 18000 23752
rect 18966 23740 18972 23752
rect 19024 23740 19030 23792
rect 19334 23740 19340 23792
rect 19392 23780 19398 23792
rect 19392 23752 19550 23780
rect 19392 23740 19398 23752
rect 20456 23712 20484 23820
rect 21634 23808 21640 23860
rect 21692 23808 21698 23860
rect 22830 23808 22836 23860
rect 22888 23848 22894 23860
rect 25133 23851 25191 23857
rect 25133 23848 25145 23851
rect 22888 23820 25145 23848
rect 22888 23808 22894 23820
rect 25133 23817 25145 23820
rect 25179 23817 25191 23851
rect 25133 23811 25191 23817
rect 20530 23740 20536 23792
rect 20588 23780 20594 23792
rect 23198 23780 23204 23792
rect 20588 23752 23204 23780
rect 20588 23740 20594 23752
rect 23198 23740 23204 23752
rect 23256 23740 23262 23792
rect 20456 23684 20944 23712
rect 18598 23604 18604 23656
rect 18656 23644 18662 23656
rect 18785 23647 18843 23653
rect 18785 23644 18797 23647
rect 18656 23616 18797 23644
rect 18656 23604 18662 23616
rect 18785 23613 18797 23616
rect 18831 23613 18843 23647
rect 18785 23607 18843 23613
rect 19058 23604 19064 23656
rect 19116 23604 19122 23656
rect 19426 23604 19432 23656
rect 19484 23644 19490 23656
rect 20809 23647 20867 23653
rect 20809 23644 20821 23647
rect 19484 23616 20821 23644
rect 19484 23604 19490 23616
rect 20809 23613 20821 23616
rect 20855 23613 20867 23647
rect 20916 23644 20944 23684
rect 22002 23672 22008 23724
rect 22060 23712 22066 23724
rect 22094 23712 22100 23724
rect 22060 23684 22100 23712
rect 22060 23672 22066 23684
rect 22094 23672 22100 23684
rect 22152 23712 22158 23724
rect 22152 23684 22232 23712
rect 22152 23672 22158 23684
rect 20916 23616 22094 23644
rect 20809 23607 20867 23613
rect 13964 23480 18000 23508
rect 13964 23468 13970 23480
rect 21082 23468 21088 23520
rect 21140 23468 21146 23520
rect 22066 23508 22094 23616
rect 22204 23576 22232 23684
rect 24302 23672 24308 23724
rect 24360 23672 24366 23724
rect 25314 23672 25320 23724
rect 25372 23672 25378 23724
rect 22925 23647 22983 23653
rect 22925 23613 22937 23647
rect 22971 23613 22983 23647
rect 22925 23607 22983 23613
rect 22940 23576 22968 23607
rect 23198 23604 23204 23656
rect 23256 23644 23262 23656
rect 23658 23644 23664 23656
rect 23256 23616 23664 23644
rect 23256 23604 23262 23616
rect 23658 23604 23664 23616
rect 23716 23604 23722 23656
rect 24486 23604 24492 23656
rect 24544 23644 24550 23656
rect 24673 23647 24731 23653
rect 24673 23644 24685 23647
rect 24544 23616 24685 23644
rect 24544 23604 24550 23616
rect 24673 23613 24685 23616
rect 24719 23613 24731 23647
rect 24673 23607 24731 23613
rect 22204 23548 22968 23576
rect 24210 23508 24216 23520
rect 22066 23480 24216 23508
rect 24210 23468 24216 23480
rect 24268 23468 24274 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 2038 23264 2044 23316
rect 2096 23264 2102 23316
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 3145 23307 3203 23313
rect 3145 23304 3157 23307
rect 2924 23276 3157 23304
rect 2924 23264 2930 23276
rect 3145 23273 3157 23276
rect 3191 23273 3203 23307
rect 3145 23267 3203 23273
rect 3878 23264 3884 23316
rect 3936 23304 3942 23316
rect 3936 23276 7144 23304
rect 3936 23264 3942 23276
rect 7116 23236 7144 23276
rect 7558 23264 7564 23316
rect 7616 23264 7622 23316
rect 12618 23304 12624 23316
rect 7668 23276 12624 23304
rect 7668 23236 7696 23276
rect 12618 23264 12624 23276
rect 12676 23304 12682 23316
rect 12802 23304 12808 23316
rect 12676 23276 12808 23304
rect 12676 23264 12682 23276
rect 12802 23264 12808 23276
rect 12860 23264 12866 23316
rect 14550 23264 14556 23316
rect 14608 23304 14614 23316
rect 16022 23304 16028 23316
rect 14608 23276 16028 23304
rect 14608 23264 14614 23276
rect 16022 23264 16028 23276
rect 16080 23264 16086 23316
rect 16390 23264 16396 23316
rect 16448 23304 16454 23316
rect 17770 23304 17776 23316
rect 16448 23276 17776 23304
rect 16448 23264 16454 23276
rect 17770 23264 17776 23276
rect 17828 23304 17834 23316
rect 18509 23307 18567 23313
rect 18509 23304 18521 23307
rect 17828 23276 18521 23304
rect 17828 23264 17834 23276
rect 18509 23273 18521 23276
rect 18555 23304 18567 23307
rect 19334 23304 19340 23316
rect 18555 23276 19340 23304
rect 18555 23273 18567 23276
rect 18509 23267 18567 23273
rect 19334 23264 19340 23276
rect 19392 23264 19398 23316
rect 20070 23264 20076 23316
rect 20128 23304 20134 23316
rect 20438 23304 20444 23316
rect 20128 23276 20444 23304
rect 20128 23264 20134 23276
rect 20438 23264 20444 23276
rect 20496 23304 20502 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 20496 23276 21189 23304
rect 20496 23264 20502 23276
rect 21177 23273 21189 23276
rect 21223 23273 21235 23307
rect 21177 23267 21235 23273
rect 7116 23208 7696 23236
rect 7834 23196 7840 23248
rect 7892 23196 7898 23248
rect 9766 23196 9772 23248
rect 9824 23236 9830 23248
rect 11333 23239 11391 23245
rect 11333 23236 11345 23239
rect 9824 23208 11345 23236
rect 9824 23196 9830 23208
rect 11333 23205 11345 23208
rect 11379 23205 11391 23239
rect 11333 23199 11391 23205
rect 12434 23196 12440 23248
rect 12492 23236 12498 23248
rect 12989 23239 13047 23245
rect 12989 23236 13001 23239
rect 12492 23208 13001 23236
rect 12492 23196 12498 23208
rect 12989 23205 13001 23208
rect 13035 23205 13047 23239
rect 12989 23199 13047 23205
rect 24486 23196 24492 23248
rect 24544 23236 24550 23248
rect 24544 23208 25176 23236
rect 24544 23196 24550 23208
rect 2866 23128 2872 23180
rect 2924 23168 2930 23180
rect 2961 23171 3019 23177
rect 2961 23168 2973 23171
rect 2924 23140 2973 23168
rect 2924 23128 2930 23140
rect 2961 23137 2973 23140
rect 3007 23168 3019 23171
rect 3418 23168 3424 23180
rect 3007 23140 3424 23168
rect 3007 23137 3019 23140
rect 2961 23131 3019 23137
rect 3418 23128 3424 23140
rect 3476 23128 3482 23180
rect 5074 23168 5080 23180
rect 3620 23140 5080 23168
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23069 2283 23103
rect 2225 23063 2283 23069
rect 2777 23103 2835 23109
rect 2777 23069 2789 23103
rect 2823 23100 2835 23103
rect 3620 23100 3648 23140
rect 5074 23128 5080 23140
rect 5132 23128 5138 23180
rect 5718 23128 5724 23180
rect 5776 23168 5782 23180
rect 5813 23171 5871 23177
rect 5813 23168 5825 23171
rect 5776 23140 5825 23168
rect 5776 23128 5782 23140
rect 5813 23137 5825 23140
rect 5859 23168 5871 23171
rect 6454 23168 6460 23180
rect 5859 23140 6460 23168
rect 5859 23137 5871 23140
rect 5813 23131 5871 23137
rect 6454 23128 6460 23140
rect 6512 23128 6518 23180
rect 7374 23168 7380 23180
rect 7208 23140 7380 23168
rect 2823 23072 3648 23100
rect 2823 23069 2835 23072
rect 2777 23063 2835 23069
rect 2240 23032 2268 23063
rect 3694 23060 3700 23112
rect 3752 23100 3758 23112
rect 4100 23103 4158 23109
rect 4100 23100 4112 23103
rect 3752 23072 4112 23100
rect 3752 23060 3758 23072
rect 4100 23069 4112 23072
rect 4146 23069 4158 23103
rect 4100 23063 4158 23069
rect 4203 23103 4261 23109
rect 4203 23069 4215 23103
rect 4249 23100 4261 23103
rect 4338 23100 4344 23112
rect 4249 23072 4344 23100
rect 4249 23069 4261 23072
rect 4203 23063 4261 23069
rect 4338 23060 4344 23072
rect 4396 23060 4402 23112
rect 7208 23086 7236 23140
rect 7374 23128 7380 23140
rect 7432 23168 7438 23180
rect 7852 23168 7880 23196
rect 7432 23140 7880 23168
rect 7432 23128 7438 23140
rect 10042 23128 10048 23180
rect 10100 23168 10106 23180
rect 10778 23168 10784 23180
rect 10100 23140 10784 23168
rect 10100 23128 10106 23140
rect 10778 23128 10784 23140
rect 10836 23128 10842 23180
rect 11606 23128 11612 23180
rect 11664 23168 11670 23180
rect 11885 23171 11943 23177
rect 11885 23168 11897 23171
rect 11664 23140 11897 23168
rect 11664 23128 11670 23140
rect 11885 23137 11897 23140
rect 11931 23137 11943 23171
rect 11885 23131 11943 23137
rect 12618 23128 12624 23180
rect 12676 23168 12682 23180
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 12676 23140 13553 23168
rect 12676 23128 12682 23140
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 13541 23131 13599 23137
rect 14274 23128 14280 23180
rect 14332 23168 14338 23180
rect 15286 23168 15292 23180
rect 14332 23140 15292 23168
rect 14332 23128 14338 23140
rect 15286 23128 15292 23140
rect 15344 23168 15350 23180
rect 16485 23171 16543 23177
rect 16485 23168 16497 23171
rect 15344 23140 16497 23168
rect 15344 23128 15350 23140
rect 16485 23137 16497 23140
rect 16531 23168 16543 23171
rect 18598 23168 18604 23180
rect 16531 23140 18604 23168
rect 16531 23137 16543 23140
rect 16485 23131 16543 23137
rect 18598 23128 18604 23140
rect 18656 23168 18662 23180
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 18656 23140 19441 23168
rect 18656 23128 18662 23140
rect 19429 23137 19441 23140
rect 19475 23137 19487 23171
rect 19429 23131 19487 23137
rect 22005 23171 22063 23177
rect 22005 23137 22017 23171
rect 22051 23168 22063 23171
rect 22051 23140 23520 23168
rect 22051 23137 22063 23140
rect 22005 23131 22063 23137
rect 9953 23103 10011 23109
rect 9953 23069 9965 23103
rect 9999 23100 10011 23103
rect 10962 23100 10968 23112
rect 9999 23072 10968 23100
rect 9999 23069 10011 23072
rect 9953 23063 10011 23069
rect 10962 23060 10968 23072
rect 11020 23060 11026 23112
rect 11698 23060 11704 23112
rect 11756 23060 11762 23112
rect 11793 23103 11851 23109
rect 11793 23069 11805 23103
rect 11839 23100 11851 23103
rect 12158 23100 12164 23112
rect 11839 23072 12164 23100
rect 11839 23069 11851 23072
rect 11793 23063 11851 23069
rect 12158 23060 12164 23072
rect 12216 23060 12222 23112
rect 13357 23103 13415 23109
rect 13357 23069 13369 23103
rect 13403 23100 13415 23103
rect 13906 23100 13912 23112
rect 13403 23072 13912 23100
rect 13403 23069 13415 23072
rect 13357 23063 13415 23069
rect 13906 23060 13912 23072
rect 13964 23060 13970 23112
rect 16114 23100 16120 23112
rect 15686 23072 16120 23100
rect 16114 23060 16120 23072
rect 16172 23100 16178 23112
rect 16390 23100 16396 23112
rect 16172 23072 16396 23100
rect 16172 23060 16178 23072
rect 16390 23060 16396 23072
rect 16448 23060 16454 23112
rect 22833 23103 22891 23109
rect 22833 23069 22845 23103
rect 22879 23069 22891 23103
rect 23492 23100 23520 23140
rect 23842 23128 23848 23180
rect 23900 23128 23906 23180
rect 24578 23128 24584 23180
rect 24636 23168 24642 23180
rect 25148 23177 25176 23208
rect 25041 23171 25099 23177
rect 25041 23168 25053 23171
rect 24636 23140 25053 23168
rect 24636 23128 24642 23140
rect 25041 23137 25053 23140
rect 25087 23137 25099 23171
rect 25041 23131 25099 23137
rect 25133 23171 25191 23177
rect 25133 23137 25145 23171
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 24949 23103 25007 23109
rect 24949 23100 24961 23103
rect 23492 23072 24961 23100
rect 22833 23063 22891 23069
rect 24949 23069 24961 23072
rect 24995 23069 25007 23103
rect 24949 23063 25007 23069
rect 3786 23032 3792 23044
rect 2240 23004 3792 23032
rect 3786 22992 3792 23004
rect 3844 22992 3850 23044
rect 6089 23035 6147 23041
rect 6089 23001 6101 23035
rect 6135 23001 6147 23035
rect 7742 23032 7748 23044
rect 6089 22995 6147 23001
rect 7484 23004 7748 23032
rect 6104 22964 6132 22995
rect 7484 22964 7512 23004
rect 7742 22992 7748 23004
rect 7800 22992 7806 23044
rect 10689 23035 10747 23041
rect 10689 23001 10701 23035
rect 10735 23001 10747 23035
rect 10689 22995 10747 23001
rect 6104 22936 7512 22964
rect 9950 22924 9956 22976
rect 10008 22964 10014 22976
rect 10704 22964 10732 22995
rect 10778 22992 10784 23044
rect 10836 23032 10842 23044
rect 12529 23035 12587 23041
rect 12529 23032 12541 23035
rect 10836 23004 12541 23032
rect 10836 22992 10842 23004
rect 12529 23001 12541 23004
rect 12575 23032 12587 23035
rect 13449 23035 13507 23041
rect 13449 23032 13461 23035
rect 12575 23004 13461 23032
rect 12575 23001 12587 23004
rect 12529 22995 12587 23001
rect 13449 23001 13461 23004
rect 13495 23001 13507 23035
rect 13449 22995 13507 23001
rect 14553 23035 14611 23041
rect 14553 23001 14565 23035
rect 14599 23001 14611 23035
rect 14553 22995 14611 23001
rect 10008 22936 10732 22964
rect 10008 22924 10014 22936
rect 12618 22924 12624 22976
rect 12676 22924 12682 22976
rect 13078 22924 13084 22976
rect 13136 22964 13142 22976
rect 14568 22964 14596 22995
rect 15930 22992 15936 23044
rect 15988 23032 15994 23044
rect 16761 23035 16819 23041
rect 16761 23032 16773 23035
rect 15988 23004 16773 23032
rect 15988 22992 15994 23004
rect 16761 23001 16773 23004
rect 16807 23001 16819 23035
rect 16761 22995 16819 23001
rect 17770 22992 17776 23044
rect 17828 22992 17834 23044
rect 19705 23035 19763 23041
rect 19705 23032 19717 23035
rect 18248 23004 19717 23032
rect 15378 22964 15384 22976
rect 13136 22936 15384 22964
rect 13136 22924 13142 22936
rect 15378 22924 15384 22936
rect 15436 22924 15442 22976
rect 15470 22924 15476 22976
rect 15528 22964 15534 22976
rect 15838 22964 15844 22976
rect 15528 22936 15844 22964
rect 15528 22924 15534 22936
rect 15838 22924 15844 22936
rect 15896 22924 15902 22976
rect 16206 22924 16212 22976
rect 16264 22964 16270 22976
rect 16482 22964 16488 22976
rect 16264 22936 16488 22964
rect 16264 22924 16270 22936
rect 16482 22924 16488 22936
rect 16540 22924 16546 22976
rect 18248 22973 18276 23004
rect 19705 23001 19717 23004
rect 19751 23032 19763 23035
rect 19978 23032 19984 23044
rect 19751 23004 19984 23032
rect 19751 23001 19763 23004
rect 19705 22995 19763 23001
rect 19978 22992 19984 23004
rect 20036 22992 20042 23044
rect 22848 23032 22876 23063
rect 25406 23032 25412 23044
rect 20088 23004 20194 23032
rect 22848 23004 25412 23032
rect 18233 22967 18291 22973
rect 18233 22933 18245 22967
rect 18279 22933 18291 22967
rect 18233 22927 18291 22933
rect 19334 22924 19340 22976
rect 19392 22964 19398 22976
rect 20088 22964 20116 23004
rect 25406 22992 25412 23004
rect 25464 22992 25470 23044
rect 21082 22964 21088 22976
rect 19392 22936 21088 22964
rect 19392 22924 19398 22936
rect 21082 22924 21088 22936
rect 21140 22964 21146 22976
rect 21453 22967 21511 22973
rect 21453 22964 21465 22967
rect 21140 22936 21465 22964
rect 21140 22924 21146 22936
rect 21453 22933 21465 22936
rect 21499 22964 21511 22967
rect 22830 22964 22836 22976
rect 21499 22936 22836 22964
rect 21499 22933 21511 22936
rect 21453 22927 21511 22933
rect 22830 22924 22836 22936
rect 22888 22924 22894 22976
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 23532 22936 24593 22964
rect 23532 22924 23538 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 1762 22720 1768 22772
rect 1820 22760 1826 22772
rect 2041 22763 2099 22769
rect 2041 22760 2053 22763
rect 1820 22732 2053 22760
rect 1820 22720 1826 22732
rect 2041 22729 2053 22732
rect 2087 22729 2099 22763
rect 2041 22723 2099 22729
rect 5629 22763 5687 22769
rect 5629 22729 5641 22763
rect 5675 22760 5687 22763
rect 6825 22763 6883 22769
rect 6825 22760 6837 22763
rect 5675 22732 6837 22760
rect 5675 22729 5687 22732
rect 5629 22723 5687 22729
rect 6825 22729 6837 22732
rect 6871 22729 6883 22763
rect 6825 22723 6883 22729
rect 7193 22763 7251 22769
rect 7193 22729 7205 22763
rect 7239 22760 7251 22763
rect 9398 22760 9404 22772
rect 7239 22732 9404 22760
rect 7239 22729 7251 22732
rect 7193 22723 7251 22729
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 10042 22720 10048 22772
rect 10100 22760 10106 22772
rect 10137 22763 10195 22769
rect 10137 22760 10149 22763
rect 10100 22732 10149 22760
rect 10100 22720 10106 22732
rect 10137 22729 10149 22732
rect 10183 22760 10195 22763
rect 10873 22763 10931 22769
rect 10873 22760 10885 22763
rect 10183 22732 10885 22760
rect 10183 22729 10195 22732
rect 10137 22723 10195 22729
rect 10873 22729 10885 22732
rect 10919 22760 10931 22763
rect 12066 22760 12072 22772
rect 10919 22732 12072 22760
rect 10919 22729 10931 22732
rect 10873 22723 10931 22729
rect 12066 22720 12072 22732
rect 12124 22720 12130 22772
rect 12345 22763 12403 22769
rect 12345 22729 12357 22763
rect 12391 22760 12403 22763
rect 12802 22760 12808 22772
rect 12391 22732 12808 22760
rect 12391 22729 12403 22732
rect 12345 22723 12403 22729
rect 12802 22720 12808 22732
rect 12860 22720 12866 22772
rect 13078 22720 13084 22772
rect 13136 22720 13142 22772
rect 15102 22720 15108 22772
rect 15160 22760 15166 22772
rect 15197 22763 15255 22769
rect 15197 22760 15209 22763
rect 15160 22732 15209 22760
rect 15160 22720 15166 22732
rect 15197 22729 15209 22732
rect 15243 22729 15255 22763
rect 15197 22723 15255 22729
rect 15378 22720 15384 22772
rect 15436 22760 15442 22772
rect 16022 22760 16028 22772
rect 15436 22732 16028 22760
rect 15436 22720 15442 22732
rect 16022 22720 16028 22732
rect 16080 22760 16086 22772
rect 16209 22763 16267 22769
rect 16209 22760 16221 22763
rect 16080 22732 16221 22760
rect 16080 22720 16086 22732
rect 16209 22729 16221 22732
rect 16255 22760 16267 22763
rect 16255 22732 16528 22760
rect 16255 22729 16267 22732
rect 16209 22723 16267 22729
rect 11514 22652 11520 22704
rect 11572 22692 11578 22704
rect 11882 22692 11888 22704
rect 11572 22664 11888 22692
rect 11572 22652 11578 22664
rect 11882 22652 11888 22664
rect 11940 22692 11946 22704
rect 12437 22695 12495 22701
rect 12437 22692 12449 22695
rect 11940 22664 12449 22692
rect 11940 22652 11946 22664
rect 12437 22661 12449 22664
rect 12483 22661 12495 22695
rect 13265 22695 13323 22701
rect 13265 22692 13277 22695
rect 12437 22655 12495 22661
rect 12728 22664 13277 22692
rect 2225 22627 2283 22633
rect 2225 22593 2237 22627
rect 2271 22624 2283 22627
rect 2866 22624 2872 22636
rect 2271 22596 2872 22624
rect 2271 22593 2283 22596
rect 2225 22587 2283 22593
rect 2866 22584 2872 22596
rect 2924 22584 2930 22636
rect 5721 22627 5779 22633
rect 5721 22593 5733 22627
rect 5767 22624 5779 22627
rect 7834 22624 7840 22636
rect 5767 22596 7840 22624
rect 5767 22593 5779 22596
rect 5721 22587 5779 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 8021 22627 8079 22633
rect 8021 22593 8033 22627
rect 8067 22624 8079 22627
rect 9217 22627 9275 22633
rect 9217 22624 9229 22627
rect 8067 22596 9229 22624
rect 8067 22593 8079 22596
rect 8021 22587 8079 22593
rect 9217 22593 9229 22596
rect 9263 22624 9275 22627
rect 9674 22624 9680 22636
rect 9263 22596 9680 22624
rect 9263 22593 9275 22596
rect 9217 22587 9275 22593
rect 9674 22584 9680 22596
rect 9732 22584 9738 22636
rect 10781 22627 10839 22633
rect 10781 22593 10793 22627
rect 10827 22624 10839 22627
rect 12728 22624 12756 22664
rect 13265 22661 13277 22664
rect 13311 22692 13323 22695
rect 15286 22692 15292 22704
rect 13311 22664 15292 22692
rect 13311 22661 13323 22664
rect 13265 22655 13323 22661
rect 15286 22652 15292 22664
rect 15344 22652 15350 22704
rect 16114 22652 16120 22704
rect 16172 22692 16178 22704
rect 16301 22695 16359 22701
rect 16301 22692 16313 22695
rect 16172 22664 16313 22692
rect 16172 22652 16178 22664
rect 16301 22661 16313 22664
rect 16347 22661 16359 22695
rect 16301 22655 16359 22661
rect 10827 22596 12296 22624
rect 10827 22593 10839 22596
rect 10781 22587 10839 22593
rect 5905 22559 5963 22565
rect 5905 22525 5917 22559
rect 5951 22556 5963 22559
rect 5994 22556 6000 22568
rect 5951 22528 6000 22556
rect 5951 22525 5963 22528
rect 5905 22519 5963 22525
rect 5994 22516 6000 22528
rect 6052 22516 6058 22568
rect 7282 22516 7288 22568
rect 7340 22516 7346 22568
rect 7469 22559 7527 22565
rect 7469 22525 7481 22559
rect 7515 22556 7527 22559
rect 7558 22556 7564 22568
rect 7515 22528 7564 22556
rect 7515 22525 7527 22528
rect 7469 22519 7527 22525
rect 7558 22516 7564 22528
rect 7616 22516 7622 22568
rect 8846 22516 8852 22568
rect 8904 22516 8910 22568
rect 10965 22559 11023 22565
rect 10965 22525 10977 22559
rect 11011 22556 11023 22559
rect 11146 22556 11152 22568
rect 11011 22528 11152 22556
rect 11011 22525 11023 22528
rect 10965 22519 11023 22525
rect 11146 22516 11152 22528
rect 11204 22516 11210 22568
rect 12268 22556 12296 22596
rect 12406 22596 12756 22624
rect 12406 22556 12434 22596
rect 13814 22584 13820 22636
rect 13872 22624 13878 22636
rect 15105 22627 15163 22633
rect 15105 22624 15117 22627
rect 13872 22596 15117 22624
rect 13872 22584 13878 22596
rect 15105 22593 15117 22596
rect 15151 22593 15163 22627
rect 16500 22624 16528 22732
rect 16574 22720 16580 22772
rect 16632 22760 16638 22772
rect 17494 22760 17500 22772
rect 16632 22732 17500 22760
rect 16632 22720 16638 22732
rect 17494 22720 17500 22732
rect 17552 22760 17558 22772
rect 20346 22760 20352 22772
rect 17552 22732 20352 22760
rect 17552 22720 17558 22732
rect 17880 22701 17908 22732
rect 20346 22720 20352 22732
rect 20404 22720 20410 22772
rect 23290 22720 23296 22772
rect 23348 22760 23354 22772
rect 23348 22732 23612 22760
rect 23348 22720 23354 22732
rect 17865 22695 17923 22701
rect 17865 22661 17877 22695
rect 17911 22661 17923 22695
rect 17865 22655 17923 22661
rect 18598 22652 18604 22704
rect 18656 22652 18662 22704
rect 19702 22652 19708 22704
rect 19760 22652 19766 22704
rect 20364 22692 20392 22720
rect 20533 22695 20591 22701
rect 20533 22692 20545 22695
rect 20364 22664 20545 22692
rect 20533 22661 20545 22664
rect 20579 22661 20591 22695
rect 23584 22692 23612 22732
rect 23658 22720 23664 22772
rect 23716 22760 23722 22772
rect 23753 22763 23811 22769
rect 23753 22760 23765 22763
rect 23716 22732 23765 22760
rect 23716 22720 23722 22732
rect 23753 22729 23765 22732
rect 23799 22729 23811 22763
rect 23753 22723 23811 22729
rect 24213 22763 24271 22769
rect 24213 22729 24225 22763
rect 24259 22760 24271 22763
rect 24302 22760 24308 22772
rect 24259 22732 24308 22760
rect 24259 22729 24271 22732
rect 24213 22723 24271 22729
rect 24228 22692 24256 22723
rect 24302 22720 24308 22732
rect 24360 22760 24366 22772
rect 24765 22763 24823 22769
rect 24765 22760 24777 22763
rect 24360 22732 24777 22760
rect 24360 22720 24366 22732
rect 24765 22729 24777 22732
rect 24811 22729 24823 22763
rect 24765 22723 24823 22729
rect 25314 22720 25320 22772
rect 25372 22760 25378 22772
rect 25409 22763 25467 22769
rect 25409 22760 25421 22763
rect 25372 22732 25421 22760
rect 25372 22720 25378 22732
rect 25409 22729 25421 22732
rect 25455 22729 25467 22763
rect 25409 22723 25467 22729
rect 23506 22664 24256 22692
rect 20533 22655 20591 22661
rect 18322 22624 18328 22636
rect 16500 22596 18328 22624
rect 15105 22587 15163 22593
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 19334 22584 19340 22636
rect 19392 22624 19398 22636
rect 19613 22627 19671 22633
rect 19613 22624 19625 22627
rect 19392 22596 19625 22624
rect 19392 22584 19398 22596
rect 19613 22593 19625 22596
rect 19659 22593 19671 22627
rect 19613 22587 19671 22593
rect 21361 22627 21419 22633
rect 21361 22593 21373 22627
rect 21407 22624 21419 22627
rect 22002 22624 22008 22636
rect 21407 22596 22008 22624
rect 21407 22593 21419 22596
rect 21361 22587 21419 22593
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 23658 22584 23664 22636
rect 23716 22624 23722 22636
rect 24486 22624 24492 22636
rect 23716 22596 24492 22624
rect 23716 22584 23722 22596
rect 24486 22584 24492 22596
rect 24544 22584 24550 22636
rect 12268 22528 12434 22556
rect 12621 22559 12679 22565
rect 12621 22525 12633 22559
rect 12667 22556 12679 22559
rect 13078 22556 13084 22568
rect 12667 22528 13084 22556
rect 12667 22525 12679 22528
rect 12621 22519 12679 22525
rect 13078 22516 13084 22528
rect 13136 22516 13142 22568
rect 13906 22516 13912 22568
rect 13964 22516 13970 22568
rect 15381 22559 15439 22565
rect 15381 22525 15393 22559
rect 15427 22556 15439 22559
rect 15930 22556 15936 22568
rect 15427 22528 15936 22556
rect 15427 22525 15439 22528
rect 15381 22519 15439 22525
rect 15930 22516 15936 22528
rect 15988 22516 15994 22568
rect 19058 22516 19064 22568
rect 19116 22556 19122 22568
rect 19797 22559 19855 22565
rect 19797 22556 19809 22559
rect 19116 22528 19809 22556
rect 19116 22516 19122 22528
rect 19797 22525 19809 22528
rect 19843 22556 19855 22559
rect 21174 22556 21180 22568
rect 19843 22528 21180 22556
rect 19843 22525 19855 22528
rect 19797 22519 19855 22525
rect 21174 22516 21180 22528
rect 21232 22516 21238 22568
rect 21634 22516 21640 22568
rect 21692 22556 21698 22568
rect 22281 22559 22339 22565
rect 22281 22556 22293 22559
rect 21692 22528 22293 22556
rect 21692 22516 21698 22528
rect 22281 22525 22293 22528
rect 22327 22525 22339 22559
rect 22281 22519 22339 22525
rect 9398 22448 9404 22500
rect 9456 22488 9462 22500
rect 10413 22491 10471 22497
rect 10413 22488 10425 22491
rect 9456 22460 10425 22488
rect 9456 22448 9462 22460
rect 10413 22457 10425 22460
rect 10459 22457 10471 22491
rect 10413 22451 10471 22457
rect 11977 22491 12035 22497
rect 11977 22457 11989 22491
rect 12023 22488 12035 22491
rect 13998 22488 14004 22500
rect 12023 22460 14004 22488
rect 12023 22457 12035 22460
rect 11977 22451 12035 22457
rect 13998 22448 14004 22460
rect 14056 22448 14062 22500
rect 4246 22380 4252 22432
rect 4304 22420 4310 22432
rect 5261 22423 5319 22429
rect 5261 22420 5273 22423
rect 4304 22392 5273 22420
rect 4304 22380 4310 22392
rect 5261 22389 5273 22392
rect 5307 22389 5319 22423
rect 5261 22383 5319 22389
rect 6914 22380 6920 22432
rect 6972 22420 6978 22432
rect 10778 22420 10784 22432
rect 6972 22392 10784 22420
rect 6972 22380 6978 22392
rect 10778 22380 10784 22392
rect 10836 22380 10842 22432
rect 11514 22380 11520 22432
rect 11572 22420 11578 22432
rect 11609 22423 11667 22429
rect 11609 22420 11621 22423
rect 11572 22392 11621 22420
rect 11572 22380 11578 22392
rect 11609 22389 11621 22392
rect 11655 22389 11667 22423
rect 11609 22383 11667 22389
rect 14737 22423 14795 22429
rect 14737 22389 14749 22423
rect 14783 22420 14795 22423
rect 15562 22420 15568 22432
rect 14783 22392 15568 22420
rect 14783 22389 14795 22392
rect 14737 22383 14795 22389
rect 15562 22380 15568 22392
rect 15620 22380 15626 22432
rect 18782 22380 18788 22432
rect 18840 22420 18846 22432
rect 18966 22420 18972 22432
rect 18840 22392 18972 22420
rect 18840 22380 18846 22392
rect 18966 22380 18972 22392
rect 19024 22380 19030 22432
rect 19242 22380 19248 22432
rect 19300 22380 19306 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 16114 22176 16120 22228
rect 16172 22216 16178 22228
rect 16301 22219 16359 22225
rect 16301 22216 16313 22219
rect 16172 22188 16313 22216
rect 16172 22176 16178 22188
rect 16301 22185 16313 22188
rect 16347 22216 16359 22219
rect 16390 22216 16396 22228
rect 16347 22188 16396 22216
rect 16347 22185 16359 22188
rect 16301 22179 16359 22185
rect 16390 22176 16396 22188
rect 16448 22176 16454 22228
rect 18598 22216 18604 22228
rect 17512 22188 18604 22216
rect 7466 22108 7472 22160
rect 7524 22148 7530 22160
rect 11514 22148 11520 22160
rect 7524 22120 11520 22148
rect 7524 22108 7530 22120
rect 11514 22108 11520 22120
rect 11572 22108 11578 22160
rect 16853 22151 16911 22157
rect 11992 22120 13768 22148
rect 11992 22089 12020 22120
rect 11977 22083 12035 22089
rect 11977 22080 11989 22083
rect 11935 22052 11989 22080
rect 11977 22049 11989 22052
rect 12023 22080 12035 22083
rect 12158 22080 12164 22092
rect 12023 22052 12164 22080
rect 12023 22049 12035 22052
rect 11977 22043 12035 22049
rect 12158 22040 12164 22052
rect 12216 22040 12222 22092
rect 11146 21972 11152 22024
rect 11204 22012 11210 22024
rect 11882 22012 11888 22024
rect 11204 21984 11888 22012
rect 11204 21972 11210 21984
rect 11882 21972 11888 21984
rect 11940 21972 11946 22024
rect 13265 22015 13323 22021
rect 13265 21981 13277 22015
rect 13311 22012 13323 22015
rect 13630 22012 13636 22024
rect 13311 21984 13636 22012
rect 13311 21981 13323 21984
rect 13265 21975 13323 21981
rect 13630 21972 13636 21984
rect 13688 21972 13694 22024
rect 11793 21947 11851 21953
rect 10888 21916 11560 21944
rect 4430 21836 4436 21888
rect 4488 21876 4494 21888
rect 4706 21876 4712 21888
rect 4488 21848 4712 21876
rect 4488 21836 4494 21848
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 8570 21836 8576 21888
rect 8628 21876 8634 21888
rect 8754 21876 8760 21888
rect 8628 21848 8760 21876
rect 8628 21836 8634 21848
rect 8754 21836 8760 21848
rect 8812 21836 8818 21888
rect 10226 21836 10232 21888
rect 10284 21876 10290 21888
rect 10888 21885 10916 21916
rect 10873 21879 10931 21885
rect 10873 21876 10885 21879
rect 10284 21848 10885 21876
rect 10284 21836 10290 21848
rect 10873 21845 10885 21848
rect 10919 21845 10931 21879
rect 10873 21839 10931 21845
rect 11422 21836 11428 21888
rect 11480 21836 11486 21888
rect 11532 21876 11560 21916
rect 11793 21913 11805 21947
rect 11839 21944 11851 21947
rect 12529 21947 12587 21953
rect 12529 21944 12541 21947
rect 11839 21916 12541 21944
rect 11839 21913 11851 21916
rect 11793 21907 11851 21913
rect 12529 21913 12541 21916
rect 12575 21944 12587 21947
rect 13538 21944 13544 21956
rect 12575 21916 13544 21944
rect 12575 21913 12587 21916
rect 12529 21907 12587 21913
rect 13538 21904 13544 21916
rect 13596 21904 13602 21956
rect 13740 21944 13768 22120
rect 16853 22117 16865 22151
rect 16899 22117 16911 22151
rect 16853 22111 16911 22117
rect 14274 22040 14280 22092
rect 14332 22040 14338 22092
rect 16025 22083 16083 22089
rect 16025 22049 16037 22083
rect 16071 22080 16083 22083
rect 16114 22080 16120 22092
rect 16071 22052 16120 22080
rect 16071 22049 16083 22052
rect 16025 22043 16083 22049
rect 16114 22040 16120 22052
rect 16172 22040 16178 22092
rect 13740 21916 14136 21944
rect 11885 21879 11943 21885
rect 11885 21876 11897 21879
rect 11532 21848 11897 21876
rect 11885 21845 11897 21848
rect 11931 21845 11943 21879
rect 11885 21839 11943 21845
rect 13081 21879 13139 21885
rect 13081 21845 13093 21879
rect 13127 21876 13139 21879
rect 13354 21876 13360 21888
rect 13127 21848 13360 21876
rect 13127 21845 13139 21848
rect 13081 21839 13139 21845
rect 13354 21836 13360 21848
rect 13412 21836 13418 21888
rect 14108 21876 14136 21916
rect 14550 21904 14556 21956
rect 14608 21904 14614 21956
rect 16390 21944 16396 21956
rect 15778 21916 16396 21944
rect 16390 21904 16396 21916
rect 16448 21904 16454 21956
rect 16868 21944 16896 22111
rect 17512 22089 17540 22188
rect 18598 22176 18604 22188
rect 18656 22176 18662 22228
rect 19686 22219 19744 22225
rect 19686 22216 19698 22219
rect 18708 22188 19698 22216
rect 18049 22151 18107 22157
rect 18049 22117 18061 22151
rect 18095 22117 18107 22151
rect 18049 22111 18107 22117
rect 17497 22083 17555 22089
rect 17497 22049 17509 22083
rect 17543 22080 17555 22083
rect 17543 22052 17577 22080
rect 17543 22049 17555 22052
rect 17497 22043 17555 22049
rect 17034 21972 17040 22024
rect 17092 22012 17098 22024
rect 17221 22015 17279 22021
rect 17221 22012 17233 22015
rect 17092 21984 17233 22012
rect 17092 21972 17098 21984
rect 17221 21981 17233 21984
rect 17267 21981 17279 22015
rect 18064 22012 18092 22111
rect 18506 22040 18512 22092
rect 18564 22040 18570 22092
rect 18708 22089 18736 22188
rect 19686 22185 19698 22188
rect 19732 22216 19744 22219
rect 20254 22216 20260 22228
rect 19732 22188 20260 22216
rect 19732 22185 19744 22188
rect 19686 22179 19744 22185
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 21174 22176 21180 22228
rect 21232 22176 21238 22228
rect 18693 22083 18751 22089
rect 18693 22049 18705 22083
rect 18739 22049 18751 22083
rect 22002 22080 22008 22092
rect 18693 22043 18751 22049
rect 19444 22052 22008 22080
rect 19444 22024 19472 22052
rect 22002 22040 22008 22052
rect 22060 22040 22066 22092
rect 22278 22040 22284 22092
rect 22336 22040 22342 22092
rect 22370 22040 22376 22092
rect 22428 22080 22434 22092
rect 23290 22080 23296 22092
rect 22428 22052 23296 22080
rect 22428 22040 22434 22052
rect 23290 22040 23296 22052
rect 23348 22040 23354 22092
rect 24029 22083 24087 22089
rect 24029 22049 24041 22083
rect 24075 22080 24087 22083
rect 24210 22080 24216 22092
rect 24075 22052 24216 22080
rect 24075 22049 24087 22052
rect 24029 22043 24087 22049
rect 24210 22040 24216 22052
rect 24268 22040 24274 22092
rect 19334 22012 19340 22024
rect 18064 21984 19340 22012
rect 17221 21975 17279 21981
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 19426 21972 19432 22024
rect 19484 21972 19490 22024
rect 24118 21972 24124 22024
rect 24176 22012 24182 22024
rect 24857 22015 24915 22021
rect 24857 22012 24869 22015
rect 24176 21984 24869 22012
rect 24176 21972 24182 21984
rect 24857 21981 24869 21984
rect 24903 21981 24915 22015
rect 24857 21975 24915 21981
rect 18417 21947 18475 21953
rect 18417 21944 18429 21947
rect 16868 21916 18429 21944
rect 18417 21913 18429 21916
rect 18463 21913 18475 21947
rect 21453 21947 21511 21953
rect 21453 21944 21465 21947
rect 20930 21916 21465 21944
rect 18417 21907 18475 21913
rect 21453 21913 21465 21916
rect 21499 21944 21511 21947
rect 22370 21944 22376 21956
rect 21499 21916 22376 21944
rect 21499 21913 21511 21916
rect 21453 21907 21511 21913
rect 22370 21904 22376 21916
rect 22428 21944 22434 21956
rect 24673 21947 24731 21953
rect 22428 21916 22770 21944
rect 22428 21904 22434 21916
rect 24673 21913 24685 21947
rect 24719 21913 24731 21947
rect 24673 21907 24731 21913
rect 15378 21876 15384 21888
rect 14108 21848 15384 21876
rect 15378 21836 15384 21848
rect 15436 21836 15442 21888
rect 15930 21836 15936 21888
rect 15988 21876 15994 21888
rect 16577 21879 16635 21885
rect 16577 21876 16589 21879
rect 15988 21848 16589 21876
rect 15988 21836 15994 21848
rect 16577 21845 16589 21848
rect 16623 21876 16635 21879
rect 17313 21879 17371 21885
rect 17313 21876 17325 21879
rect 16623 21848 17325 21876
rect 16623 21845 16635 21848
rect 16577 21839 16635 21845
rect 17313 21845 17325 21848
rect 17359 21876 17371 21879
rect 19978 21876 19984 21888
rect 17359 21848 19984 21876
rect 17359 21845 17371 21848
rect 17313 21839 17371 21845
rect 19978 21836 19984 21848
rect 20036 21836 20042 21888
rect 21542 21836 21548 21888
rect 21600 21876 21606 21888
rect 24688 21876 24716 21907
rect 21600 21848 24716 21876
rect 21600 21836 21606 21848
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 7098 21632 7104 21684
rect 7156 21632 7162 21684
rect 7469 21675 7527 21681
rect 7469 21641 7481 21675
rect 7515 21672 7527 21675
rect 8297 21675 8355 21681
rect 8297 21672 8309 21675
rect 7515 21644 8309 21672
rect 7515 21641 7527 21644
rect 7469 21635 7527 21641
rect 8297 21641 8309 21644
rect 8343 21641 8355 21675
rect 8297 21635 8355 21641
rect 8665 21675 8723 21681
rect 8665 21641 8677 21675
rect 8711 21672 8723 21675
rect 9766 21672 9772 21684
rect 8711 21644 9772 21672
rect 8711 21641 8723 21644
rect 8665 21635 8723 21641
rect 9766 21632 9772 21644
rect 9824 21632 9830 21684
rect 9861 21675 9919 21681
rect 9861 21641 9873 21675
rect 9907 21672 9919 21675
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 9907 21644 11713 21672
rect 9907 21641 9919 21644
rect 9861 21635 9919 21641
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 11701 21635 11759 21641
rect 11974 21632 11980 21684
rect 12032 21672 12038 21684
rect 12069 21675 12127 21681
rect 12069 21672 12081 21675
rect 12032 21644 12081 21672
rect 12032 21632 12038 21644
rect 12069 21641 12081 21644
rect 12115 21641 12127 21675
rect 12069 21635 12127 21641
rect 13541 21675 13599 21681
rect 13541 21641 13553 21675
rect 13587 21672 13599 21675
rect 13814 21672 13820 21684
rect 13587 21644 13820 21672
rect 13587 21641 13599 21644
rect 13541 21635 13599 21641
rect 13814 21632 13820 21644
rect 13872 21632 13878 21684
rect 13906 21632 13912 21684
rect 13964 21632 13970 21684
rect 13998 21632 14004 21684
rect 14056 21632 14062 21684
rect 14734 21632 14740 21684
rect 14792 21672 14798 21684
rect 14792 21644 18736 21672
rect 14792 21632 14798 21644
rect 7650 21564 7656 21616
rect 7708 21604 7714 21616
rect 7708 21576 10088 21604
rect 7708 21564 7714 21576
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21536 1823 21539
rect 1854 21536 1860 21548
rect 1811 21508 1860 21536
rect 1811 21505 1823 21508
rect 1765 21499 1823 21505
rect 1854 21496 1860 21508
rect 1912 21496 1918 21548
rect 3421 21539 3479 21545
rect 3421 21505 3433 21539
rect 3467 21536 3479 21539
rect 4430 21536 4436 21548
rect 3467 21508 4436 21536
rect 3467 21505 3479 21508
rect 3421 21499 3479 21505
rect 4430 21496 4436 21508
rect 4488 21496 4494 21548
rect 4525 21539 4583 21545
rect 4525 21505 4537 21539
rect 4571 21536 4583 21539
rect 4706 21536 4712 21548
rect 4571 21508 4712 21536
rect 4571 21505 4583 21508
rect 4525 21499 4583 21505
rect 4706 21496 4712 21508
rect 4764 21496 4770 21548
rect 7561 21539 7619 21545
rect 7561 21505 7573 21539
rect 7607 21536 7619 21539
rect 8938 21536 8944 21548
rect 7607 21508 8944 21536
rect 7607 21505 7619 21508
rect 7561 21499 7619 21505
rect 8938 21496 8944 21508
rect 8996 21496 9002 21548
rect 1302 21428 1308 21480
rect 1360 21468 1366 21480
rect 2041 21471 2099 21477
rect 2041 21468 2053 21471
rect 1360 21440 2053 21468
rect 1360 21428 1366 21440
rect 2041 21437 2053 21440
rect 2087 21437 2099 21471
rect 2041 21431 2099 21437
rect 3602 21428 3608 21480
rect 3660 21468 3666 21480
rect 4062 21468 4068 21480
rect 3660 21440 4068 21468
rect 3660 21428 3666 21440
rect 4062 21428 4068 21440
rect 4120 21468 4126 21480
rect 4985 21471 5043 21477
rect 4985 21468 4997 21471
rect 4120 21440 4997 21468
rect 4120 21428 4126 21440
rect 4985 21437 4997 21440
rect 5031 21437 5043 21471
rect 4985 21431 5043 21437
rect 7650 21428 7656 21480
rect 7708 21428 7714 21480
rect 8754 21428 8760 21480
rect 8812 21428 8818 21480
rect 8849 21471 8907 21477
rect 8849 21437 8861 21471
rect 8895 21468 8907 21471
rect 9030 21468 9036 21480
rect 8895 21440 9036 21468
rect 8895 21437 8907 21440
rect 8849 21431 8907 21437
rect 9030 21428 9036 21440
rect 9088 21428 9094 21480
rect 10060 21477 10088 21576
rect 12250 21564 12256 21616
rect 12308 21604 12314 21616
rect 12308 21576 17080 21604
rect 12308 21564 12314 21576
rect 12161 21539 12219 21545
rect 12161 21505 12173 21539
rect 12207 21536 12219 21539
rect 13630 21536 13636 21548
rect 12207 21508 13636 21536
rect 12207 21505 12219 21508
rect 12161 21499 12219 21505
rect 13630 21496 13636 21508
rect 13688 21496 13694 21548
rect 15197 21539 15255 21545
rect 15197 21505 15209 21539
rect 15243 21536 15255 21539
rect 16114 21536 16120 21548
rect 15243 21508 16120 21536
rect 15243 21505 15255 21508
rect 15197 21499 15255 21505
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 16206 21496 16212 21548
rect 16264 21496 16270 21548
rect 17052 21545 17080 21576
rect 17218 21564 17224 21616
rect 17276 21604 17282 21616
rect 17678 21604 17684 21616
rect 17276 21576 17684 21604
rect 17276 21564 17282 21576
rect 17678 21564 17684 21576
rect 17736 21564 17742 21616
rect 18708 21545 18736 21644
rect 22554 21632 22560 21684
rect 22612 21632 22618 21684
rect 22002 21564 22008 21616
rect 22060 21604 22066 21616
rect 22060 21576 23428 21604
rect 22060 21564 22066 21576
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21505 17095 21539
rect 17037 21499 17095 21505
rect 18693 21539 18751 21545
rect 18693 21505 18705 21539
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 20162 21496 20168 21548
rect 20220 21536 20226 21548
rect 20438 21536 20444 21548
rect 20220 21508 20444 21536
rect 20220 21496 20226 21508
rect 20438 21496 20444 21508
rect 20496 21496 20502 21548
rect 22465 21539 22523 21545
rect 22465 21505 22477 21539
rect 22511 21536 22523 21539
rect 23290 21536 23296 21548
rect 22511 21508 23296 21536
rect 22511 21505 22523 21508
rect 22465 21499 22523 21505
rect 23290 21496 23296 21508
rect 23348 21496 23354 21548
rect 23400 21545 23428 21576
rect 23658 21564 23664 21616
rect 23716 21564 23722 21616
rect 24210 21564 24216 21616
rect 24268 21564 24274 21616
rect 23385 21539 23443 21545
rect 23385 21505 23397 21539
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 9953 21471 10011 21477
rect 9953 21437 9965 21471
rect 9999 21437 10011 21471
rect 9953 21431 10011 21437
rect 10045 21471 10103 21477
rect 10045 21437 10057 21471
rect 10091 21437 10103 21471
rect 10045 21431 10103 21437
rect 3786 21360 3792 21412
rect 3844 21360 3850 21412
rect 3970 21360 3976 21412
rect 4028 21400 4034 21412
rect 7466 21400 7472 21412
rect 4028 21372 7472 21400
rect 4028 21360 4034 21372
rect 7466 21360 7472 21372
rect 7524 21360 7530 21412
rect 7834 21360 7840 21412
rect 7892 21400 7898 21412
rect 9493 21403 9551 21409
rect 9493 21400 9505 21403
rect 7892 21372 9505 21400
rect 7892 21360 7898 21372
rect 9493 21369 9505 21372
rect 9539 21369 9551 21403
rect 9968 21400 9996 21431
rect 12250 21428 12256 21480
rect 12308 21428 12314 21480
rect 14185 21471 14243 21477
rect 14185 21437 14197 21471
rect 14231 21468 14243 21471
rect 14550 21468 14556 21480
rect 14231 21440 14556 21468
rect 14231 21437 14243 21440
rect 14185 21431 14243 21437
rect 14550 21428 14556 21440
rect 14608 21428 14614 21480
rect 14642 21428 14648 21480
rect 14700 21468 14706 21480
rect 15289 21471 15347 21477
rect 15289 21468 15301 21471
rect 14700 21440 15301 21468
rect 14700 21428 14706 21440
rect 15289 21437 15301 21440
rect 15335 21437 15347 21471
rect 15289 21431 15347 21437
rect 15378 21428 15384 21480
rect 15436 21428 15442 21480
rect 17586 21428 17592 21480
rect 17644 21468 17650 21480
rect 17681 21471 17739 21477
rect 17681 21468 17693 21471
rect 17644 21440 17693 21468
rect 17644 21428 17650 21440
rect 17681 21437 17693 21440
rect 17727 21437 17739 21471
rect 17681 21431 17739 21437
rect 22278 21428 22284 21480
rect 22336 21468 22342 21480
rect 22741 21471 22799 21477
rect 22741 21468 22753 21471
rect 22336 21440 22753 21468
rect 22336 21428 22342 21440
rect 22741 21437 22753 21440
rect 22787 21468 22799 21471
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 22787 21440 25145 21468
rect 22787 21437 22799 21440
rect 22741 21431 22799 21437
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 11054 21400 11060 21412
rect 9968 21372 11060 21400
rect 9493 21363 9551 21369
rect 11054 21360 11060 21372
rect 11112 21360 11118 21412
rect 15930 21400 15936 21412
rect 12406 21372 15936 21400
rect 4801 21335 4859 21341
rect 4801 21301 4813 21335
rect 4847 21332 4859 21335
rect 5810 21332 5816 21344
rect 4847 21304 5816 21332
rect 4847 21301 4859 21304
rect 4801 21295 4859 21301
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 5902 21292 5908 21344
rect 5960 21332 5966 21344
rect 12406 21332 12434 21372
rect 15930 21360 15936 21372
rect 15988 21360 15994 21412
rect 16025 21403 16083 21409
rect 16025 21369 16037 21403
rect 16071 21400 16083 21403
rect 17218 21400 17224 21412
rect 16071 21372 17224 21400
rect 16071 21369 16083 21372
rect 16025 21363 16083 21369
rect 17218 21360 17224 21372
rect 17276 21360 17282 21412
rect 20254 21400 20260 21412
rect 17328 21372 20260 21400
rect 5960 21304 12434 21332
rect 5960 21292 5966 21304
rect 13814 21292 13820 21344
rect 13872 21332 13878 21344
rect 14829 21335 14887 21341
rect 14829 21332 14841 21335
rect 13872 21304 14841 21332
rect 13872 21292 13878 21304
rect 14829 21301 14841 21304
rect 14875 21301 14887 21335
rect 14829 21295 14887 21301
rect 16850 21292 16856 21344
rect 16908 21292 16914 21344
rect 17034 21292 17040 21344
rect 17092 21332 17098 21344
rect 17328 21332 17356 21372
rect 20254 21360 20260 21372
rect 20312 21360 20318 21412
rect 17092 21304 17356 21332
rect 17092 21292 17098 21304
rect 18414 21292 18420 21344
rect 18472 21332 18478 21344
rect 18509 21335 18567 21341
rect 18509 21332 18521 21335
rect 18472 21304 18521 21332
rect 18472 21292 18478 21304
rect 18509 21301 18521 21304
rect 18555 21301 18567 21335
rect 18509 21295 18567 21301
rect 20438 21292 20444 21344
rect 20496 21292 20502 21344
rect 21266 21292 21272 21344
rect 21324 21332 21330 21344
rect 22097 21335 22155 21341
rect 22097 21332 22109 21335
rect 21324 21304 22109 21332
rect 21324 21292 21330 21304
rect 22097 21301 22109 21304
rect 22143 21301 22155 21335
rect 22097 21295 22155 21301
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 2866 21088 2872 21140
rect 2924 21128 2930 21140
rect 3145 21131 3203 21137
rect 3145 21128 3157 21131
rect 2924 21100 3157 21128
rect 2924 21088 2930 21100
rect 3145 21097 3157 21100
rect 3191 21097 3203 21131
rect 3145 21091 3203 21097
rect 7282 21088 7288 21140
rect 7340 21128 7346 21140
rect 7837 21131 7895 21137
rect 7837 21128 7849 21131
rect 7340 21100 7849 21128
rect 7340 21088 7346 21100
rect 7837 21097 7849 21100
rect 7883 21097 7895 21131
rect 7837 21091 7895 21097
rect 10502 21088 10508 21140
rect 10560 21128 10566 21140
rect 11885 21131 11943 21137
rect 11885 21128 11897 21131
rect 10560 21100 11897 21128
rect 10560 21088 10566 21100
rect 11885 21097 11897 21100
rect 11931 21097 11943 21131
rect 11885 21091 11943 21097
rect 13725 21131 13783 21137
rect 13725 21097 13737 21131
rect 13771 21128 13783 21131
rect 14182 21128 14188 21140
rect 13771 21100 14188 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 14182 21088 14188 21100
rect 14240 21088 14246 21140
rect 16850 21088 16856 21140
rect 16908 21128 16914 21140
rect 22005 21131 22063 21137
rect 16908 21100 21220 21128
rect 16908 21088 16914 21100
rect 4065 21063 4123 21069
rect 4065 21029 4077 21063
rect 4111 21029 4123 21063
rect 12250 21060 12256 21072
rect 4065 21023 4123 21029
rect 11532 21032 12256 21060
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20992 2835 20995
rect 4080 20992 4108 21023
rect 2823 20964 4108 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 7742 20952 7748 21004
rect 7800 20992 7806 21004
rect 8481 20995 8539 21001
rect 8481 20992 8493 20995
rect 7800 20964 8493 20992
rect 7800 20952 7806 20964
rect 8481 20961 8493 20964
rect 8527 20992 8539 20995
rect 10410 20992 10416 21004
rect 8527 20964 10416 20992
rect 8527 20961 8539 20964
rect 8481 20955 8539 20961
rect 10410 20952 10416 20964
rect 10468 20992 10474 21004
rect 11532 21001 11560 21032
rect 12250 21020 12256 21032
rect 12308 21020 12314 21072
rect 12342 21020 12348 21072
rect 12400 21060 12406 21072
rect 16206 21060 16212 21072
rect 12400 21032 16212 21060
rect 12400 21020 12406 21032
rect 16206 21020 16212 21032
rect 16264 21020 16270 21072
rect 16301 21063 16359 21069
rect 16301 21029 16313 21063
rect 16347 21060 16359 21063
rect 17034 21060 17040 21072
rect 16347 21032 17040 21060
rect 16347 21029 16359 21032
rect 16301 21023 16359 21029
rect 11517 20995 11575 21001
rect 11517 20992 11529 20995
rect 10468 20964 11529 20992
rect 10468 20952 10474 20964
rect 11517 20961 11529 20964
rect 11563 20961 11575 20995
rect 13817 20995 13875 21001
rect 13817 20992 13829 20995
rect 11517 20955 11575 20961
rect 12268 20964 13829 20992
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20893 2283 20927
rect 2225 20887 2283 20893
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20924 3019 20927
rect 3694 20924 3700 20936
rect 3007 20896 3700 20924
rect 3007 20893 3019 20896
rect 2961 20887 3019 20893
rect 1854 20816 1860 20868
rect 1912 20856 1918 20868
rect 2240 20856 2268 20887
rect 3694 20884 3700 20896
rect 3752 20924 3758 20936
rect 4062 20924 4068 20936
rect 3752 20896 4068 20924
rect 3752 20884 3758 20896
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 4246 20884 4252 20936
rect 4304 20884 4310 20936
rect 9769 20927 9827 20933
rect 9769 20893 9781 20927
rect 9815 20893 9827 20927
rect 9769 20887 9827 20893
rect 2866 20856 2872 20868
rect 1912 20828 2176 20856
rect 2240 20828 2872 20856
rect 1912 20816 1918 20828
rect 1762 20748 1768 20800
rect 1820 20788 1826 20800
rect 2041 20791 2099 20797
rect 2041 20788 2053 20791
rect 1820 20760 2053 20788
rect 1820 20748 1826 20760
rect 2041 20757 2053 20760
rect 2087 20757 2099 20791
rect 2148 20788 2176 20828
rect 2866 20816 2872 20828
rect 2924 20816 2930 20868
rect 7742 20816 7748 20868
rect 7800 20856 7806 20868
rect 8297 20859 8355 20865
rect 8297 20856 8309 20859
rect 7800 20828 8309 20856
rect 7800 20816 7806 20828
rect 8297 20825 8309 20828
rect 8343 20825 8355 20859
rect 9784 20856 9812 20887
rect 11882 20884 11888 20936
rect 11940 20924 11946 20936
rect 12268 20924 12296 20964
rect 13817 20961 13829 20964
rect 13863 20992 13875 20995
rect 14921 20995 14979 21001
rect 14921 20992 14933 20995
rect 13863 20964 14933 20992
rect 13863 20961 13875 20964
rect 13817 20955 13875 20961
rect 14921 20961 14933 20964
rect 14967 20961 14979 20995
rect 16316 20992 16344 21023
rect 17034 21020 17040 21032
rect 17092 21020 17098 21072
rect 17221 21063 17279 21069
rect 17221 21029 17233 21063
rect 17267 21060 17279 21063
rect 19334 21060 19340 21072
rect 17267 21032 19340 21060
rect 17267 21029 17279 21032
rect 17221 21023 17279 21029
rect 19334 21020 19340 21032
rect 19392 21020 19398 21072
rect 21192 21060 21220 21100
rect 22005 21097 22017 21131
rect 22051 21128 22063 21131
rect 22370 21128 22376 21140
rect 22051 21100 22376 21128
rect 22051 21097 22063 21100
rect 22005 21091 22063 21097
rect 22370 21088 22376 21100
rect 22428 21128 22434 21140
rect 24210 21128 24216 21140
rect 22428 21100 24216 21128
rect 22428 21088 22434 21100
rect 24210 21088 24216 21100
rect 24268 21088 24274 21140
rect 23474 21060 23480 21072
rect 21192 21032 23480 21060
rect 23474 21020 23480 21032
rect 23532 21020 23538 21072
rect 14921 20955 14979 20961
rect 15672 20964 16344 20992
rect 11940 20896 12296 20924
rect 11940 20884 11946 20896
rect 12342 20884 12348 20936
rect 12400 20924 12406 20936
rect 12618 20924 12624 20936
rect 12400 20896 12624 20924
rect 12400 20884 12406 20896
rect 12618 20884 12624 20896
rect 12676 20884 12682 20936
rect 14182 20884 14188 20936
rect 14240 20924 14246 20936
rect 14829 20927 14887 20933
rect 14829 20924 14841 20927
rect 14240 20896 14841 20924
rect 14240 20884 14246 20896
rect 14829 20893 14841 20896
rect 14875 20893 14887 20927
rect 15672 20924 15700 20964
rect 17310 20952 17316 21004
rect 17368 20992 17374 21004
rect 17865 20995 17923 21001
rect 17368 20964 17724 20992
rect 17368 20952 17374 20964
rect 14829 20887 14887 20893
rect 15120 20896 15700 20924
rect 9950 20856 9956 20868
rect 9784 20828 9956 20856
rect 8297 20819 8355 20825
rect 9950 20816 9956 20828
rect 10008 20816 10014 20868
rect 10045 20859 10103 20865
rect 10045 20825 10057 20859
rect 10091 20856 10103 20859
rect 10318 20856 10324 20868
rect 10091 20828 10324 20856
rect 10091 20825 10103 20828
rect 10045 20819 10103 20825
rect 10318 20816 10324 20828
rect 10376 20816 10382 20868
rect 10502 20856 10508 20868
rect 10428 20828 10508 20856
rect 7469 20791 7527 20797
rect 7469 20788 7481 20791
rect 2148 20760 7481 20788
rect 2041 20751 2099 20757
rect 7469 20757 7481 20760
rect 7515 20788 7527 20791
rect 8205 20791 8263 20797
rect 8205 20788 8217 20791
rect 7515 20760 8217 20788
rect 7515 20757 7527 20760
rect 7469 20751 7527 20757
rect 8205 20757 8217 20760
rect 8251 20788 8263 20791
rect 8570 20788 8576 20800
rect 8251 20760 8576 20788
rect 8251 20757 8263 20760
rect 8205 20751 8263 20757
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 9582 20748 9588 20800
rect 9640 20788 9646 20800
rect 10428 20788 10456 20828
rect 10502 20816 10508 20828
rect 10560 20816 10566 20868
rect 11348 20828 12388 20856
rect 9640 20760 10456 20788
rect 9640 20748 9646 20760
rect 10686 20748 10692 20800
rect 10744 20788 10750 20800
rect 11348 20788 11376 20828
rect 10744 20760 11376 20788
rect 12360 20788 12388 20828
rect 14200 20788 14228 20884
rect 14737 20859 14795 20865
rect 14737 20825 14749 20859
rect 14783 20856 14795 20859
rect 15120 20856 15148 20896
rect 15746 20884 15752 20936
rect 15804 20884 15810 20936
rect 16114 20884 16120 20936
rect 16172 20924 16178 20936
rect 16172 20896 17540 20924
rect 16172 20884 16178 20896
rect 14783 20828 15148 20856
rect 14783 20825 14795 20828
rect 14737 20819 14795 20825
rect 15194 20816 15200 20868
rect 15252 20856 15258 20868
rect 16942 20856 16948 20868
rect 15252 20828 16948 20856
rect 15252 20816 15258 20828
rect 16942 20816 16948 20828
rect 17000 20816 17006 20868
rect 17512 20856 17540 20896
rect 17586 20884 17592 20936
rect 17644 20884 17650 20936
rect 17696 20924 17724 20964
rect 17865 20961 17877 20995
rect 17911 20992 17923 20995
rect 17911 20964 19380 20992
rect 17911 20961 17923 20964
rect 17865 20955 17923 20961
rect 18877 20927 18935 20933
rect 18877 20924 18889 20927
rect 17696 20896 18889 20924
rect 18877 20893 18889 20896
rect 18923 20893 18935 20927
rect 18877 20887 18935 20893
rect 19150 20856 19156 20868
rect 17512 20828 19156 20856
rect 19150 20816 19156 20828
rect 19208 20816 19214 20868
rect 19352 20856 19380 20964
rect 19426 20952 19432 21004
rect 19484 20992 19490 21004
rect 19889 20995 19947 21001
rect 19889 20992 19901 20995
rect 19484 20964 19901 20992
rect 19484 20952 19490 20964
rect 19889 20961 19901 20964
rect 19935 20961 19947 20995
rect 19889 20955 19947 20961
rect 23845 20995 23903 21001
rect 23845 20961 23857 20995
rect 23891 20992 23903 20995
rect 24854 20992 24860 21004
rect 23891 20964 24860 20992
rect 23891 20961 23903 20964
rect 23845 20955 23903 20961
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 22370 20924 22376 20936
rect 21298 20896 22376 20924
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 22646 20884 22652 20936
rect 22704 20884 22710 20936
rect 20162 20856 20168 20868
rect 19352 20828 20168 20856
rect 20162 20816 20168 20828
rect 20220 20816 20226 20868
rect 25038 20856 25044 20868
rect 21468 20828 25044 20856
rect 12360 20760 14228 20788
rect 10744 20748 10750 20760
rect 14274 20748 14280 20800
rect 14332 20788 14338 20800
rect 14369 20791 14427 20797
rect 14369 20788 14381 20791
rect 14332 20760 14381 20788
rect 14332 20748 14338 20760
rect 14369 20757 14381 20760
rect 14415 20757 14427 20791
rect 14369 20751 14427 20757
rect 15565 20791 15623 20797
rect 15565 20757 15577 20791
rect 15611 20788 15623 20791
rect 15654 20788 15660 20800
rect 15611 20760 15660 20788
rect 15611 20757 15623 20760
rect 15565 20751 15623 20757
rect 15654 20748 15660 20760
rect 15712 20748 15718 20800
rect 16850 20748 16856 20800
rect 16908 20788 16914 20800
rect 17681 20791 17739 20797
rect 17681 20788 17693 20791
rect 16908 20760 17693 20788
rect 16908 20748 16914 20760
rect 17681 20757 17693 20760
rect 17727 20757 17739 20791
rect 17681 20751 17739 20757
rect 18693 20791 18751 20797
rect 18693 20757 18705 20791
rect 18739 20788 18751 20791
rect 21468 20788 21496 20828
rect 25038 20816 25044 20828
rect 25096 20816 25102 20868
rect 18739 20760 21496 20788
rect 18739 20757 18751 20760
rect 18693 20751 18751 20757
rect 21634 20748 21640 20800
rect 21692 20748 21698 20800
rect 22370 20748 22376 20800
rect 22428 20748 22434 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 5718 20584 5724 20596
rect 3988 20556 5724 20584
rect 3988 20457 4016 20556
rect 5718 20544 5724 20556
rect 5776 20544 5782 20596
rect 8846 20584 8852 20596
rect 6656 20556 8852 20584
rect 4249 20519 4307 20525
rect 4249 20485 4261 20519
rect 4295 20516 4307 20519
rect 4338 20516 4344 20528
rect 4295 20488 4344 20516
rect 4295 20485 4307 20488
rect 4249 20479 4307 20485
rect 4338 20476 4344 20488
rect 4396 20476 4402 20528
rect 5997 20519 6055 20525
rect 5997 20516 6009 20519
rect 5474 20488 6009 20516
rect 5997 20485 6009 20488
rect 6043 20516 6055 20519
rect 6454 20516 6460 20528
rect 6043 20488 6460 20516
rect 6043 20485 6055 20488
rect 5997 20479 6055 20485
rect 6454 20476 6460 20488
rect 6512 20476 6518 20528
rect 6656 20516 6684 20556
rect 8846 20544 8852 20556
rect 8904 20544 8910 20596
rect 8938 20544 8944 20596
rect 8996 20584 9002 20596
rect 9953 20587 10011 20593
rect 9953 20584 9965 20587
rect 8996 20556 9965 20584
rect 8996 20544 9002 20556
rect 9953 20553 9965 20556
rect 9999 20553 10011 20587
rect 9953 20547 10011 20553
rect 12437 20587 12495 20593
rect 12437 20553 12449 20587
rect 12483 20584 12495 20587
rect 13265 20587 13323 20593
rect 13265 20584 13277 20587
rect 12483 20556 13277 20584
rect 12483 20553 12495 20556
rect 12437 20547 12495 20553
rect 13265 20553 13277 20556
rect 13311 20553 13323 20587
rect 13265 20547 13323 20553
rect 17310 20544 17316 20596
rect 17368 20584 17374 20596
rect 17368 20556 17724 20584
rect 17368 20544 17374 20556
rect 6564 20488 6684 20516
rect 3973 20451 4031 20457
rect 3973 20417 3985 20451
rect 4019 20417 4031 20451
rect 3973 20411 4031 20417
rect 5718 20408 5724 20460
rect 5776 20448 5782 20460
rect 6564 20457 6592 20488
rect 7282 20476 7288 20528
rect 7340 20476 7346 20528
rect 9030 20476 9036 20528
rect 9088 20516 9094 20528
rect 10413 20519 10471 20525
rect 9088 20488 9628 20516
rect 9088 20476 9094 20488
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 5776 20420 6561 20448
rect 5776 20408 5782 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 8662 20408 8668 20460
rect 8720 20448 8726 20460
rect 9125 20451 9183 20457
rect 9125 20448 9137 20451
rect 8720 20420 9137 20448
rect 8720 20408 8726 20420
rect 9125 20417 9137 20420
rect 9171 20417 9183 20451
rect 9125 20411 9183 20417
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 9217 20383 9275 20389
rect 6871 20352 9168 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 8754 20272 8760 20324
rect 8812 20272 8818 20324
rect 9140 20312 9168 20352
rect 9217 20349 9229 20383
rect 9263 20380 9275 20383
rect 9306 20380 9312 20392
rect 9263 20352 9312 20380
rect 9263 20349 9275 20352
rect 9217 20343 9275 20349
rect 9306 20340 9312 20352
rect 9364 20340 9370 20392
rect 9401 20383 9459 20389
rect 9401 20349 9413 20383
rect 9447 20349 9459 20383
rect 9600 20380 9628 20488
rect 10413 20485 10425 20519
rect 10459 20516 10471 20519
rect 11514 20516 11520 20528
rect 10459 20488 11520 20516
rect 10459 20485 10471 20488
rect 10413 20479 10471 20485
rect 11514 20476 11520 20488
rect 11572 20476 11578 20528
rect 16850 20516 16856 20528
rect 12406 20488 16856 20516
rect 10321 20451 10379 20457
rect 10321 20417 10333 20451
rect 10367 20448 10379 20451
rect 11698 20448 11704 20460
rect 10367 20420 11704 20448
rect 10367 20417 10379 20420
rect 10321 20411 10379 20417
rect 11698 20408 11704 20420
rect 11756 20408 11762 20460
rect 10505 20383 10563 20389
rect 10505 20380 10517 20383
rect 9600 20352 10517 20380
rect 9401 20343 9459 20349
rect 10505 20349 10517 20352
rect 10551 20349 10563 20383
rect 10505 20343 10563 20349
rect 9416 20312 9444 20343
rect 10594 20340 10600 20392
rect 10652 20380 10658 20392
rect 12406 20380 12434 20488
rect 16850 20476 16856 20488
rect 16908 20476 16914 20528
rect 17696 20525 17724 20556
rect 19334 20544 19340 20596
rect 19392 20544 19398 20596
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 19518 20584 19524 20596
rect 19475 20556 19524 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 17681 20519 17739 20525
rect 17681 20485 17693 20519
rect 17727 20485 17739 20519
rect 17681 20479 17739 20485
rect 17954 20476 17960 20528
rect 18012 20516 18018 20528
rect 18598 20516 18604 20528
rect 18012 20488 18604 20516
rect 18012 20476 18018 20488
rect 18598 20476 18604 20488
rect 18656 20516 18662 20528
rect 19610 20516 19616 20528
rect 18656 20488 19616 20516
rect 18656 20476 18662 20488
rect 19610 20476 19616 20488
rect 19668 20476 19674 20528
rect 23293 20519 23351 20525
rect 23293 20485 23305 20519
rect 23339 20516 23351 20519
rect 23382 20516 23388 20528
rect 23339 20488 23388 20516
rect 23339 20485 23351 20488
rect 23293 20479 23351 20485
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 25130 20516 25136 20528
rect 23584 20488 25136 20516
rect 13446 20408 13452 20460
rect 13504 20448 13510 20460
rect 15657 20451 15715 20457
rect 15657 20448 15669 20451
rect 13504 20420 15669 20448
rect 13504 20408 13510 20420
rect 15657 20417 15669 20420
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 18506 20408 18512 20460
rect 18564 20408 18570 20460
rect 22281 20451 22339 20457
rect 22281 20417 22293 20451
rect 22327 20448 22339 20451
rect 23584 20448 23612 20488
rect 25130 20476 25136 20488
rect 25188 20476 25194 20528
rect 22327 20420 23612 20448
rect 24121 20451 24179 20457
rect 22327 20417 22339 20420
rect 22281 20411 22339 20417
rect 24121 20417 24133 20451
rect 24167 20448 24179 20451
rect 25222 20448 25228 20460
rect 24167 20420 25228 20448
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 25222 20408 25228 20420
rect 25280 20408 25286 20460
rect 10652 20352 12434 20380
rect 12529 20383 12587 20389
rect 10652 20340 10658 20352
rect 12529 20349 12541 20383
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 11606 20312 11612 20324
rect 9140 20284 11612 20312
rect 11606 20272 11612 20284
rect 11664 20272 11670 20324
rect 5721 20247 5779 20253
rect 5721 20213 5733 20247
rect 5767 20244 5779 20247
rect 5810 20244 5816 20256
rect 5767 20216 5816 20244
rect 5767 20213 5779 20216
rect 5721 20207 5779 20213
rect 5810 20204 5816 20216
rect 5868 20204 5874 20256
rect 6454 20204 6460 20256
rect 6512 20244 6518 20256
rect 7282 20244 7288 20256
rect 6512 20216 7288 20244
rect 6512 20204 6518 20216
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 9030 20244 9036 20256
rect 8352 20216 9036 20244
rect 8352 20204 8358 20216
rect 9030 20204 9036 20216
rect 9088 20204 9094 20256
rect 12066 20204 12072 20256
rect 12124 20204 12130 20256
rect 12544 20244 12572 20343
rect 12710 20340 12716 20392
rect 12768 20340 12774 20392
rect 19613 20383 19671 20389
rect 19613 20349 19625 20383
rect 19659 20380 19671 20383
rect 21634 20380 21640 20392
rect 19659 20352 21640 20380
rect 19659 20349 19671 20352
rect 19613 20343 19671 20349
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 24670 20340 24676 20392
rect 24728 20340 24734 20392
rect 17862 20272 17868 20324
rect 17920 20272 17926 20324
rect 13354 20244 13360 20256
rect 12544 20216 13360 20244
rect 13354 20204 13360 20216
rect 13412 20244 13418 20256
rect 13725 20247 13783 20253
rect 13725 20244 13737 20247
rect 13412 20216 13737 20244
rect 13412 20204 13418 20216
rect 13725 20213 13737 20216
rect 13771 20244 13783 20247
rect 13998 20244 14004 20256
rect 13771 20216 14004 20244
rect 13771 20213 13783 20216
rect 13725 20207 13783 20213
rect 13998 20204 14004 20216
rect 14056 20204 14062 20256
rect 14090 20204 14096 20256
rect 14148 20244 14154 20256
rect 14642 20244 14648 20256
rect 14148 20216 14648 20244
rect 14148 20204 14154 20216
rect 14642 20204 14648 20216
rect 14700 20204 14706 20256
rect 15473 20247 15531 20253
rect 15473 20213 15485 20247
rect 15519 20244 15531 20247
rect 17310 20244 17316 20256
rect 15519 20216 17316 20244
rect 15519 20213 15531 20216
rect 15473 20207 15531 20213
rect 17310 20204 17316 20216
rect 17368 20204 17374 20256
rect 18325 20247 18383 20253
rect 18325 20213 18337 20247
rect 18371 20244 18383 20247
rect 18782 20244 18788 20256
rect 18371 20216 18788 20244
rect 18371 20213 18383 20216
rect 18325 20207 18383 20213
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 18969 20247 19027 20253
rect 18969 20213 18981 20247
rect 19015 20244 19027 20247
rect 19794 20244 19800 20256
rect 19015 20216 19800 20244
rect 19015 20213 19027 20216
rect 18969 20207 19027 20213
rect 19794 20204 19800 20216
rect 19852 20204 19858 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 5074 20000 5080 20052
rect 5132 20000 5138 20052
rect 11698 20000 11704 20052
rect 11756 20000 11762 20052
rect 13630 20000 13636 20052
rect 13688 20040 13694 20052
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 13688 20012 14289 20040
rect 13688 20000 13694 20012
rect 14277 20009 14289 20012
rect 14323 20009 14335 20043
rect 14277 20003 14335 20009
rect 20349 20043 20407 20049
rect 20349 20009 20361 20043
rect 20395 20040 20407 20043
rect 20530 20040 20536 20052
rect 20395 20012 20536 20040
rect 20395 20009 20407 20012
rect 20349 20003 20407 20009
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 12158 19972 12164 19984
rect 11164 19944 12164 19972
rect 5718 19864 5724 19916
rect 5776 19864 5782 19916
rect 5997 19907 6055 19913
rect 5997 19873 6009 19907
rect 6043 19904 6055 19907
rect 8294 19904 8300 19916
rect 6043 19876 8300 19904
rect 6043 19873 6055 19876
rect 5997 19867 6055 19873
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 8846 19864 8852 19916
rect 8904 19904 8910 19916
rect 11164 19913 11192 19944
rect 12158 19932 12164 19944
rect 12216 19932 12222 19984
rect 14642 19932 14648 19984
rect 14700 19972 14706 19984
rect 15381 19975 15439 19981
rect 15381 19972 15393 19975
rect 14700 19944 15393 19972
rect 14700 19932 14706 19944
rect 15381 19941 15393 19944
rect 15427 19972 15439 19975
rect 17954 19972 17960 19984
rect 15427 19944 17960 19972
rect 15427 19941 15439 19944
rect 15381 19935 15439 19941
rect 17954 19932 17960 19944
rect 18012 19932 18018 19984
rect 9125 19907 9183 19913
rect 9125 19904 9137 19907
rect 8904 19876 9137 19904
rect 8904 19864 8910 19876
rect 9125 19873 9137 19876
rect 9171 19873 9183 19907
rect 9125 19867 9183 19873
rect 11149 19907 11207 19913
rect 11149 19873 11161 19907
rect 11195 19873 11207 19907
rect 12253 19907 12311 19913
rect 12253 19904 12265 19907
rect 11149 19867 11207 19873
rect 11900 19876 12265 19904
rect 5261 19839 5319 19845
rect 5261 19805 5273 19839
rect 5307 19805 5319 19839
rect 5261 19799 5319 19805
rect 5276 19700 5304 19799
rect 7282 19796 7288 19848
rect 7340 19836 7346 19848
rect 7745 19839 7803 19845
rect 7745 19836 7757 19839
rect 7340 19808 7757 19836
rect 7340 19796 7346 19808
rect 7745 19805 7757 19808
rect 7791 19836 7803 19839
rect 8389 19839 8447 19845
rect 8389 19836 8401 19839
rect 7791 19808 8401 19836
rect 7791 19805 7803 19808
rect 7745 19799 7803 19805
rect 8389 19805 8401 19808
rect 8435 19836 8447 19839
rect 8938 19836 8944 19848
rect 8435 19808 8944 19836
rect 8435 19805 8447 19808
rect 8389 19799 8447 19805
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 11606 19796 11612 19848
rect 11664 19836 11670 19848
rect 11900 19836 11928 19876
rect 12253 19873 12265 19876
rect 12299 19873 12311 19907
rect 12253 19867 12311 19873
rect 14458 19864 14464 19916
rect 14516 19904 14522 19916
rect 14829 19907 14887 19913
rect 14829 19904 14841 19907
rect 14516 19876 14841 19904
rect 14516 19864 14522 19876
rect 14829 19873 14841 19876
rect 14875 19873 14887 19907
rect 14829 19867 14887 19873
rect 17402 19864 17408 19916
rect 17460 19904 17466 19916
rect 23845 19907 23903 19913
rect 17460 19876 22048 19904
rect 17460 19864 17466 19876
rect 11664 19808 11928 19836
rect 12069 19839 12127 19845
rect 11664 19796 11670 19808
rect 12069 19805 12081 19839
rect 12115 19836 12127 19839
rect 12434 19836 12440 19848
rect 12115 19808 12440 19836
rect 12115 19805 12127 19808
rect 12069 19799 12127 19805
rect 12434 19796 12440 19808
rect 12492 19796 12498 19848
rect 13909 19839 13967 19845
rect 13909 19805 13921 19839
rect 13955 19836 13967 19839
rect 17221 19839 17279 19845
rect 13955 19808 14780 19836
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 6454 19728 6460 19780
rect 6512 19728 6518 19780
rect 7650 19768 7656 19780
rect 7484 19740 7656 19768
rect 7374 19700 7380 19712
rect 5276 19672 7380 19700
rect 7374 19660 7380 19672
rect 7432 19660 7438 19712
rect 7484 19709 7512 19740
rect 7650 19728 7656 19740
rect 7708 19768 7714 19780
rect 9401 19771 9459 19777
rect 9401 19768 9413 19771
rect 7708 19740 9413 19768
rect 7708 19728 7714 19740
rect 9401 19737 9413 19740
rect 9447 19737 9459 19771
rect 12161 19771 12219 19777
rect 9401 19731 9459 19737
rect 9508 19740 9890 19768
rect 7469 19703 7527 19709
rect 7469 19669 7481 19703
rect 7515 19669 7527 19703
rect 7469 19663 7527 19669
rect 8662 19660 8668 19712
rect 8720 19660 8726 19712
rect 8938 19660 8944 19712
rect 8996 19700 9002 19712
rect 9508 19700 9536 19740
rect 12161 19737 12173 19771
rect 12207 19768 12219 19771
rect 14182 19768 14188 19780
rect 12207 19740 14188 19768
rect 12207 19737 12219 19740
rect 12161 19731 12219 19737
rect 14182 19728 14188 19740
rect 14240 19728 14246 19780
rect 14642 19728 14648 19780
rect 14700 19728 14706 19780
rect 14752 19768 14780 19808
rect 17221 19805 17233 19839
rect 17267 19836 17279 19839
rect 17770 19836 17776 19848
rect 17267 19808 17776 19836
rect 17267 19805 17279 19808
rect 17221 19799 17279 19805
rect 17770 19796 17776 19808
rect 17828 19796 17834 19848
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19836 18751 19839
rect 18874 19836 18880 19848
rect 18739 19808 18880 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 18874 19796 18880 19808
rect 18932 19796 18938 19848
rect 22020 19845 22048 19876
rect 23845 19873 23857 19907
rect 23891 19904 23903 19907
rect 24946 19904 24952 19916
rect 23891 19876 24952 19904
rect 23891 19873 23903 19876
rect 23845 19867 23903 19873
rect 24946 19864 24952 19876
rect 25004 19864 25010 19916
rect 22005 19839 22063 19845
rect 22005 19805 22017 19839
rect 22051 19805 22063 19839
rect 22005 19799 22063 19805
rect 22833 19839 22891 19845
rect 22833 19805 22845 19839
rect 22879 19836 22891 19839
rect 25590 19836 25596 19848
rect 22879 19808 25596 19836
rect 22879 19805 22891 19808
rect 22833 19799 22891 19805
rect 25590 19796 25596 19808
rect 25648 19796 25654 19848
rect 17313 19771 17371 19777
rect 17313 19768 17325 19771
rect 14752 19740 17325 19768
rect 14752 19712 14780 19740
rect 17313 19737 17325 19740
rect 17359 19768 17371 19771
rect 17586 19768 17592 19780
rect 17359 19740 17592 19768
rect 17359 19737 17371 19740
rect 17313 19731 17371 19737
rect 17586 19728 17592 19740
rect 17644 19728 17650 19780
rect 17957 19771 18015 19777
rect 17957 19737 17969 19771
rect 18003 19768 18015 19771
rect 18414 19768 18420 19780
rect 18003 19740 18420 19768
rect 18003 19737 18015 19740
rect 17957 19731 18015 19737
rect 18414 19728 18420 19740
rect 18472 19728 18478 19780
rect 22189 19771 22247 19777
rect 22189 19737 22201 19771
rect 22235 19768 22247 19771
rect 23842 19768 23848 19780
rect 22235 19740 23848 19768
rect 22235 19737 22247 19740
rect 22189 19731 22247 19737
rect 23842 19728 23848 19740
rect 23900 19728 23906 19780
rect 9582 19700 9588 19712
rect 8996 19672 9588 19700
rect 8996 19660 9002 19672
rect 9582 19660 9588 19672
rect 9640 19660 9646 19712
rect 14734 19660 14740 19712
rect 14792 19660 14798 19712
rect 18509 19703 18567 19709
rect 18509 19669 18521 19703
rect 18555 19700 18567 19703
rect 19058 19700 19064 19712
rect 18555 19672 19064 19700
rect 18555 19669 18567 19672
rect 18509 19663 18567 19669
rect 19058 19660 19064 19672
rect 19116 19660 19122 19712
rect 19334 19660 19340 19712
rect 19392 19660 19398 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 1486 19456 1492 19508
rect 1544 19496 1550 19508
rect 2041 19499 2099 19505
rect 2041 19496 2053 19499
rect 1544 19468 2053 19496
rect 1544 19456 1550 19468
rect 2041 19465 2053 19468
rect 2087 19465 2099 19499
rect 3602 19496 3608 19508
rect 2041 19459 2099 19465
rect 2746 19468 3608 19496
rect 2746 19428 2774 19468
rect 3602 19456 3608 19468
rect 3660 19456 3666 19508
rect 4430 19456 4436 19508
rect 4488 19496 4494 19508
rect 4709 19499 4767 19505
rect 4709 19496 4721 19499
rect 4488 19468 4721 19496
rect 4488 19456 4494 19468
rect 4709 19465 4721 19468
rect 4755 19465 4767 19499
rect 4709 19459 4767 19465
rect 9217 19499 9275 19505
rect 9217 19465 9229 19499
rect 9263 19496 9275 19499
rect 9398 19496 9404 19508
rect 9263 19468 9404 19496
rect 9263 19465 9275 19468
rect 9217 19459 9275 19465
rect 9398 19456 9404 19468
rect 9456 19456 9462 19508
rect 11701 19499 11759 19505
rect 11701 19465 11713 19499
rect 11747 19465 11759 19499
rect 11701 19459 11759 19465
rect 12069 19499 12127 19505
rect 12069 19465 12081 19499
rect 12115 19496 12127 19499
rect 13446 19496 13452 19508
rect 12115 19468 13452 19496
rect 12115 19465 12127 19468
rect 12069 19459 12127 19465
rect 4522 19428 4528 19440
rect 2240 19400 2774 19428
rect 3068 19400 4528 19428
rect 2240 19369 2268 19400
rect 3068 19369 3096 19400
rect 4522 19388 4528 19400
rect 4580 19388 4586 19440
rect 7282 19388 7288 19440
rect 7340 19388 7346 19440
rect 9306 19388 9312 19440
rect 9364 19428 9370 19440
rect 11716 19428 11744 19459
rect 13446 19456 13452 19468
rect 13504 19456 13510 19508
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 17497 19499 17555 19505
rect 17497 19465 17509 19499
rect 17543 19496 17555 19499
rect 18690 19496 18696 19508
rect 17543 19468 18696 19496
rect 17543 19465 17555 19468
rect 17497 19459 17555 19465
rect 9364 19400 11744 19428
rect 9364 19388 9370 19400
rect 13998 19388 14004 19440
rect 14056 19428 14062 19440
rect 16298 19428 16304 19440
rect 14056 19400 16304 19428
rect 14056 19388 14062 19400
rect 16298 19388 16304 19400
rect 16356 19388 16362 19440
rect 16868 19428 16896 19459
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 19429 19499 19487 19505
rect 19429 19465 19441 19499
rect 19475 19465 19487 19499
rect 19429 19459 19487 19465
rect 18785 19431 18843 19437
rect 16868 19400 18736 19428
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19329 2283 19363
rect 2225 19323 2283 19329
rect 3053 19363 3111 19369
rect 3053 19329 3065 19363
rect 3099 19329 3111 19363
rect 3053 19323 3111 19329
rect 3878 19320 3884 19372
rect 3936 19320 3942 19372
rect 4893 19363 4951 19369
rect 4893 19329 4905 19363
rect 4939 19360 4951 19363
rect 6270 19360 6276 19372
rect 4939 19332 6276 19360
rect 4939 19329 4951 19332
rect 4893 19323 4951 19329
rect 6270 19320 6276 19332
rect 6328 19320 6334 19372
rect 6546 19320 6552 19372
rect 6604 19320 6610 19372
rect 8386 19320 8392 19372
rect 8444 19360 8450 19372
rect 8662 19360 8668 19372
rect 8444 19332 8668 19360
rect 8444 19320 8450 19332
rect 8662 19320 8668 19332
rect 8720 19360 8726 19372
rect 9125 19363 9183 19369
rect 9125 19360 9137 19363
rect 8720 19332 9137 19360
rect 8720 19320 8726 19332
rect 9125 19329 9137 19332
rect 9171 19329 9183 19363
rect 9125 19323 9183 19329
rect 12158 19320 12164 19372
rect 12216 19320 12222 19372
rect 13909 19363 13967 19369
rect 13909 19329 13921 19363
rect 13955 19360 13967 19363
rect 14642 19360 14648 19372
rect 13955 19332 14648 19360
rect 13955 19329 13967 19332
rect 13909 19323 13967 19329
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 14826 19320 14832 19372
rect 14884 19360 14890 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 14884 19332 17049 19360
rect 14884 19320 14890 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 17586 19320 17592 19372
rect 17644 19360 17650 19372
rect 17865 19363 17923 19369
rect 17865 19360 17877 19363
rect 17644 19332 17877 19360
rect 17644 19320 17650 19332
rect 17865 19329 17877 19332
rect 17911 19329 17923 19363
rect 18708 19360 18736 19400
rect 18785 19397 18797 19431
rect 18831 19428 18843 19431
rect 19242 19428 19248 19440
rect 18831 19400 19248 19428
rect 18831 19397 18843 19400
rect 18785 19391 18843 19397
rect 19242 19388 19248 19400
rect 19300 19388 19306 19440
rect 19444 19428 19472 19459
rect 19518 19456 19524 19508
rect 19576 19496 19582 19508
rect 19797 19499 19855 19505
rect 19797 19496 19809 19499
rect 19576 19468 19809 19496
rect 19576 19456 19582 19468
rect 19797 19465 19809 19468
rect 19843 19465 19855 19499
rect 19797 19459 19855 19465
rect 19889 19499 19947 19505
rect 19889 19465 19901 19499
rect 19935 19496 19947 19499
rect 20530 19496 20536 19508
rect 19935 19468 20536 19496
rect 19935 19465 19947 19468
rect 19889 19459 19947 19465
rect 20530 19456 20536 19468
rect 20588 19456 20594 19508
rect 20717 19499 20775 19505
rect 20717 19465 20729 19499
rect 20763 19465 20775 19499
rect 20717 19459 20775 19465
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 21358 19496 21364 19508
rect 21223 19468 21364 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 20732 19428 20760 19459
rect 21358 19456 21364 19468
rect 21416 19456 21422 19508
rect 21910 19456 21916 19508
rect 21968 19496 21974 19508
rect 23753 19499 23811 19505
rect 23753 19496 23765 19499
rect 21968 19468 23765 19496
rect 21968 19456 21974 19468
rect 23753 19465 23765 19468
rect 23799 19465 23811 19499
rect 23753 19459 23811 19465
rect 22554 19428 22560 19440
rect 19444 19400 20668 19428
rect 20732 19400 22560 19428
rect 20640 19360 20668 19400
rect 22554 19388 22560 19400
rect 22612 19388 22618 19440
rect 20806 19360 20812 19372
rect 18708 19332 19748 19360
rect 20640 19332 20812 19360
rect 17865 19323 17923 19329
rect 6822 19252 6828 19304
rect 6880 19252 6886 19304
rect 9030 19252 9036 19304
rect 9088 19292 9094 19304
rect 9309 19295 9367 19301
rect 9309 19292 9321 19295
rect 9088 19264 9321 19292
rect 9088 19252 9094 19264
rect 9309 19261 9321 19264
rect 9355 19261 9367 19295
rect 9309 19255 9367 19261
rect 9582 19252 9588 19304
rect 9640 19292 9646 19304
rect 11149 19295 11207 19301
rect 11149 19292 11161 19295
rect 9640 19264 11161 19292
rect 9640 19252 9646 19264
rect 11149 19261 11161 19264
rect 11195 19292 11207 19295
rect 12253 19295 12311 19301
rect 12253 19292 12265 19295
rect 11195 19264 12265 19292
rect 11195 19261 11207 19264
rect 11149 19255 11207 19261
rect 12253 19261 12265 19264
rect 12299 19292 12311 19295
rect 12342 19292 12348 19304
rect 12299 19264 12348 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12342 19252 12348 19264
rect 12400 19292 12406 19304
rect 13265 19295 13323 19301
rect 12400 19252 12434 19292
rect 13265 19261 13277 19295
rect 13311 19292 13323 19295
rect 13998 19292 14004 19304
rect 13311 19264 14004 19292
rect 13311 19261 13323 19264
rect 13265 19255 13323 19261
rect 13998 19252 14004 19264
rect 14056 19252 14062 19304
rect 14185 19295 14243 19301
rect 14185 19261 14197 19295
rect 14231 19292 14243 19295
rect 14458 19292 14464 19304
rect 14231 19264 14464 19292
rect 14231 19261 14243 19264
rect 14185 19255 14243 19261
rect 14458 19252 14464 19264
rect 14516 19252 14522 19304
rect 16574 19252 16580 19304
rect 16632 19292 16638 19304
rect 17770 19292 17776 19304
rect 16632 19264 17776 19292
rect 16632 19252 16638 19264
rect 17770 19252 17776 19264
rect 17828 19292 17834 19304
rect 17957 19295 18015 19301
rect 17957 19292 17969 19295
rect 17828 19264 17969 19292
rect 17828 19252 17834 19264
rect 17957 19261 17969 19264
rect 18003 19261 18015 19295
rect 17957 19255 18015 19261
rect 18141 19295 18199 19301
rect 18141 19261 18153 19295
rect 18187 19292 18199 19295
rect 19150 19292 19156 19304
rect 18187 19264 19156 19292
rect 18187 19261 18199 19264
rect 18141 19255 18199 19261
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 10318 19184 10324 19236
rect 10376 19224 10382 19236
rect 10962 19224 10968 19236
rect 10376 19196 10968 19224
rect 10376 19184 10382 19196
rect 10962 19184 10968 19196
rect 11020 19184 11026 19236
rect 12406 19224 12434 19252
rect 18969 19227 19027 19233
rect 12406 19196 14872 19224
rect 14844 19168 14872 19196
rect 18969 19193 18981 19227
rect 19015 19224 19027 19227
rect 19242 19224 19248 19236
rect 19015 19196 19248 19224
rect 19015 19193 19027 19196
rect 18969 19187 19027 19193
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 19720 19224 19748 19332
rect 20806 19320 20812 19332
rect 20864 19320 20870 19372
rect 21082 19320 21088 19372
rect 21140 19320 21146 19372
rect 20073 19295 20131 19301
rect 20073 19261 20085 19295
rect 20119 19292 20131 19295
rect 20622 19292 20628 19304
rect 20119 19264 20628 19292
rect 20119 19261 20131 19264
rect 20073 19255 20131 19261
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 21361 19295 21419 19301
rect 21361 19261 21373 19295
rect 21407 19292 21419 19295
rect 21910 19292 21916 19304
rect 21407 19264 21916 19292
rect 21407 19261 21419 19264
rect 21361 19255 21419 19261
rect 21910 19252 21916 19264
rect 21968 19252 21974 19304
rect 22002 19252 22008 19304
rect 22060 19252 22066 19304
rect 22278 19252 22284 19304
rect 22336 19252 22342 19304
rect 22830 19252 22836 19304
rect 22888 19292 22894 19304
rect 23400 19292 23428 19346
rect 22888 19264 24072 19292
rect 22888 19252 22894 19264
rect 20990 19224 20996 19236
rect 19720 19196 20996 19224
rect 20990 19184 20996 19196
rect 21048 19184 21054 19236
rect 24044 19168 24072 19264
rect 7834 19116 7840 19168
rect 7892 19156 7898 19168
rect 8297 19159 8355 19165
rect 8297 19156 8309 19159
rect 7892 19128 8309 19156
rect 7892 19116 7898 19128
rect 8297 19125 8309 19128
rect 8343 19125 8355 19159
rect 8297 19119 8355 19125
rect 8754 19116 8760 19168
rect 8812 19116 8818 19168
rect 10778 19116 10784 19168
rect 10836 19156 10842 19168
rect 10873 19159 10931 19165
rect 10873 19156 10885 19159
rect 10836 19128 10885 19156
rect 10836 19116 10842 19128
rect 10873 19125 10885 19128
rect 10919 19125 10931 19159
rect 10873 19119 10931 19125
rect 11146 19116 11152 19168
rect 11204 19156 11210 19168
rect 11241 19159 11299 19165
rect 11241 19156 11253 19159
rect 11204 19128 11253 19156
rect 11204 19116 11210 19128
rect 11241 19125 11253 19128
rect 11287 19125 11299 19159
rect 11241 19119 11299 19125
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 13541 19159 13599 19165
rect 13541 19156 13553 19159
rect 12492 19128 13553 19156
rect 12492 19116 12498 19128
rect 13541 19125 13553 19128
rect 13587 19125 13599 19159
rect 13541 19119 13599 19125
rect 14642 19116 14648 19168
rect 14700 19116 14706 19168
rect 14826 19116 14832 19168
rect 14884 19116 14890 19168
rect 24026 19116 24032 19168
rect 24084 19116 24090 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 8938 18912 8944 18964
rect 8996 18912 9002 18964
rect 10594 18952 10600 18964
rect 9048 18924 10600 18952
rect 3786 18844 3792 18896
rect 3844 18884 3850 18896
rect 9048 18884 9076 18924
rect 10594 18912 10600 18924
rect 10652 18912 10658 18964
rect 10778 18912 10784 18964
rect 10836 18952 10842 18964
rect 12158 18952 12164 18964
rect 10836 18924 12164 18952
rect 10836 18912 10842 18924
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 14182 18912 14188 18964
rect 14240 18952 14246 18964
rect 14277 18955 14335 18961
rect 14277 18952 14289 18955
rect 14240 18924 14289 18952
rect 14240 18912 14246 18924
rect 14277 18921 14289 18924
rect 14323 18921 14335 18955
rect 14277 18915 14335 18921
rect 17957 18955 18015 18961
rect 17957 18921 17969 18955
rect 18003 18952 18015 18955
rect 18322 18952 18328 18964
rect 18003 18924 18328 18952
rect 18003 18921 18015 18924
rect 17957 18915 18015 18921
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 18966 18912 18972 18964
rect 19024 18912 19030 18964
rect 22278 18912 22284 18964
rect 22336 18952 22342 18964
rect 24029 18955 24087 18961
rect 24029 18952 24041 18955
rect 22336 18924 24041 18952
rect 22336 18912 22342 18924
rect 24029 18921 24041 18924
rect 24075 18921 24087 18955
rect 24029 18915 24087 18921
rect 3844 18856 9076 18884
rect 3844 18844 3850 18856
rect 13354 18844 13360 18896
rect 13412 18884 13418 18896
rect 13906 18884 13912 18896
rect 13412 18856 13912 18884
rect 13412 18844 13418 18856
rect 13906 18844 13912 18856
rect 13964 18844 13970 18896
rect 19058 18884 19064 18896
rect 17512 18856 19064 18884
rect 1302 18776 1308 18828
rect 1360 18816 1366 18828
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 1360 18788 2053 18816
rect 1360 18776 1366 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 4890 18776 4896 18828
rect 4948 18816 4954 18828
rect 5077 18819 5135 18825
rect 5077 18816 5089 18819
rect 4948 18788 5089 18816
rect 4948 18776 4954 18788
rect 5077 18785 5089 18788
rect 5123 18816 5135 18819
rect 5902 18816 5908 18828
rect 5123 18788 5908 18816
rect 5123 18785 5135 18788
rect 5077 18779 5135 18785
rect 5902 18776 5908 18788
rect 5960 18776 5966 18828
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 12768 18788 13553 18816
rect 12768 18776 12774 18788
rect 13541 18785 13553 18788
rect 13587 18816 13599 18819
rect 14182 18816 14188 18828
rect 13587 18788 14188 18816
rect 13587 18785 13599 18788
rect 13541 18779 13599 18785
rect 14182 18776 14188 18788
rect 14240 18776 14246 18828
rect 14826 18776 14832 18828
rect 14884 18776 14890 18828
rect 17512 18816 17540 18856
rect 19058 18844 19064 18856
rect 19116 18844 19122 18896
rect 16132 18788 17540 18816
rect 1762 18708 1768 18760
rect 1820 18708 1826 18760
rect 4065 18751 4123 18757
rect 4065 18717 4077 18751
rect 4111 18748 4123 18751
rect 5166 18748 5172 18760
rect 4111 18720 5172 18748
rect 4111 18717 4123 18720
rect 4065 18711 4123 18717
rect 5166 18708 5172 18720
rect 5224 18708 5230 18760
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 9232 18720 9781 18748
rect 9232 18689 9260 18720
rect 9769 18717 9781 18720
rect 9815 18717 9827 18751
rect 9769 18711 9827 18717
rect 11146 18708 11152 18760
rect 11204 18748 11210 18760
rect 11885 18751 11943 18757
rect 11885 18748 11897 18751
rect 11204 18720 11897 18748
rect 11204 18708 11210 18720
rect 11885 18717 11897 18720
rect 11931 18748 11943 18751
rect 12802 18748 12808 18760
rect 11931 18720 12808 18748
rect 11931 18717 11943 18720
rect 11885 18711 11943 18717
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 13449 18751 13507 18757
rect 13449 18717 13461 18751
rect 13495 18748 13507 18751
rect 13814 18748 13820 18760
rect 13495 18720 13820 18748
rect 13495 18717 13507 18720
rect 13449 18711 13507 18717
rect 13814 18708 13820 18720
rect 13872 18708 13878 18760
rect 14645 18751 14703 18757
rect 14645 18717 14657 18751
rect 14691 18748 14703 18751
rect 16132 18748 16160 18788
rect 17770 18776 17776 18828
rect 17828 18816 17834 18828
rect 18325 18819 18383 18825
rect 18325 18816 18337 18819
rect 17828 18788 18337 18816
rect 17828 18776 17834 18788
rect 18325 18785 18337 18788
rect 18371 18785 18383 18819
rect 18325 18779 18383 18785
rect 14691 18720 16160 18748
rect 14691 18717 14703 18720
rect 14645 18711 14703 18717
rect 16206 18708 16212 18760
rect 16264 18708 16270 18760
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19024 18720 19625 18748
rect 19024 18708 19030 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18748 20407 18751
rect 20438 18748 20444 18760
rect 20395 18720 20444 18748
rect 20395 18717 20407 18720
rect 20349 18711 20407 18717
rect 20438 18708 20444 18720
rect 20496 18748 20502 18760
rect 21545 18751 21603 18757
rect 21545 18748 21557 18751
rect 20496 18720 21557 18748
rect 20496 18708 20502 18720
rect 21545 18717 21557 18720
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 22002 18708 22008 18760
rect 22060 18748 22066 18760
rect 22281 18751 22339 18757
rect 22281 18748 22293 18751
rect 22060 18720 22293 18748
rect 22060 18708 22094 18720
rect 22281 18717 22293 18720
rect 22327 18717 22339 18751
rect 22281 18711 22339 18717
rect 9217 18683 9275 18689
rect 9217 18680 9229 18683
rect 8496 18652 9229 18680
rect 8496 18624 8524 18652
rect 9217 18649 9229 18652
rect 9263 18649 9275 18683
rect 9217 18643 9275 18649
rect 10045 18683 10103 18689
rect 10045 18649 10057 18683
rect 10091 18649 10103 18683
rect 10045 18643 10103 18649
rect 11348 18652 13032 18680
rect 8478 18572 8484 18624
rect 8536 18572 8542 18624
rect 8662 18572 8668 18624
rect 8720 18572 8726 18624
rect 9306 18572 9312 18624
rect 9364 18612 9370 18624
rect 9401 18615 9459 18621
rect 9401 18612 9413 18615
rect 9364 18584 9413 18612
rect 9364 18572 9370 18584
rect 9401 18581 9413 18584
rect 9447 18612 9459 18615
rect 9582 18612 9588 18624
rect 9447 18584 9588 18612
rect 9447 18581 9459 18584
rect 9401 18575 9459 18581
rect 9582 18572 9588 18584
rect 9640 18612 9646 18624
rect 10060 18612 10088 18643
rect 9640 18584 10088 18612
rect 9640 18572 9646 18584
rect 10870 18572 10876 18624
rect 10928 18612 10934 18624
rect 11348 18612 11376 18652
rect 10928 18584 11376 18612
rect 11517 18615 11575 18621
rect 10928 18572 10934 18584
rect 11517 18581 11529 18615
rect 11563 18612 11575 18615
rect 11606 18612 11612 18624
rect 11563 18584 11612 18612
rect 11563 18581 11575 18584
rect 11517 18575 11575 18581
rect 11606 18572 11612 18584
rect 11664 18572 11670 18624
rect 11974 18572 11980 18624
rect 12032 18612 12038 18624
rect 13004 18621 13032 18652
rect 13630 18640 13636 18692
rect 13688 18680 13694 18692
rect 14737 18683 14795 18689
rect 14737 18680 14749 18683
rect 13688 18652 14749 18680
rect 13688 18640 13694 18652
rect 14737 18649 14749 18652
rect 14783 18649 14795 18683
rect 14737 18643 14795 18649
rect 16485 18683 16543 18689
rect 16485 18649 16497 18683
rect 16531 18649 16543 18683
rect 18509 18683 18567 18689
rect 18509 18680 18521 18683
rect 17710 18652 18521 18680
rect 16485 18643 16543 18649
rect 18509 18649 18521 18652
rect 18555 18680 18567 18683
rect 19426 18680 19432 18692
rect 18555 18652 19432 18680
rect 18555 18649 18567 18652
rect 18509 18643 18567 18649
rect 12069 18615 12127 18621
rect 12069 18612 12081 18615
rect 12032 18584 12081 18612
rect 12032 18572 12038 18584
rect 12069 18581 12081 18584
rect 12115 18581 12127 18615
rect 12069 18575 12127 18581
rect 12989 18615 13047 18621
rect 12989 18581 13001 18615
rect 13035 18581 13047 18615
rect 12989 18575 13047 18581
rect 13354 18572 13360 18624
rect 13412 18572 13418 18624
rect 16500 18612 16528 18643
rect 19426 18640 19432 18652
rect 19484 18640 19490 18692
rect 20898 18640 20904 18692
rect 20956 18680 20962 18692
rect 21085 18683 21143 18689
rect 21085 18680 21097 18683
rect 20956 18652 21097 18680
rect 20956 18640 20962 18652
rect 21085 18649 21097 18652
rect 21131 18680 21143 18683
rect 22066 18680 22094 18708
rect 21131 18652 22094 18680
rect 21131 18649 21143 18652
rect 21085 18643 21143 18649
rect 22554 18640 22560 18692
rect 22612 18640 22618 18692
rect 22940 18652 23046 18680
rect 22940 18624 22968 18652
rect 18414 18612 18420 18624
rect 16500 18584 18420 18612
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 19518 18572 19524 18624
rect 19576 18612 19582 18624
rect 19705 18615 19763 18621
rect 19705 18612 19717 18615
rect 19576 18584 19717 18612
rect 19576 18572 19582 18584
rect 19705 18581 19717 18584
rect 19751 18581 19763 18615
rect 19705 18575 19763 18581
rect 20714 18572 20720 18624
rect 20772 18612 20778 18624
rect 21729 18615 21787 18621
rect 21729 18612 21741 18615
rect 20772 18584 21741 18612
rect 20772 18572 20778 18584
rect 21729 18581 21741 18584
rect 21775 18612 21787 18615
rect 22370 18612 22376 18624
rect 21775 18584 22376 18612
rect 21775 18581 21787 18584
rect 21729 18575 21787 18581
rect 22370 18572 22376 18584
rect 22428 18612 22434 18624
rect 22922 18612 22928 18624
rect 22428 18584 22928 18612
rect 22428 18572 22434 18584
rect 22922 18572 22928 18584
rect 22980 18612 22986 18624
rect 24397 18615 24455 18621
rect 24397 18612 24409 18615
rect 22980 18584 24409 18612
rect 22980 18572 22986 18584
rect 24397 18581 24409 18584
rect 24443 18581 24455 18615
rect 24397 18575 24455 18581
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 7745 18411 7803 18417
rect 7745 18408 7757 18411
rect 7616 18380 7757 18408
rect 7616 18368 7622 18380
rect 7745 18377 7757 18380
rect 7791 18377 7803 18411
rect 9674 18408 9680 18420
rect 7745 18371 7803 18377
rect 8496 18380 9680 18408
rect 8496 18349 8524 18380
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 11054 18368 11060 18420
rect 11112 18408 11118 18420
rect 11701 18411 11759 18417
rect 11701 18408 11713 18411
rect 11112 18380 11713 18408
rect 11112 18368 11118 18380
rect 11701 18377 11713 18380
rect 11747 18377 11759 18411
rect 12894 18408 12900 18420
rect 11701 18371 11759 18377
rect 12636 18380 12900 18408
rect 8481 18343 8539 18349
rect 8481 18309 8493 18343
rect 8527 18309 8539 18343
rect 8481 18303 8539 18309
rect 12069 18343 12127 18349
rect 12069 18309 12081 18343
rect 12115 18340 12127 18343
rect 12434 18340 12440 18352
rect 12115 18312 12440 18340
rect 12115 18309 12127 18312
rect 12069 18303 12127 18309
rect 12434 18300 12440 18312
rect 12492 18300 12498 18352
rect 3329 18275 3387 18281
rect 3329 18241 3341 18275
rect 3375 18272 3387 18275
rect 5258 18272 5264 18284
rect 3375 18244 5264 18272
rect 3375 18241 3387 18244
rect 3329 18235 3387 18241
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 7653 18275 7711 18281
rect 7653 18272 7665 18275
rect 6932 18244 7665 18272
rect 3786 18164 3792 18216
rect 3844 18164 3850 18216
rect 4982 18028 4988 18080
rect 5040 18068 5046 18080
rect 6932 18077 6960 18244
rect 7653 18241 7665 18244
rect 7699 18241 7711 18275
rect 7653 18235 7711 18241
rect 7742 18232 7748 18284
rect 7800 18272 7806 18284
rect 10781 18275 10839 18281
rect 7800 18244 10456 18272
rect 7800 18232 7806 18244
rect 7098 18164 7104 18216
rect 7156 18204 7162 18216
rect 7834 18204 7840 18216
rect 7156 18176 7840 18204
rect 7156 18164 7162 18176
rect 7834 18164 7840 18176
rect 7892 18164 7898 18216
rect 9217 18207 9275 18213
rect 9217 18173 9229 18207
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 8478 18096 8484 18148
rect 8536 18136 8542 18148
rect 9232 18136 9260 18167
rect 10428 18145 10456 18244
rect 10781 18241 10793 18275
rect 10827 18272 10839 18275
rect 11974 18272 11980 18284
rect 10827 18244 11980 18272
rect 10827 18241 10839 18244
rect 10781 18235 10839 18241
rect 11974 18232 11980 18244
rect 12032 18272 12038 18284
rect 12636 18272 12664 18380
rect 12894 18368 12900 18380
rect 12952 18368 12958 18420
rect 13354 18368 13360 18420
rect 13412 18408 13418 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 13412 18380 14289 18408
rect 13412 18368 13418 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 14645 18411 14703 18417
rect 14645 18377 14657 18411
rect 14691 18408 14703 18411
rect 15381 18411 15439 18417
rect 15381 18408 15393 18411
rect 14691 18380 15393 18408
rect 14691 18377 14703 18380
rect 14645 18371 14703 18377
rect 15381 18377 15393 18380
rect 15427 18408 15439 18411
rect 18322 18408 18328 18420
rect 15427 18380 18328 18408
rect 15427 18377 15439 18380
rect 15381 18371 15439 18377
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 21821 18411 21879 18417
rect 21821 18408 21833 18411
rect 19536 18380 21833 18408
rect 13817 18343 13875 18349
rect 13817 18309 13829 18343
rect 13863 18340 13875 18343
rect 13863 18312 14780 18340
rect 13863 18309 13875 18312
rect 13817 18303 13875 18309
rect 12032 18244 12664 18272
rect 12032 18232 12038 18244
rect 12710 18232 12716 18284
rect 12768 18272 12774 18284
rect 14752 18281 14780 18312
rect 19150 18300 19156 18352
rect 19208 18300 19214 18352
rect 19426 18300 19432 18352
rect 19484 18340 19490 18352
rect 19536 18340 19564 18380
rect 21821 18377 21833 18380
rect 21867 18408 21879 18411
rect 21867 18380 22094 18408
rect 21867 18377 21879 18380
rect 21821 18371 21879 18377
rect 19484 18312 19642 18340
rect 19484 18300 19490 18312
rect 14737 18275 14795 18281
rect 12768 18244 14596 18272
rect 12768 18232 12774 18244
rect 10686 18164 10692 18216
rect 10744 18204 10750 18216
rect 10873 18207 10931 18213
rect 10873 18204 10885 18207
rect 10744 18176 10885 18204
rect 10744 18164 10750 18176
rect 10873 18173 10885 18176
rect 10919 18173 10931 18207
rect 10873 18167 10931 18173
rect 10962 18164 10968 18216
rect 11020 18164 11026 18216
rect 12158 18164 12164 18216
rect 12216 18164 12222 18216
rect 12250 18164 12256 18216
rect 12308 18164 12314 18216
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 14458 18204 14464 18216
rect 12492 18176 14464 18204
rect 12492 18164 12498 18176
rect 14458 18164 14464 18176
rect 14516 18164 14522 18216
rect 14568 18204 14596 18244
rect 14737 18241 14749 18275
rect 14783 18272 14795 18275
rect 15010 18272 15016 18284
rect 14783 18244 15016 18272
rect 14783 18241 14795 18244
rect 14737 18235 14795 18241
rect 15010 18232 15016 18244
rect 15068 18232 15074 18284
rect 17494 18232 17500 18284
rect 17552 18232 17558 18284
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 22066 18272 22094 18380
rect 22373 18275 22431 18281
rect 22373 18272 22385 18275
rect 22066 18244 22385 18272
rect 21269 18235 21327 18241
rect 22373 18241 22385 18244
rect 22419 18272 22431 18275
rect 24026 18272 24032 18284
rect 22419 18244 24032 18272
rect 22419 18241 22431 18244
rect 22373 18235 22431 18241
rect 14921 18207 14979 18213
rect 14921 18204 14933 18207
rect 14568 18176 14933 18204
rect 14921 18173 14933 18176
rect 14967 18204 14979 18207
rect 15378 18204 15384 18216
rect 14967 18176 15384 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 15378 18164 15384 18176
rect 15436 18204 15442 18216
rect 16022 18204 16028 18216
rect 15436 18176 16028 18204
rect 15436 18164 15442 18176
rect 16022 18164 16028 18176
rect 16080 18164 16086 18216
rect 16206 18164 16212 18216
rect 16264 18204 16270 18216
rect 16482 18204 16488 18216
rect 16264 18176 16488 18204
rect 16264 18164 16270 18176
rect 16482 18164 16488 18176
rect 16540 18204 16546 18216
rect 18325 18207 18383 18213
rect 18325 18204 18337 18207
rect 16540 18176 18337 18204
rect 16540 18164 16546 18176
rect 18325 18173 18337 18176
rect 18371 18204 18383 18207
rect 18877 18207 18935 18213
rect 18877 18204 18889 18207
rect 18371 18176 18889 18204
rect 18371 18173 18383 18176
rect 18325 18167 18383 18173
rect 18877 18173 18889 18176
rect 18923 18173 18935 18207
rect 21284 18204 21312 18235
rect 24026 18232 24032 18244
rect 24084 18232 24090 18284
rect 18877 18167 18935 18173
rect 18984 18176 21312 18204
rect 8536 18108 9260 18136
rect 10413 18139 10471 18145
rect 8536 18096 8542 18108
rect 10413 18105 10425 18139
rect 10459 18105 10471 18139
rect 10413 18099 10471 18105
rect 12342 18096 12348 18148
rect 12400 18136 12406 18148
rect 12526 18136 12532 18148
rect 12400 18108 12532 18136
rect 12400 18096 12406 18108
rect 12526 18096 12532 18108
rect 12584 18136 12590 18148
rect 13630 18136 13636 18148
rect 12584 18108 13636 18136
rect 12584 18096 12590 18108
rect 13630 18096 13636 18108
rect 13688 18136 13694 18148
rect 13909 18139 13967 18145
rect 13909 18136 13921 18139
rect 13688 18108 13921 18136
rect 13688 18096 13694 18108
rect 13909 18105 13921 18108
rect 13955 18105 13967 18139
rect 13909 18099 13967 18105
rect 18506 18096 18512 18148
rect 18564 18136 18570 18148
rect 18984 18136 19012 18176
rect 22922 18164 22928 18216
rect 22980 18204 22986 18216
rect 23385 18207 23443 18213
rect 23385 18204 23397 18207
rect 22980 18176 23397 18204
rect 22980 18164 22986 18176
rect 23385 18173 23397 18176
rect 23431 18204 23443 18207
rect 23658 18204 23664 18216
rect 23431 18176 23664 18204
rect 23431 18173 23443 18176
rect 23385 18167 23443 18173
rect 23658 18164 23664 18176
rect 23716 18164 23722 18216
rect 18564 18108 19012 18136
rect 18564 18096 18570 18108
rect 21450 18096 21456 18148
rect 21508 18096 21514 18148
rect 6917 18071 6975 18077
rect 6917 18068 6929 18071
rect 5040 18040 6929 18068
rect 5040 18028 5046 18040
rect 6917 18037 6929 18040
rect 6963 18037 6975 18071
rect 6917 18031 6975 18037
rect 7285 18071 7343 18077
rect 7285 18037 7297 18071
rect 7331 18068 7343 18071
rect 7742 18068 7748 18080
rect 7331 18040 7748 18068
rect 7331 18037 7343 18040
rect 7285 18031 7343 18037
rect 7742 18028 7748 18040
rect 7800 18028 7806 18080
rect 10137 18071 10195 18077
rect 10137 18037 10149 18071
rect 10183 18068 10195 18071
rect 10686 18068 10692 18080
rect 10183 18040 10692 18068
rect 10183 18037 10195 18040
rect 10137 18031 10195 18037
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 11606 18028 11612 18080
rect 11664 18068 11670 18080
rect 12250 18068 12256 18080
rect 11664 18040 12256 18068
rect 11664 18028 11670 18040
rect 12250 18028 12256 18040
rect 12308 18028 12314 18080
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 13998 18068 14004 18080
rect 13596 18040 14004 18068
rect 13596 18028 13602 18040
rect 13998 18028 14004 18040
rect 14056 18068 14062 18080
rect 14734 18068 14740 18080
rect 14056 18040 14740 18068
rect 14056 18028 14062 18040
rect 14734 18028 14740 18040
rect 14792 18028 14798 18080
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 17129 18071 17187 18077
rect 17129 18068 17141 18071
rect 16632 18040 17141 18068
rect 16632 18028 16638 18040
rect 17129 18037 17141 18040
rect 17175 18068 17187 18071
rect 17494 18068 17500 18080
rect 17175 18040 17500 18068
rect 17175 18037 17187 18040
rect 17129 18031 17187 18037
rect 17494 18028 17500 18040
rect 17552 18028 17558 18080
rect 20162 18028 20168 18080
rect 20220 18068 20226 18080
rect 20625 18071 20683 18077
rect 20625 18068 20637 18071
rect 20220 18040 20637 18068
rect 20220 18028 20226 18040
rect 20625 18037 20637 18040
rect 20671 18037 20683 18071
rect 20625 18031 20683 18037
rect 23937 18071 23995 18077
rect 23937 18037 23949 18071
rect 23983 18068 23995 18071
rect 24026 18068 24032 18080
rect 23983 18040 24032 18068
rect 23983 18037 23995 18040
rect 23937 18031 23995 18037
rect 24026 18028 24032 18040
rect 24084 18028 24090 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 6270 17824 6276 17876
rect 6328 17824 6334 17876
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 9125 17867 9183 17873
rect 9125 17864 9137 17867
rect 7432 17836 9137 17864
rect 7432 17824 7438 17836
rect 9125 17833 9137 17836
rect 9171 17833 9183 17867
rect 9125 17827 9183 17833
rect 11882 17824 11888 17876
rect 11940 17864 11946 17876
rect 12526 17864 12532 17876
rect 11940 17836 12532 17864
rect 11940 17824 11946 17836
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 12710 17824 12716 17876
rect 12768 17864 12774 17876
rect 12894 17864 12900 17876
rect 12768 17836 12900 17864
rect 12768 17824 12774 17836
rect 12894 17824 12900 17836
rect 12952 17824 12958 17876
rect 15102 17824 15108 17876
rect 15160 17864 15166 17876
rect 19242 17864 19248 17876
rect 15160 17836 19248 17864
rect 15160 17824 15166 17836
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 20622 17824 20628 17876
rect 20680 17864 20686 17876
rect 21637 17867 21695 17873
rect 21637 17864 21649 17867
rect 20680 17836 21649 17864
rect 20680 17824 20686 17836
rect 21637 17833 21649 17836
rect 21683 17864 21695 17867
rect 21683 17836 22232 17864
rect 21683 17833 21695 17836
rect 21637 17827 21695 17833
rect 17221 17799 17279 17805
rect 17221 17796 17233 17799
rect 16684 17768 17233 17796
rect 6825 17731 6883 17737
rect 6825 17697 6837 17731
rect 6871 17728 6883 17731
rect 6914 17728 6920 17740
rect 6871 17700 6920 17728
rect 6871 17697 6883 17700
rect 6825 17691 6883 17697
rect 6914 17688 6920 17700
rect 6972 17688 6978 17740
rect 8113 17731 8171 17737
rect 8113 17697 8125 17731
rect 8159 17728 8171 17731
rect 8386 17728 8392 17740
rect 8159 17700 8392 17728
rect 8159 17697 8171 17700
rect 8113 17691 8171 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9456 17700 9689 17728
rect 9456 17688 9462 17700
rect 9677 17697 9689 17700
rect 9723 17697 9735 17731
rect 9677 17691 9735 17697
rect 11974 17688 11980 17740
rect 12032 17728 12038 17740
rect 12713 17731 12771 17737
rect 12713 17728 12725 17731
rect 12032 17700 12725 17728
rect 12032 17688 12038 17700
rect 12713 17697 12725 17700
rect 12759 17728 12771 17731
rect 13541 17731 13599 17737
rect 13541 17728 13553 17731
rect 12759 17700 13553 17728
rect 12759 17697 12771 17700
rect 12713 17691 12771 17697
rect 13541 17697 13553 17700
rect 13587 17697 13599 17731
rect 13541 17691 13599 17697
rect 14458 17688 14464 17740
rect 14516 17728 14522 17740
rect 14826 17728 14832 17740
rect 14516 17700 14832 17728
rect 14516 17688 14522 17700
rect 14826 17688 14832 17700
rect 14884 17688 14890 17740
rect 16390 17688 16396 17740
rect 16448 17728 16454 17740
rect 16684 17737 16712 17768
rect 17221 17765 17233 17768
rect 17267 17765 17279 17799
rect 17221 17759 17279 17765
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 16448 17700 16681 17728
rect 16448 17688 16454 17700
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 16853 17731 16911 17737
rect 16853 17697 16865 17731
rect 16899 17728 16911 17731
rect 17034 17728 17040 17740
rect 16899 17700 17040 17728
rect 16899 17697 16911 17700
rect 16853 17691 16911 17697
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 19889 17731 19947 17737
rect 19889 17697 19901 17731
rect 19935 17728 19947 17731
rect 20898 17728 20904 17740
rect 19935 17700 20904 17728
rect 19935 17697 19947 17700
rect 19889 17691 19947 17697
rect 20898 17688 20904 17700
rect 20956 17728 20962 17740
rect 22097 17731 22155 17737
rect 22097 17728 22109 17731
rect 20956 17700 22109 17728
rect 20956 17688 20962 17700
rect 22097 17697 22109 17700
rect 22143 17697 22155 17731
rect 22204 17728 22232 17836
rect 22554 17824 22560 17876
rect 22612 17864 22618 17876
rect 23845 17867 23903 17873
rect 23845 17864 23857 17867
rect 22612 17836 23857 17864
rect 22612 17824 22618 17836
rect 23845 17833 23857 17836
rect 23891 17833 23903 17867
rect 23845 17827 23903 17833
rect 22373 17731 22431 17737
rect 22373 17728 22385 17731
rect 22204 17700 22385 17728
rect 22097 17691 22155 17697
rect 22373 17697 22385 17700
rect 22419 17697 22431 17731
rect 22373 17691 22431 17697
rect 4706 17620 4712 17672
rect 4764 17660 4770 17672
rect 7929 17663 7987 17669
rect 4764 17632 7604 17660
rect 4764 17620 4770 17632
rect 6641 17595 6699 17601
rect 6641 17561 6653 17595
rect 6687 17592 6699 17595
rect 7576 17592 7604 17632
rect 7929 17629 7941 17663
rect 7975 17660 7987 17663
rect 8754 17660 8760 17672
rect 7975 17632 8760 17660
rect 7975 17629 7987 17632
rect 7929 17623 7987 17629
rect 8754 17620 8760 17632
rect 8812 17620 8818 17672
rect 9582 17620 9588 17672
rect 9640 17660 9646 17672
rect 11885 17663 11943 17669
rect 11885 17660 11897 17663
rect 9640 17632 11897 17660
rect 9640 17620 9646 17632
rect 11885 17629 11897 17632
rect 11931 17629 11943 17663
rect 11885 17623 11943 17629
rect 12526 17620 12532 17672
rect 12584 17660 12590 17672
rect 13449 17663 13507 17669
rect 13449 17660 13461 17663
rect 12584 17632 13461 17660
rect 12584 17620 12590 17632
rect 13449 17629 13461 17632
rect 13495 17629 13507 17663
rect 13449 17623 13507 17629
rect 14642 17620 14648 17672
rect 14700 17660 14706 17672
rect 15102 17660 15108 17672
rect 14700 17632 15108 17660
rect 14700 17620 14706 17632
rect 15102 17620 15108 17632
rect 15160 17620 15166 17672
rect 15562 17620 15568 17672
rect 15620 17620 15626 17672
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 16206 17660 16212 17672
rect 15712 17632 16212 17660
rect 15712 17620 15718 17632
rect 16206 17620 16212 17632
rect 16264 17620 16270 17672
rect 24857 17663 24915 17669
rect 24857 17629 24869 17663
rect 24903 17660 24915 17663
rect 25038 17660 25044 17672
rect 24903 17632 25044 17660
rect 24903 17629 24915 17632
rect 24857 17623 24915 17629
rect 25038 17620 25044 17632
rect 25096 17620 25102 17672
rect 6687 17564 7512 17592
rect 7576 17564 8800 17592
rect 6687 17561 6699 17564
rect 6641 17555 6699 17561
rect 6733 17527 6791 17533
rect 6733 17493 6745 17527
rect 6779 17524 6791 17527
rect 7282 17524 7288 17536
rect 6779 17496 7288 17524
rect 6779 17493 6791 17496
rect 6733 17487 6791 17493
rect 7282 17484 7288 17496
rect 7340 17484 7346 17536
rect 7484 17533 7512 17564
rect 8772 17536 8800 17564
rect 9674 17552 9680 17604
rect 9732 17592 9738 17604
rect 10502 17592 10508 17604
rect 9732 17564 10508 17592
rect 9732 17552 9738 17564
rect 10502 17552 10508 17564
rect 10560 17552 10566 17604
rect 11330 17552 11336 17604
rect 11388 17552 11394 17604
rect 13357 17595 13415 17601
rect 13357 17561 13369 17595
rect 13403 17592 13415 17595
rect 15672 17592 15700 17620
rect 18874 17592 18880 17604
rect 13403 17564 15700 17592
rect 16224 17564 18880 17592
rect 13403 17561 13415 17564
rect 13357 17555 13415 17561
rect 7469 17527 7527 17533
rect 7469 17493 7481 17527
rect 7515 17493 7527 17527
rect 7469 17487 7527 17493
rect 7837 17527 7895 17533
rect 7837 17493 7849 17527
rect 7883 17524 7895 17527
rect 8570 17524 8576 17536
rect 7883 17496 8576 17524
rect 7883 17493 7895 17496
rect 7837 17487 7895 17493
rect 8570 17484 8576 17496
rect 8628 17484 8634 17536
rect 8754 17484 8760 17536
rect 8812 17484 8818 17536
rect 9490 17484 9496 17536
rect 9548 17484 9554 17536
rect 9585 17527 9643 17533
rect 9585 17493 9597 17527
rect 9631 17524 9643 17527
rect 10134 17524 10140 17536
rect 9631 17496 10140 17524
rect 9631 17493 9643 17496
rect 9585 17487 9643 17493
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 12989 17527 13047 17533
rect 12989 17524 13001 17527
rect 12768 17496 13001 17524
rect 12768 17484 12774 17496
rect 12989 17493 13001 17496
rect 13035 17493 13047 17527
rect 12989 17487 13047 17493
rect 13538 17484 13544 17536
rect 13596 17524 13602 17536
rect 14277 17527 14335 17533
rect 14277 17524 14289 17527
rect 13596 17496 14289 17524
rect 13596 17484 13602 17496
rect 14277 17493 14289 17496
rect 14323 17493 14335 17527
rect 14277 17487 14335 17493
rect 14734 17484 14740 17536
rect 14792 17484 14798 17536
rect 15378 17484 15384 17536
rect 15436 17524 15442 17536
rect 16224 17533 16252 17564
rect 18874 17552 18880 17564
rect 18932 17552 18938 17604
rect 20162 17552 20168 17604
rect 20220 17552 20226 17604
rect 20714 17552 20720 17604
rect 20772 17552 20778 17604
rect 23658 17592 23664 17604
rect 23598 17564 23664 17592
rect 23658 17552 23664 17564
rect 23716 17592 23722 17604
rect 24121 17595 24179 17601
rect 24121 17592 24133 17595
rect 23716 17564 24133 17592
rect 23716 17552 23722 17564
rect 24121 17561 24133 17564
rect 24167 17561 24179 17595
rect 24121 17555 24179 17561
rect 15657 17527 15715 17533
rect 15657 17524 15669 17527
rect 15436 17496 15669 17524
rect 15436 17484 15442 17496
rect 15657 17493 15669 17496
rect 15703 17493 15715 17527
rect 15657 17487 15715 17493
rect 16209 17527 16267 17533
rect 16209 17493 16221 17527
rect 16255 17493 16267 17527
rect 16209 17487 16267 17493
rect 16390 17484 16396 17536
rect 16448 17524 16454 17536
rect 16577 17527 16635 17533
rect 16577 17524 16589 17527
rect 16448 17496 16589 17524
rect 16448 17484 16454 17496
rect 16577 17493 16589 17496
rect 16623 17493 16635 17527
rect 16577 17487 16635 17493
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 24673 17527 24731 17533
rect 24673 17524 24685 17527
rect 24268 17496 24685 17524
rect 24268 17484 24274 17496
rect 24673 17493 24685 17496
rect 24719 17493 24731 17527
rect 24673 17487 24731 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 8846 17280 8852 17332
rect 8904 17320 8910 17332
rect 8904 17292 9444 17320
rect 8904 17280 8910 17292
rect 3694 17212 3700 17264
rect 3752 17252 3758 17264
rect 3970 17252 3976 17264
rect 3752 17224 3976 17252
rect 3752 17212 3758 17224
rect 3970 17212 3976 17224
rect 4028 17212 4034 17264
rect 8110 17252 8116 17264
rect 8050 17224 8116 17252
rect 8110 17212 8116 17224
rect 8168 17252 8174 17264
rect 8938 17252 8944 17264
rect 8168 17224 8944 17252
rect 8168 17212 8174 17224
rect 8938 17212 8944 17224
rect 8996 17212 9002 17264
rect 9416 17252 9444 17292
rect 9490 17280 9496 17332
rect 9548 17320 9554 17332
rect 10045 17323 10103 17329
rect 10045 17320 10057 17323
rect 9548 17292 10057 17320
rect 9548 17280 9554 17292
rect 10045 17289 10057 17292
rect 10091 17289 10103 17323
rect 10045 17283 10103 17289
rect 10502 17280 10508 17332
rect 10560 17320 10566 17332
rect 11517 17323 11575 17329
rect 11517 17320 11529 17323
rect 10560 17292 11529 17320
rect 10560 17280 10566 17292
rect 11517 17289 11529 17292
rect 11563 17320 11575 17323
rect 16574 17320 16580 17332
rect 11563 17292 16580 17320
rect 11563 17289 11575 17292
rect 11517 17283 11575 17289
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 20898 17320 20904 17332
rect 17696 17292 20904 17320
rect 10413 17255 10471 17261
rect 9416 17224 9674 17252
rect 3145 17187 3203 17193
rect 3145 17153 3157 17187
rect 3191 17184 3203 17187
rect 4614 17184 4620 17196
rect 3191 17156 4620 17184
rect 3191 17153 3203 17156
rect 3145 17147 3203 17153
rect 4614 17144 4620 17156
rect 4672 17144 4678 17196
rect 8754 17144 8760 17196
rect 8812 17184 8818 17196
rect 9033 17187 9091 17193
rect 9033 17184 9045 17187
rect 8812 17156 9045 17184
rect 8812 17144 8818 17156
rect 9033 17153 9045 17156
rect 9079 17153 9091 17187
rect 9033 17147 9091 17153
rect 6546 17076 6552 17128
rect 6604 17076 6610 17128
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 6914 17116 6920 17128
rect 6871 17088 6920 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 6914 17076 6920 17088
rect 6972 17076 6978 17128
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 8846 17116 8852 17128
rect 8619 17088 8852 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 8846 17076 8852 17088
rect 8904 17076 8910 17128
rect 9646 17116 9674 17224
rect 10413 17221 10425 17255
rect 10459 17252 10471 17255
rect 12066 17252 12072 17264
rect 10459 17224 12072 17252
rect 10459 17221 10471 17224
rect 10413 17215 10471 17221
rect 12066 17212 12072 17224
rect 12124 17212 12130 17264
rect 12802 17212 12808 17264
rect 12860 17252 12866 17264
rect 13354 17252 13360 17264
rect 12860 17224 13360 17252
rect 12860 17212 12866 17224
rect 13354 17212 13360 17224
rect 13412 17212 13418 17264
rect 15102 17212 15108 17264
rect 15160 17212 15166 17264
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17184 17095 17187
rect 17126 17184 17132 17196
rect 17083 17156 17132 17184
rect 17083 17153 17095 17156
rect 17037 17147 17095 17153
rect 17126 17144 17132 17156
rect 17184 17144 17190 17196
rect 17696 17193 17724 17292
rect 20898 17280 20904 17292
rect 20956 17280 20962 17332
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 19797 17255 19855 17261
rect 18012 17224 18446 17252
rect 18012 17212 18018 17224
rect 19797 17221 19809 17255
rect 19843 17252 19855 17255
rect 20714 17252 20720 17264
rect 19843 17224 20720 17252
rect 19843 17221 19855 17224
rect 19797 17215 19855 17221
rect 20714 17212 20720 17224
rect 20772 17212 20778 17264
rect 23293 17255 23351 17261
rect 23293 17221 23305 17255
rect 23339 17252 23351 17255
rect 24854 17252 24860 17264
rect 23339 17224 24860 17252
rect 23339 17221 23351 17224
rect 23293 17215 23351 17221
rect 24854 17212 24860 17224
rect 24912 17212 24918 17264
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17153 21327 17187
rect 21269 17147 21327 17153
rect 9140 17088 9444 17116
rect 9646 17088 10456 17116
rect 9140 16989 9168 17088
rect 9416 17048 9444 17088
rect 9950 17048 9956 17060
rect 9416 17020 9956 17048
rect 9950 17008 9956 17020
rect 10008 17008 10014 17060
rect 10428 17048 10456 17088
rect 10502 17076 10508 17128
rect 10560 17076 10566 17128
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 10962 17116 10968 17128
rect 10735 17088 10968 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 10962 17076 10968 17088
rect 11020 17076 11026 17128
rect 11330 17076 11336 17128
rect 11388 17116 11394 17128
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 11388 17088 12633 17116
rect 11388 17076 11394 17088
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 12894 17076 12900 17128
rect 12952 17076 12958 17128
rect 13354 17076 13360 17128
rect 13412 17116 13418 17128
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 13412 17088 14933 17116
rect 13412 17076 13418 17088
rect 14921 17085 14933 17088
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 17957 17119 18015 17125
rect 17957 17085 17969 17119
rect 18003 17116 18015 17119
rect 18598 17116 18604 17128
rect 18003 17088 18604 17116
rect 18003 17085 18015 17088
rect 17957 17079 18015 17085
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 19150 17076 19156 17128
rect 19208 17116 19214 17128
rect 19429 17119 19487 17125
rect 19429 17116 19441 17119
rect 19208 17088 19441 17116
rect 19208 17076 19214 17088
rect 19429 17085 19441 17088
rect 19475 17085 19487 17119
rect 19429 17079 19487 17085
rect 20438 17076 20444 17128
rect 20496 17076 20502 17128
rect 11054 17048 11060 17060
rect 10428 17020 11060 17048
rect 11054 17008 11060 17020
rect 11112 17048 11118 17060
rect 12434 17048 12440 17060
rect 11112 17020 12440 17048
rect 11112 17008 11118 17020
rect 12434 17008 12440 17020
rect 12492 17008 12498 17060
rect 14182 17008 14188 17060
rect 14240 17048 14246 17060
rect 14369 17051 14427 17057
rect 14369 17048 14381 17051
rect 14240 17020 14381 17048
rect 14240 17008 14246 17020
rect 14369 17017 14381 17020
rect 14415 17017 14427 17051
rect 14369 17011 14427 17017
rect 15010 17008 15016 17060
rect 15068 17048 15074 17060
rect 16025 17051 16083 17057
rect 16025 17048 16037 17051
rect 15068 17020 16037 17048
rect 15068 17008 15074 17020
rect 16025 17017 16037 17020
rect 16071 17048 16083 17051
rect 16390 17048 16396 17060
rect 16071 17020 16396 17048
rect 16071 17017 16083 17020
rect 16025 17011 16083 17017
rect 16390 17008 16396 17020
rect 16448 17008 16454 17060
rect 9125 16983 9183 16989
rect 9125 16949 9137 16983
rect 9171 16949 9183 16983
rect 9125 16943 9183 16949
rect 9490 16940 9496 16992
rect 9548 16940 9554 16992
rect 9968 16980 9996 17008
rect 11606 16980 11612 16992
rect 9968 16952 11612 16980
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 14458 16940 14464 16992
rect 14516 16980 14522 16992
rect 14737 16983 14795 16989
rect 14737 16980 14749 16983
rect 14516 16952 14749 16980
rect 14516 16940 14522 16952
rect 14737 16949 14749 16952
rect 14783 16949 14795 16983
rect 14737 16943 14795 16949
rect 16850 16940 16856 16992
rect 16908 16940 16914 16992
rect 17218 16940 17224 16992
rect 17276 16980 17282 16992
rect 21284 16980 21312 17147
rect 22094 17144 22100 17196
rect 22152 17144 22158 17196
rect 23934 17144 23940 17196
rect 23992 17144 23998 17196
rect 23290 17076 23296 17128
rect 23348 17116 23354 17128
rect 24397 17119 24455 17125
rect 24397 17116 24409 17119
rect 23348 17088 24409 17116
rect 23348 17076 23354 17088
rect 24397 17085 24409 17088
rect 24443 17085 24455 17119
rect 24397 17079 24455 17085
rect 21453 17051 21511 17057
rect 21453 17017 21465 17051
rect 21499 17048 21511 17051
rect 21726 17048 21732 17060
rect 21499 17020 21732 17048
rect 21499 17017 21511 17020
rect 21453 17011 21511 17017
rect 21726 17008 21732 17020
rect 21784 17008 21790 17060
rect 17276 16952 21312 16980
rect 17276 16940 17282 16952
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 5616 16779 5674 16785
rect 5616 16745 5628 16779
rect 5662 16776 5674 16779
rect 5662 16748 6868 16776
rect 5662 16745 5674 16748
rect 5616 16739 5674 16745
rect 6840 16708 6868 16748
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7101 16779 7159 16785
rect 7101 16776 7113 16779
rect 6972 16748 7113 16776
rect 6972 16736 6978 16748
rect 7101 16745 7113 16748
rect 7147 16745 7159 16779
rect 7101 16739 7159 16745
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 7469 16779 7527 16785
rect 7469 16776 7481 16779
rect 7248 16748 7481 16776
rect 7248 16736 7254 16748
rect 7469 16745 7481 16748
rect 7515 16776 7527 16779
rect 8110 16776 8116 16788
rect 7515 16748 8116 16776
rect 7515 16745 7527 16748
rect 7469 16739 7527 16745
rect 8110 16736 8116 16748
rect 8168 16776 8174 16788
rect 8168 16748 8524 16776
rect 8168 16736 8174 16748
rect 8386 16708 8392 16720
rect 6840 16680 8392 16708
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 8496 16708 8524 16748
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 8628 16748 9137 16776
rect 8628 16736 8634 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9125 16739 9183 16745
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 10505 16779 10563 16785
rect 10505 16776 10517 16779
rect 10192 16748 10517 16776
rect 10192 16736 10198 16748
rect 10505 16745 10517 16748
rect 10551 16745 10563 16779
rect 12802 16776 12808 16788
rect 10505 16739 10563 16745
rect 10612 16748 12808 16776
rect 8665 16711 8723 16717
rect 8665 16708 8677 16711
rect 8496 16680 8677 16708
rect 8665 16677 8677 16680
rect 8711 16708 8723 16711
rect 8754 16708 8760 16720
rect 8711 16680 8760 16708
rect 8711 16677 8723 16680
rect 8665 16671 8723 16677
rect 8754 16668 8760 16680
rect 8812 16668 8818 16720
rect 9950 16668 9956 16720
rect 10008 16708 10014 16720
rect 10229 16711 10287 16717
rect 10229 16708 10241 16711
rect 10008 16680 10241 16708
rect 10008 16668 10014 16680
rect 10229 16677 10241 16680
rect 10275 16677 10287 16711
rect 10229 16671 10287 16677
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16640 5411 16643
rect 6638 16640 6644 16652
rect 5399 16612 6644 16640
rect 5399 16609 5411 16612
rect 5353 16603 5411 16609
rect 6638 16600 6644 16612
rect 6696 16640 6702 16652
rect 7653 16643 7711 16649
rect 7653 16640 7665 16643
rect 6696 16612 7665 16640
rect 6696 16600 6702 16612
rect 7653 16609 7665 16612
rect 7699 16640 7711 16643
rect 8478 16640 8484 16652
rect 7699 16612 8484 16640
rect 7699 16609 7711 16612
rect 7653 16603 7711 16609
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 9416 16612 9689 16640
rect 1486 16532 1492 16584
rect 1544 16572 1550 16584
rect 1581 16575 1639 16581
rect 1581 16572 1593 16575
rect 1544 16544 1593 16572
rect 1544 16532 1550 16544
rect 1581 16541 1593 16544
rect 1627 16541 1639 16575
rect 1581 16535 1639 16541
rect 8294 16532 8300 16584
rect 8352 16572 8358 16584
rect 9030 16572 9036 16584
rect 8352 16544 9036 16572
rect 8352 16532 8358 16544
rect 9030 16532 9036 16544
rect 9088 16572 9094 16584
rect 9416 16572 9444 16612
rect 9677 16609 9689 16612
rect 9723 16640 9735 16643
rect 10612 16640 10640 16748
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 19337 16779 19395 16785
rect 19337 16776 19349 16779
rect 15764 16748 19349 16776
rect 14274 16708 14280 16720
rect 12268 16680 14280 16708
rect 9723 16612 10640 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 10962 16600 10968 16652
rect 11020 16640 11026 16652
rect 12268 16649 12296 16680
rect 14274 16668 14280 16680
rect 14332 16668 14338 16720
rect 11057 16643 11115 16649
rect 11057 16640 11069 16643
rect 11020 16612 11069 16640
rect 11020 16600 11026 16612
rect 11057 16609 11069 16612
rect 11103 16609 11115 16643
rect 11057 16603 11115 16609
rect 12253 16643 12311 16649
rect 12253 16609 12265 16643
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16640 12403 16643
rect 12802 16640 12808 16652
rect 12391 16612 12808 16640
rect 12391 16609 12403 16612
rect 12345 16603 12403 16609
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 14918 16600 14924 16652
rect 14976 16640 14982 16652
rect 15764 16649 15792 16748
rect 19337 16745 19349 16748
rect 19383 16776 19395 16779
rect 19702 16776 19708 16788
rect 19383 16748 19708 16776
rect 19383 16745 19395 16748
rect 19337 16739 19395 16745
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 20162 16736 20168 16788
rect 20220 16776 20226 16788
rect 20220 16748 20668 16776
rect 20220 16736 20226 16748
rect 18690 16668 18696 16720
rect 18748 16708 18754 16720
rect 18748 16680 20576 16708
rect 18748 16668 18754 16680
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 14976 16612 15761 16640
rect 14976 16600 14982 16612
rect 15749 16609 15761 16612
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16022 16640 16028 16652
rect 15979 16612 16028 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16022 16600 16028 16612
rect 16080 16600 16086 16652
rect 9088 16544 9444 16572
rect 9493 16575 9551 16581
rect 9088 16532 9094 16544
rect 9493 16541 9505 16575
rect 9539 16572 9551 16575
rect 9582 16572 9588 16584
rect 9539 16544 9588 16572
rect 9539 16541 9551 16544
rect 9493 16535 9551 16541
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 10318 16572 10324 16584
rect 9876 16544 10324 16572
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 7190 16504 7196 16516
rect 6854 16476 7196 16504
rect 2501 16467 2559 16473
rect 7190 16464 7196 16476
rect 7248 16464 7254 16516
rect 9876 16504 9904 16544
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 10870 16532 10876 16584
rect 10928 16532 10934 16584
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16572 12219 16575
rect 12710 16572 12716 16584
rect 12207 16544 12716 16572
rect 12207 16541 12219 16544
rect 12161 16535 12219 16541
rect 12710 16532 12716 16544
rect 12768 16532 12774 16584
rect 20438 16532 20444 16584
rect 20496 16532 20502 16584
rect 20548 16581 20576 16680
rect 20640 16649 20668 16748
rect 20625 16643 20683 16649
rect 20625 16609 20637 16643
rect 20671 16609 20683 16643
rect 20625 16603 20683 16609
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 21729 16643 21787 16649
rect 21729 16640 21741 16643
rect 20956 16612 21741 16640
rect 20956 16600 20962 16612
rect 21729 16609 21741 16612
rect 21775 16609 21787 16643
rect 21729 16603 21787 16609
rect 22002 16600 22008 16652
rect 22060 16600 22066 16652
rect 22646 16600 22652 16652
rect 22704 16640 22710 16652
rect 23658 16640 23664 16652
rect 22704 16612 23664 16640
rect 22704 16600 22710 16612
rect 23658 16600 23664 16612
rect 23716 16640 23722 16652
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 23716 16612 23765 16640
rect 23716 16600 23722 16612
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 20533 16575 20591 16581
rect 20533 16541 20545 16575
rect 20579 16541 20591 16575
rect 20533 16535 20591 16541
rect 10226 16504 10232 16516
rect 7300 16476 9904 16504
rect 9968 16476 10232 16504
rect 5166 16396 5172 16448
rect 5224 16436 5230 16448
rect 7300 16436 7328 16476
rect 9968 16448 9996 16476
rect 10226 16464 10232 16476
rect 10284 16464 10290 16516
rect 22646 16464 22652 16516
rect 22704 16464 22710 16516
rect 5224 16408 7328 16436
rect 5224 16396 5230 16408
rect 8478 16396 8484 16448
rect 8536 16396 8542 16448
rect 9585 16439 9643 16445
rect 9585 16405 9597 16439
rect 9631 16436 9643 16439
rect 9950 16436 9956 16448
rect 9631 16408 9956 16436
rect 9631 16405 9643 16408
rect 9585 16399 9643 16405
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10965 16439 11023 16445
rect 10965 16405 10977 16439
rect 11011 16436 11023 16439
rect 11698 16436 11704 16448
rect 11011 16408 11704 16436
rect 11011 16405 11023 16408
rect 10965 16399 11023 16405
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 11790 16396 11796 16448
rect 11848 16396 11854 16448
rect 15286 16396 15292 16448
rect 15344 16396 15350 16448
rect 15657 16439 15715 16445
rect 15657 16405 15669 16439
rect 15703 16436 15715 16439
rect 16298 16436 16304 16448
rect 15703 16408 16304 16436
rect 15703 16405 15715 16408
rect 15657 16399 15715 16405
rect 16298 16396 16304 16408
rect 16356 16436 16362 16448
rect 16393 16439 16451 16445
rect 16393 16436 16405 16439
rect 16356 16408 16405 16436
rect 16356 16396 16362 16408
rect 16393 16405 16405 16408
rect 16439 16436 16451 16439
rect 17126 16436 17132 16448
rect 16439 16408 17132 16436
rect 16439 16405 16451 16408
rect 16393 16399 16451 16405
rect 17126 16396 17132 16408
rect 17184 16396 17190 16448
rect 17218 16396 17224 16448
rect 17276 16436 17282 16448
rect 17954 16436 17960 16448
rect 17276 16408 17960 16436
rect 17276 16396 17282 16408
rect 17954 16396 17960 16408
rect 18012 16436 18018 16448
rect 18690 16436 18696 16448
rect 18012 16408 18696 16436
rect 18012 16396 18018 16408
rect 18690 16396 18696 16408
rect 18748 16396 18754 16448
rect 20073 16439 20131 16445
rect 20073 16405 20085 16439
rect 20119 16436 20131 16439
rect 20162 16436 20168 16448
rect 20119 16408 20168 16436
rect 20119 16405 20131 16408
rect 20073 16399 20131 16405
rect 20162 16396 20168 16408
rect 20220 16396 20226 16448
rect 21174 16396 21180 16448
rect 21232 16436 21238 16448
rect 23477 16439 23535 16445
rect 23477 16436 23489 16439
rect 21232 16408 23489 16436
rect 21232 16396 21238 16408
rect 23477 16405 23489 16408
rect 23523 16405 23535 16439
rect 23477 16399 23535 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 8941 16235 8999 16241
rect 8941 16232 8953 16235
rect 7340 16204 8953 16232
rect 7340 16192 7346 16204
rect 8941 16201 8953 16204
rect 8987 16201 8999 16235
rect 8941 16195 8999 16201
rect 10137 16235 10195 16241
rect 10137 16201 10149 16235
rect 10183 16232 10195 16235
rect 10502 16232 10508 16244
rect 10183 16204 10508 16232
rect 10183 16201 10195 16204
rect 10137 16195 10195 16201
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 10597 16235 10655 16241
rect 10597 16201 10609 16235
rect 10643 16232 10655 16235
rect 11422 16232 11428 16244
rect 10643 16204 11428 16232
rect 10643 16201 10655 16204
rect 10597 16195 10655 16201
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 11701 16235 11759 16241
rect 11701 16232 11713 16235
rect 11572 16204 11713 16232
rect 11572 16192 11578 16204
rect 11701 16201 11713 16204
rect 11747 16201 11759 16235
rect 11701 16195 11759 16201
rect 12069 16235 12127 16241
rect 12069 16201 12081 16235
rect 12115 16232 12127 16235
rect 13538 16232 13544 16244
rect 12115 16204 13544 16232
rect 12115 16201 12127 16204
rect 12069 16195 12127 16201
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 13722 16192 13728 16244
rect 13780 16192 13786 16244
rect 14734 16192 14740 16244
rect 14792 16192 14798 16244
rect 17310 16192 17316 16244
rect 17368 16232 17374 16244
rect 17368 16204 18460 16232
rect 17368 16192 17374 16204
rect 2498 16124 2504 16176
rect 2556 16124 2562 16176
rect 7190 16124 7196 16176
rect 7248 16164 7254 16176
rect 9309 16167 9367 16173
rect 7248 16136 7406 16164
rect 7248 16124 7254 16136
rect 9309 16133 9321 16167
rect 9355 16164 9367 16167
rect 11790 16164 11796 16176
rect 9355 16136 11796 16164
rect 9355 16133 9367 16136
rect 9309 16127 9367 16133
rect 11790 16124 11796 16136
rect 11848 16124 11854 16176
rect 13081 16167 13139 16173
rect 13081 16133 13093 16167
rect 13127 16164 13139 16167
rect 13354 16164 13360 16176
rect 13127 16136 13360 16164
rect 13127 16133 13139 16136
rect 13081 16127 13139 16133
rect 13354 16124 13360 16136
rect 13412 16124 13418 16176
rect 14185 16167 14243 16173
rect 14185 16133 14197 16167
rect 14231 16164 14243 16167
rect 14752 16164 14780 16192
rect 14231 16136 14780 16164
rect 14231 16133 14243 16136
rect 14185 16127 14243 16133
rect 15930 16124 15936 16176
rect 15988 16164 15994 16176
rect 16393 16167 16451 16173
rect 16393 16164 16405 16167
rect 15988 16136 16405 16164
rect 15988 16124 15994 16136
rect 16393 16133 16405 16136
rect 16439 16133 16451 16167
rect 16393 16127 16451 16133
rect 17034 16124 17040 16176
rect 17092 16164 17098 16176
rect 17129 16167 17187 16173
rect 17129 16164 17141 16167
rect 17092 16136 17141 16164
rect 17092 16124 17098 16136
rect 17129 16133 17141 16136
rect 17175 16133 17187 16167
rect 17129 16127 17187 16133
rect 17218 16124 17224 16176
rect 17276 16164 17282 16176
rect 18432 16164 18460 16204
rect 18598 16192 18604 16244
rect 18656 16192 18662 16244
rect 18690 16192 18696 16244
rect 18748 16232 18754 16244
rect 18877 16235 18935 16241
rect 18877 16232 18889 16235
rect 18748 16204 18889 16232
rect 18748 16192 18754 16204
rect 18877 16201 18889 16204
rect 18923 16201 18935 16235
rect 18877 16195 18935 16201
rect 19245 16235 19303 16241
rect 19245 16201 19257 16235
rect 19291 16232 19303 16235
rect 21082 16232 21088 16244
rect 19291 16204 21088 16232
rect 19291 16201 19303 16204
rect 19245 16195 19303 16201
rect 21082 16192 21088 16204
rect 21140 16192 21146 16244
rect 17276 16136 17618 16164
rect 18432 16136 20576 16164
rect 17276 16124 17282 16136
rect 6638 16056 6644 16108
rect 6696 16056 6702 16108
rect 8404 16068 9536 16096
rect 8404 16040 8432 16068
rect 3786 15988 3792 16040
rect 3844 16028 3850 16040
rect 4062 16028 4068 16040
rect 3844 16000 4068 16028
rect 3844 15988 3850 16000
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 16028 6975 16031
rect 8294 16028 8300 16040
rect 6963 16000 8300 16028
rect 6963 15997 6975 16000
rect 6917 15991 6975 15997
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 8386 15988 8392 16040
rect 8444 15988 8450 16040
rect 9508 16037 9536 16068
rect 10318 16056 10324 16108
rect 10376 16096 10382 16108
rect 10505 16099 10563 16105
rect 10505 16096 10517 16099
rect 10376 16068 10517 16096
rect 10376 16056 10382 16068
rect 10505 16065 10517 16068
rect 10551 16065 10563 16099
rect 10505 16059 10563 16065
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12710 16096 12716 16108
rect 12207 16068 12716 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16632 16068 16865 16096
rect 16632 16056 16638 16068
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16096 19671 16099
rect 20441 16099 20499 16105
rect 20441 16096 20453 16099
rect 19659 16068 20453 16096
rect 19659 16065 19671 16068
rect 19613 16059 19671 16065
rect 20441 16065 20453 16068
rect 20487 16065 20499 16099
rect 20548 16096 20576 16136
rect 20806 16124 20812 16176
rect 20864 16164 20870 16176
rect 22465 16167 22523 16173
rect 22465 16164 22477 16167
rect 20864 16136 22477 16164
rect 20864 16124 20870 16136
rect 22465 16133 22477 16136
rect 22511 16133 22523 16167
rect 24394 16164 24400 16176
rect 22465 16127 22523 16133
rect 24136 16136 24400 16164
rect 21269 16099 21327 16105
rect 21269 16096 21281 16099
rect 20548 16068 21281 16096
rect 20441 16059 20499 16065
rect 21269 16065 21281 16068
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 22370 16056 22376 16108
rect 22428 16056 22434 16108
rect 23474 16056 23480 16108
rect 23532 16056 23538 16108
rect 24136 16105 24164 16136
rect 24394 16124 24400 16136
rect 24452 16124 24458 16176
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16065 24179 16099
rect 24121 16059 24179 16065
rect 9401 16031 9459 16037
rect 9401 15997 9413 16031
rect 9447 15997 9459 16031
rect 9401 15991 9459 15997
rect 9493 16031 9551 16037
rect 9493 15997 9505 16031
rect 9539 15997 9551 16031
rect 9493 15991 9551 15997
rect 9416 15960 9444 15991
rect 10226 15988 10232 16040
rect 10284 16028 10290 16040
rect 10689 16031 10747 16037
rect 10689 16028 10701 16031
rect 10284 16000 10701 16028
rect 10284 15988 10290 16000
rect 10689 15997 10701 16000
rect 10735 16028 10747 16031
rect 11422 16028 11428 16040
rect 10735 16000 11428 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 11422 15988 11428 16000
rect 11480 15988 11486 16040
rect 12250 15988 12256 16040
rect 12308 15988 12314 16040
rect 19702 15988 19708 16040
rect 19760 15988 19766 16040
rect 19889 16031 19947 16037
rect 19889 15997 19901 16031
rect 19935 15997 19947 16031
rect 22278 16028 22284 16040
rect 19889 15991 19947 15997
rect 20548 16000 22284 16028
rect 12066 15960 12072 15972
rect 9416 15932 12072 15960
rect 12066 15920 12072 15932
rect 12124 15920 12130 15972
rect 19904 15960 19932 15991
rect 20548 15960 20576 16000
rect 22278 15988 22284 16000
rect 22336 15988 22342 16040
rect 22554 15988 22560 16040
rect 22612 15988 22618 16040
rect 23382 15988 23388 16040
rect 23440 16028 23446 16040
rect 24397 16031 24455 16037
rect 24397 16028 24409 16031
rect 23440 16000 24409 16028
rect 23440 15988 23446 16000
rect 24397 15997 24409 16000
rect 24443 15997 24455 16031
rect 24397 15991 24455 15997
rect 19904 15932 20576 15960
rect 21453 15963 21511 15969
rect 21453 15929 21465 15963
rect 21499 15960 21511 15963
rect 23658 15960 23664 15972
rect 21499 15932 23664 15960
rect 21499 15929 21511 15932
rect 21453 15923 21511 15929
rect 23658 15920 23664 15932
rect 23716 15920 23722 15972
rect 1762 15852 1768 15904
rect 1820 15892 1826 15904
rect 2593 15895 2651 15901
rect 2593 15892 2605 15895
rect 1820 15864 2605 15892
rect 1820 15852 1826 15864
rect 2593 15861 2605 15864
rect 2639 15861 2651 15895
rect 2593 15855 2651 15861
rect 14274 15852 14280 15904
rect 14332 15852 14338 15904
rect 15562 15852 15568 15904
rect 15620 15892 15626 15904
rect 16025 15895 16083 15901
rect 16025 15892 16037 15895
rect 15620 15864 16037 15892
rect 15620 15852 15626 15864
rect 16025 15861 16037 15864
rect 16071 15861 16083 15895
rect 16025 15855 16083 15861
rect 22005 15895 22063 15901
rect 22005 15861 22017 15895
rect 22051 15892 22063 15895
rect 22186 15892 22192 15904
rect 22051 15864 22192 15892
rect 22051 15861 22063 15864
rect 22005 15855 22063 15861
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 22462 15852 22468 15904
rect 22520 15892 22526 15904
rect 23293 15895 23351 15901
rect 23293 15892 23305 15895
rect 22520 15864 23305 15892
rect 22520 15852 22526 15864
rect 23293 15861 23305 15864
rect 23339 15861 23351 15895
rect 23293 15855 23351 15861
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 8754 15648 8760 15700
rect 8812 15648 8818 15700
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10134 15688 10140 15700
rect 10008 15660 10140 15688
rect 10008 15648 10014 15660
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 11756 15660 14289 15688
rect 11756 15648 11762 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 21085 15691 21143 15697
rect 21085 15688 21097 15691
rect 14277 15651 14335 15657
rect 19996 15660 21097 15688
rect 17313 15623 17371 15629
rect 17313 15589 17325 15623
rect 17359 15620 17371 15623
rect 19886 15620 19892 15632
rect 17359 15592 19892 15620
rect 17359 15589 17371 15592
rect 17313 15583 17371 15589
rect 19886 15580 19892 15592
rect 19944 15580 19950 15632
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15552 11115 15555
rect 11330 15552 11336 15564
rect 11103 15524 11336 15552
rect 11103 15521 11115 15524
rect 11057 15515 11115 15521
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 11422 15512 11428 15564
rect 11480 15552 11486 15564
rect 14182 15552 14188 15564
rect 11480 15524 14188 15552
rect 11480 15512 11486 15524
rect 14182 15512 14188 15524
rect 14240 15552 14246 15564
rect 14829 15555 14887 15561
rect 14829 15552 14841 15555
rect 14240 15524 14841 15552
rect 14240 15512 14246 15524
rect 14829 15521 14841 15524
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 17402 15512 17408 15564
rect 17460 15552 17466 15564
rect 17865 15555 17923 15561
rect 17865 15552 17877 15555
rect 17460 15524 17877 15552
rect 17460 15512 17466 15524
rect 17865 15521 17877 15524
rect 17911 15521 17923 15555
rect 19996 15552 20024 15660
rect 21085 15657 21097 15660
rect 21131 15657 21143 15691
rect 21085 15651 21143 15657
rect 20990 15580 20996 15632
rect 21048 15620 21054 15632
rect 21048 15592 21864 15620
rect 21048 15580 21054 15592
rect 17865 15515 17923 15521
rect 19904 15524 20024 15552
rect 20073 15555 20131 15561
rect 13354 15484 13360 15496
rect 12466 15470 13360 15484
rect 12452 15456 13360 15470
rect 11333 15419 11391 15425
rect 11333 15385 11345 15419
rect 11379 15385 11391 15419
rect 11333 15379 11391 15385
rect 8478 15308 8484 15360
rect 8536 15308 8542 15360
rect 10229 15351 10287 15357
rect 10229 15317 10241 15351
rect 10275 15348 10287 15351
rect 10318 15348 10324 15360
rect 10275 15320 10324 15348
rect 10275 15317 10287 15320
rect 10229 15311 10287 15317
rect 10318 15308 10324 15320
rect 10376 15308 10382 15360
rect 10781 15351 10839 15357
rect 10781 15317 10793 15351
rect 10827 15348 10839 15351
rect 10870 15348 10876 15360
rect 10827 15320 10876 15348
rect 10827 15317 10839 15320
rect 10781 15311 10839 15317
rect 10870 15308 10876 15320
rect 10928 15348 10934 15360
rect 11348 15348 11376 15379
rect 11974 15348 11980 15360
rect 10928 15320 11980 15348
rect 10928 15308 10934 15320
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12250 15308 12256 15360
rect 12308 15348 12314 15360
rect 12452 15348 12480 15456
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 13449 15487 13507 15493
rect 13449 15453 13461 15487
rect 13495 15484 13507 15487
rect 13722 15484 13728 15496
rect 13495 15456 13728 15484
rect 13495 15453 13507 15456
rect 13449 15447 13507 15453
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15484 14703 15487
rect 15286 15484 15292 15496
rect 14691 15456 15292 15484
rect 14691 15453 14703 15456
rect 14645 15447 14703 15453
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 17678 15444 17684 15496
rect 17736 15484 17742 15496
rect 19904 15493 19932 15524
rect 20073 15521 20085 15555
rect 20119 15552 20131 15555
rect 21174 15552 21180 15564
rect 20119 15524 21180 15552
rect 20119 15521 20131 15524
rect 20073 15515 20131 15521
rect 21174 15512 21180 15524
rect 21232 15512 21238 15564
rect 19889 15487 19947 15493
rect 19889 15484 19901 15487
rect 17736 15456 19901 15484
rect 17736 15444 17742 15456
rect 19889 15453 19901 15456
rect 19935 15453 19947 15487
rect 19889 15447 19947 15453
rect 20809 15487 20867 15493
rect 20809 15453 20821 15487
rect 20855 15484 20867 15487
rect 21266 15484 21272 15496
rect 20855 15456 21272 15484
rect 20855 15453 20867 15456
rect 20809 15447 20867 15453
rect 21266 15444 21272 15456
rect 21324 15444 21330 15496
rect 21836 15493 21864 15592
rect 21821 15487 21879 15493
rect 21821 15453 21833 15487
rect 21867 15453 21879 15487
rect 21821 15447 21879 15453
rect 22833 15487 22891 15493
rect 22833 15453 22845 15487
rect 22879 15484 22891 15487
rect 24210 15484 24216 15496
rect 22879 15456 24216 15484
rect 22879 15453 22891 15456
rect 22833 15447 22891 15453
rect 24210 15444 24216 15456
rect 24268 15444 24274 15496
rect 12618 15376 12624 15428
rect 12676 15416 12682 15428
rect 13633 15419 13691 15425
rect 13633 15416 13645 15419
rect 12676 15388 13645 15416
rect 12676 15376 12682 15388
rect 13633 15385 13645 15388
rect 13679 15385 13691 15419
rect 13633 15379 13691 15385
rect 15470 15376 15476 15428
rect 15528 15416 15534 15428
rect 17773 15419 17831 15425
rect 17773 15416 17785 15419
rect 15528 15388 17785 15416
rect 15528 15376 15534 15388
rect 17773 15385 17785 15388
rect 17819 15416 17831 15419
rect 18325 15419 18383 15425
rect 18325 15416 18337 15419
rect 17819 15388 18337 15416
rect 17819 15385 17831 15388
rect 17773 15379 17831 15385
rect 18325 15385 18337 15388
rect 18371 15385 18383 15419
rect 21542 15416 21548 15428
rect 18325 15379 18383 15385
rect 19444 15388 21548 15416
rect 12308 15320 12480 15348
rect 12308 15308 12314 15320
rect 12802 15308 12808 15360
rect 12860 15308 12866 15360
rect 14737 15351 14795 15357
rect 14737 15317 14749 15351
rect 14783 15348 14795 15351
rect 15654 15348 15660 15360
rect 14783 15320 15660 15348
rect 14783 15317 14795 15320
rect 14737 15311 14795 15317
rect 15654 15308 15660 15320
rect 15712 15308 15718 15360
rect 16758 15308 16764 15360
rect 16816 15348 16822 15360
rect 17037 15351 17095 15357
rect 17037 15348 17049 15351
rect 16816 15320 17049 15348
rect 16816 15308 16822 15320
rect 17037 15317 17049 15320
rect 17083 15348 17095 15351
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 17083 15320 17693 15348
rect 17083 15317 17095 15320
rect 17037 15311 17095 15317
rect 17681 15317 17693 15320
rect 17727 15317 17739 15351
rect 17681 15311 17739 15317
rect 18690 15308 18696 15360
rect 18748 15308 18754 15360
rect 19444 15357 19472 15388
rect 21542 15376 21548 15388
rect 21600 15376 21606 15428
rect 23845 15419 23903 15425
rect 23845 15385 23857 15419
rect 23891 15416 23903 15419
rect 24946 15416 24952 15428
rect 23891 15388 24952 15416
rect 23891 15385 23903 15388
rect 23845 15379 23903 15385
rect 24946 15376 24952 15388
rect 25004 15376 25010 15428
rect 19429 15351 19487 15357
rect 19429 15317 19441 15351
rect 19475 15317 19487 15351
rect 19429 15311 19487 15317
rect 19702 15308 19708 15360
rect 19760 15348 19766 15360
rect 19797 15351 19855 15357
rect 19797 15348 19809 15351
rect 19760 15320 19809 15348
rect 19760 15308 19766 15320
rect 19797 15317 19809 15320
rect 19843 15317 19855 15351
rect 19797 15311 19855 15317
rect 20622 15308 20628 15360
rect 20680 15308 20686 15360
rect 21910 15308 21916 15360
rect 21968 15308 21974 15360
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 8754 15104 8760 15156
rect 8812 15144 8818 15156
rect 9582 15144 9588 15156
rect 8812 15116 9588 15144
rect 8812 15104 8818 15116
rect 9582 15104 9588 15116
rect 9640 15144 9646 15156
rect 9640 15116 10732 15144
rect 9640 15104 9646 15116
rect 9398 15036 9404 15088
rect 9456 15036 9462 15088
rect 10704 15076 10732 15116
rect 12158 15104 12164 15156
rect 12216 15144 12222 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12216 15116 13001 15144
rect 12216 15104 12222 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 14185 15147 14243 15153
rect 14185 15113 14197 15147
rect 14231 15144 14243 15147
rect 17310 15144 17316 15156
rect 14231 15116 17316 15144
rect 14231 15113 14243 15116
rect 14185 15107 14243 15113
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 18748 15116 18797 15144
rect 18748 15104 18754 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 18785 15107 18843 15113
rect 18874 15104 18880 15156
rect 18932 15104 18938 15156
rect 22281 15147 22339 15153
rect 22281 15113 22293 15147
rect 22327 15144 22339 15147
rect 22370 15144 22376 15156
rect 22327 15116 22376 15144
rect 22327 15113 22339 15116
rect 22281 15107 22339 15113
rect 22370 15104 22376 15116
rect 22428 15104 22434 15156
rect 11609 15079 11667 15085
rect 11609 15076 11621 15079
rect 10626 15048 11621 15076
rect 11609 15045 11621 15048
rect 11655 15076 11667 15079
rect 12250 15076 12256 15088
rect 11655 15048 12256 15076
rect 11655 15045 11667 15048
rect 11609 15039 11667 15045
rect 12250 15036 12256 15048
rect 12308 15036 12314 15088
rect 13357 15079 13415 15085
rect 13357 15045 13369 15079
rect 13403 15076 13415 15079
rect 15378 15076 15384 15088
rect 13403 15048 15384 15076
rect 13403 15045 13415 15048
rect 13357 15039 13415 15045
rect 15378 15036 15384 15048
rect 15436 15036 15442 15088
rect 15657 15079 15715 15085
rect 15657 15045 15669 15079
rect 15703 15076 15715 15079
rect 16114 15076 16120 15088
rect 15703 15048 16120 15076
rect 15703 15045 15715 15048
rect 15657 15039 15715 15045
rect 16114 15036 16120 15048
rect 16172 15036 16178 15088
rect 16298 15036 16304 15088
rect 16356 15076 16362 15088
rect 19702 15076 19708 15088
rect 16356 15048 19708 15076
rect 16356 15036 16362 15048
rect 19702 15036 19708 15048
rect 19760 15076 19766 15088
rect 20073 15079 20131 15085
rect 20073 15076 20085 15079
rect 19760 15048 20085 15076
rect 19760 15036 19766 15048
rect 20073 15045 20085 15048
rect 20119 15045 20131 15079
rect 20073 15039 20131 15045
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 12492 14980 13584 15008
rect 12492 14968 12498 14980
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14909 9183 14943
rect 9125 14903 9183 14909
rect 9140 14804 9168 14903
rect 10870 14900 10876 14952
rect 10928 14940 10934 14952
rect 13556 14949 13584 14980
rect 14550 14968 14556 15020
rect 14608 14968 14614 15020
rect 14645 15011 14703 15017
rect 14645 14977 14657 15011
rect 14691 15008 14703 15011
rect 15289 15011 15347 15017
rect 15289 15008 15301 15011
rect 14691 14980 15301 15008
rect 14691 14977 14703 14980
rect 14645 14971 14703 14977
rect 15289 14977 15301 14980
rect 15335 15008 15347 15011
rect 15470 15008 15476 15020
rect 15335 14980 15476 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 16758 14968 16764 15020
rect 16816 14968 16822 15020
rect 16942 14968 16948 15020
rect 17000 15008 17006 15020
rect 17221 15011 17279 15017
rect 17221 15008 17233 15011
rect 17000 14980 17233 15008
rect 17000 14968 17006 14980
rect 17221 14977 17233 14980
rect 17267 15008 17279 15011
rect 17681 15011 17739 15017
rect 17681 15008 17693 15011
rect 17267 14980 17693 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 17681 14977 17693 14980
rect 17727 14977 17739 15011
rect 17681 14971 17739 14977
rect 18598 14968 18604 15020
rect 18656 15008 18662 15020
rect 18656 14980 19012 15008
rect 18656 14968 18662 14980
rect 11149 14943 11207 14949
rect 11149 14940 11161 14943
rect 10928 14912 11161 14940
rect 10928 14900 10934 14912
rect 11149 14909 11161 14912
rect 11195 14909 11207 14943
rect 11149 14903 11207 14909
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 12713 14875 12771 14881
rect 12713 14841 12725 14875
rect 12759 14872 12771 14875
rect 13464 14872 13492 14903
rect 14826 14900 14832 14952
rect 14884 14900 14890 14952
rect 16776 14940 16804 14968
rect 14936 14912 16804 14940
rect 13630 14872 13636 14884
rect 12759 14844 13636 14872
rect 12759 14841 12771 14844
rect 12713 14835 12771 14841
rect 13630 14832 13636 14844
rect 13688 14872 13694 14884
rect 14936 14872 14964 14912
rect 17862 14900 17868 14952
rect 17920 14940 17926 14952
rect 18782 14940 18788 14952
rect 17920 14912 18788 14940
rect 17920 14900 17926 14912
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 18984 14949 19012 14980
rect 19794 14968 19800 15020
rect 19852 14968 19858 15020
rect 23385 15011 23443 15017
rect 23385 14977 23397 15011
rect 23431 15008 23443 15011
rect 23566 15008 23572 15020
rect 23431 14980 23572 15008
rect 23431 14977 23443 14980
rect 23385 14971 23443 14977
rect 23566 14968 23572 14980
rect 23624 14968 23630 15020
rect 24118 14968 24124 15020
rect 24176 14968 24182 15020
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14909 19027 14943
rect 18969 14903 19027 14909
rect 24762 14900 24768 14952
rect 24820 14900 24826 14952
rect 13688 14844 14964 14872
rect 17405 14875 17463 14881
rect 13688 14832 13694 14844
rect 17405 14841 17417 14875
rect 17451 14872 17463 14875
rect 17586 14872 17592 14884
rect 17451 14844 17592 14872
rect 17451 14841 17463 14844
rect 17405 14835 17463 14841
rect 17586 14832 17592 14844
rect 17644 14832 17650 14884
rect 9950 14804 9956 14816
rect 9140 14776 9956 14804
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 15749 14807 15807 14813
rect 15749 14773 15761 14807
rect 15795 14804 15807 14807
rect 16666 14804 16672 14816
rect 15795 14776 16672 14804
rect 15795 14773 15807 14776
rect 15749 14767 15807 14773
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 18417 14807 18475 14813
rect 18417 14773 18429 14807
rect 18463 14804 18475 14807
rect 18874 14804 18880 14816
rect 18463 14776 18880 14804
rect 18463 14773 18475 14776
rect 18417 14767 18475 14773
rect 18874 14764 18880 14776
rect 18932 14764 18938 14816
rect 19613 14807 19671 14813
rect 19613 14773 19625 14807
rect 19659 14804 19671 14807
rect 19794 14804 19800 14816
rect 19659 14776 19800 14804
rect 19659 14773 19671 14776
rect 19613 14767 19671 14773
rect 19794 14764 19800 14776
rect 19852 14764 19858 14816
rect 21266 14764 21272 14816
rect 21324 14804 21330 14816
rect 23201 14807 23259 14813
rect 23201 14804 23213 14807
rect 21324 14776 23213 14804
rect 21324 14764 21330 14776
rect 23201 14773 23213 14776
rect 23247 14773 23259 14807
rect 23201 14767 23259 14773
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 10410 14560 10416 14612
rect 10468 14600 10474 14612
rect 10686 14600 10692 14612
rect 10468 14572 10692 14600
rect 10468 14560 10474 14572
rect 10686 14560 10692 14572
rect 10744 14600 10750 14612
rect 10744 14572 12434 14600
rect 10744 14560 10750 14572
rect 11330 14492 11336 14544
rect 11388 14492 11394 14544
rect 12069 14535 12127 14541
rect 12069 14501 12081 14535
rect 12115 14532 12127 14535
rect 12250 14532 12256 14544
rect 12115 14504 12256 14532
rect 12115 14501 12127 14504
rect 12069 14495 12127 14501
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 11348 14464 11376 14492
rect 10008 14436 11376 14464
rect 10008 14424 10014 14436
rect 11974 14396 11980 14408
rect 11362 14368 11980 14396
rect 11974 14356 11980 14368
rect 12032 14396 12038 14408
rect 12084 14396 12112 14495
rect 12250 14492 12256 14504
rect 12308 14492 12314 14544
rect 12406 14532 12434 14572
rect 12710 14560 12716 14612
rect 12768 14600 12774 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12768 14572 13001 14600
rect 12768 14560 12774 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 14369 14603 14427 14609
rect 14369 14569 14381 14603
rect 14415 14600 14427 14603
rect 14461 14603 14519 14609
rect 14461 14600 14473 14603
rect 14415 14572 14473 14600
rect 14415 14569 14427 14572
rect 14369 14563 14427 14569
rect 14461 14569 14473 14572
rect 14507 14600 14519 14603
rect 15378 14600 15384 14612
rect 14507 14572 15384 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 14093 14535 14151 14541
rect 14093 14532 14105 14535
rect 12406 14504 14105 14532
rect 14093 14501 14105 14504
rect 14139 14532 14151 14535
rect 14550 14532 14556 14544
rect 14139 14504 14556 14532
rect 14139 14501 14151 14504
rect 14093 14495 14151 14501
rect 14550 14492 14556 14504
rect 14608 14492 14614 14544
rect 12713 14467 12771 14473
rect 12713 14433 12725 14467
rect 12759 14464 12771 14467
rect 13541 14467 13599 14473
rect 13541 14464 13553 14467
rect 12759 14436 13553 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 13541 14433 13553 14436
rect 13587 14464 13599 14467
rect 14458 14464 14464 14476
rect 13587 14436 14464 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 12032 14368 12112 14396
rect 13357 14399 13415 14405
rect 12032 14356 12038 14368
rect 13357 14365 13369 14399
rect 13403 14396 13415 14399
rect 14660 14396 14688 14572
rect 15378 14560 15384 14572
rect 15436 14600 15442 14612
rect 15838 14600 15844 14612
rect 15436 14572 15844 14600
rect 15436 14560 15442 14572
rect 15838 14560 15844 14572
rect 15896 14560 15902 14612
rect 17034 14560 17040 14612
rect 17092 14600 17098 14612
rect 17129 14603 17187 14609
rect 17129 14600 17141 14603
rect 17092 14572 17141 14600
rect 17092 14560 17098 14572
rect 17129 14569 17141 14572
rect 17175 14569 17187 14603
rect 17129 14563 17187 14569
rect 18693 14603 18751 14609
rect 18693 14569 18705 14603
rect 18739 14600 18751 14603
rect 21634 14600 21640 14612
rect 18739 14572 21640 14600
rect 18739 14569 18751 14572
rect 18693 14563 18751 14569
rect 21634 14560 21640 14572
rect 21692 14560 21698 14612
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 16390 14464 16396 14476
rect 15436 14436 16396 14464
rect 15436 14424 15442 14436
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 17126 14424 17132 14476
rect 17184 14464 17190 14476
rect 20806 14464 20812 14476
rect 17184 14436 20812 14464
rect 17184 14424 17190 14436
rect 20806 14424 20812 14436
rect 20864 14424 20870 14476
rect 21174 14424 21180 14476
rect 21232 14424 21238 14476
rect 13403 14368 14688 14396
rect 18233 14399 18291 14405
rect 13403 14365 13415 14368
rect 13357 14359 13415 14365
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 18506 14396 18512 14408
rect 18279 14368 18512 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18506 14356 18512 14368
rect 18564 14396 18570 14408
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 18564 14368 18613 14396
rect 18564 14356 18570 14368
rect 18601 14365 18613 14368
rect 18647 14365 18659 14399
rect 18601 14359 18659 14365
rect 20898 14356 20904 14408
rect 20956 14356 20962 14408
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 22646 14396 22652 14408
rect 22336 14368 22652 14396
rect 22336 14356 22342 14368
rect 22646 14356 22652 14368
rect 22704 14396 22710 14408
rect 22925 14399 22983 14405
rect 22925 14396 22937 14399
rect 22704 14368 22937 14396
rect 22704 14356 22710 14368
rect 22925 14365 22937 14368
rect 22971 14365 22983 14399
rect 22925 14359 22983 14365
rect 10226 14288 10232 14340
rect 10284 14288 10290 14340
rect 12526 14288 12532 14340
rect 12584 14328 12590 14340
rect 13449 14331 13507 14337
rect 13449 14328 13461 14331
rect 12584 14300 13461 14328
rect 12584 14288 12590 14300
rect 13449 14297 13461 14300
rect 13495 14328 13507 14331
rect 13630 14328 13636 14340
rect 13495 14300 13636 14328
rect 13495 14297 13507 14300
rect 13449 14291 13507 14297
rect 13630 14288 13636 14300
rect 13688 14288 13694 14340
rect 15657 14331 15715 14337
rect 15657 14297 15669 14331
rect 15703 14328 15715 14331
rect 15930 14328 15936 14340
rect 15703 14300 15936 14328
rect 15703 14297 15715 14300
rect 15657 14291 15715 14297
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 16040 14300 16146 14328
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 10962 14260 10968 14272
rect 9916 14232 10968 14260
rect 9916 14220 9922 14232
rect 10962 14220 10968 14232
rect 11020 14260 11026 14272
rect 11701 14263 11759 14269
rect 11701 14260 11713 14263
rect 11020 14232 11713 14260
rect 11020 14220 11026 14232
rect 11701 14229 11713 14232
rect 11747 14229 11759 14263
rect 11701 14223 11759 14229
rect 15746 14220 15752 14272
rect 15804 14260 15810 14272
rect 16040 14260 16068 14300
rect 17218 14260 17224 14272
rect 15804 14232 17224 14260
rect 15804 14220 15810 14232
rect 17218 14220 17224 14232
rect 17276 14260 17282 14272
rect 17405 14263 17463 14269
rect 17405 14260 17417 14263
rect 17276 14232 17417 14260
rect 17276 14220 17282 14232
rect 17405 14229 17417 14232
rect 17451 14229 17463 14263
rect 17405 14223 17463 14229
rect 19426 14220 19432 14272
rect 19484 14220 19490 14272
rect 19702 14220 19708 14272
rect 19760 14260 19766 14272
rect 19981 14263 20039 14269
rect 19981 14260 19993 14263
rect 19760 14232 19993 14260
rect 19760 14220 19766 14232
rect 19981 14229 19993 14232
rect 20027 14229 20039 14263
rect 19981 14223 20039 14229
rect 21818 14220 21824 14272
rect 21876 14260 21882 14272
rect 22649 14263 22707 14269
rect 22649 14260 22661 14263
rect 21876 14232 22661 14260
rect 21876 14220 21882 14232
rect 22649 14229 22661 14232
rect 22695 14229 22707 14263
rect 22649 14223 22707 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 9950 14056 9956 14068
rect 8128 14028 9956 14056
rect 8128 13988 8156 14028
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10318 14056 10324 14068
rect 10192 14028 10324 14056
rect 10192 14016 10198 14028
rect 10318 14016 10324 14028
rect 10376 14056 10382 14068
rect 11885 14059 11943 14065
rect 11885 14056 11897 14059
rect 10376 14028 11897 14056
rect 10376 14016 10382 14028
rect 11885 14025 11897 14028
rect 11931 14025 11943 14059
rect 11885 14019 11943 14025
rect 9582 13988 9588 14000
rect 8036 13960 8156 13988
rect 9522 13960 9588 13988
rect 1762 13880 1768 13932
rect 1820 13880 1826 13932
rect 8036 13929 8064 13960
rect 9582 13948 9588 13960
rect 9640 13988 9646 14000
rect 10045 13991 10103 13997
rect 10045 13988 10057 13991
rect 9640 13960 10057 13988
rect 9640 13948 9646 13960
rect 10045 13957 10057 13960
rect 10091 13957 10103 13991
rect 10045 13951 10103 13957
rect 8021 13923 8079 13929
rect 8021 13889 8033 13923
rect 8067 13889 8079 13923
rect 8021 13883 8079 13889
rect 10318 13880 10324 13932
rect 10376 13920 10382 13932
rect 10594 13920 10600 13932
rect 10376 13892 10600 13920
rect 10376 13880 10382 13892
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 11900 13920 11928 14019
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 12713 14059 12771 14065
rect 12713 14056 12725 14059
rect 12492 14028 12725 14056
rect 12492 14016 12498 14028
rect 12713 14025 12725 14028
rect 12759 14025 12771 14059
rect 12713 14019 12771 14025
rect 17218 14016 17224 14068
rect 17276 14056 17282 14068
rect 17276 14028 17540 14056
rect 17276 14016 17282 14028
rect 13538 13948 13544 14000
rect 13596 13988 13602 14000
rect 14001 13991 14059 13997
rect 14001 13988 14013 13991
rect 13596 13960 14013 13988
rect 13596 13948 13602 13960
rect 14001 13957 14013 13960
rect 14047 13957 14059 13991
rect 14001 13951 14059 13957
rect 17402 13948 17408 14000
rect 17460 13948 17466 14000
rect 17512 13988 17540 14028
rect 18414 14016 18420 14068
rect 18472 14056 18478 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 18472 14028 18889 14056
rect 18472 14016 18478 14028
rect 18877 14025 18889 14028
rect 18923 14056 18935 14059
rect 19242 14056 19248 14068
rect 18923 14028 19248 14056
rect 18923 14025 18935 14028
rect 18877 14019 18935 14025
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 19797 14059 19855 14065
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 22370 14056 22376 14068
rect 19843 14028 22376 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 22370 14016 22376 14028
rect 22428 14016 22434 14068
rect 22646 14016 22652 14068
rect 22704 14056 22710 14068
rect 23017 14059 23075 14065
rect 23017 14056 23029 14059
rect 22704 14028 23029 14056
rect 22704 14016 22710 14028
rect 23017 14025 23029 14028
rect 23063 14025 23075 14059
rect 23017 14019 23075 14025
rect 17862 13988 17868 14000
rect 17512 13960 17868 13988
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 19702 13948 19708 14000
rect 19760 13948 19766 14000
rect 19978 13948 19984 14000
rect 20036 13988 20042 14000
rect 21177 13991 21235 13997
rect 21177 13988 21189 13991
rect 20036 13960 21189 13988
rect 20036 13948 20042 13960
rect 21177 13957 21189 13960
rect 21223 13988 21235 13991
rect 21821 13991 21879 13997
rect 21821 13988 21833 13991
rect 21223 13960 21833 13988
rect 21223 13957 21235 13960
rect 21177 13951 21235 13957
rect 21821 13957 21833 13960
rect 21867 13957 21879 13991
rect 21821 13951 21879 13957
rect 12621 13923 12679 13929
rect 12621 13920 12633 13923
rect 11900 13892 12633 13920
rect 12621 13889 12633 13892
rect 12667 13889 12679 13923
rect 12621 13883 12679 13889
rect 16574 13880 16580 13932
rect 16632 13920 16638 13932
rect 17126 13920 17132 13932
rect 16632 13892 17132 13920
rect 16632 13880 16638 13892
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 20254 13880 20260 13932
rect 20312 13920 20318 13932
rect 20441 13923 20499 13929
rect 20441 13920 20453 13923
rect 20312 13892 20453 13920
rect 20312 13880 20318 13892
rect 20441 13889 20453 13892
rect 20487 13920 20499 13923
rect 20714 13920 20720 13932
rect 20487 13892 20720 13920
rect 20487 13889 20499 13892
rect 20441 13883 20499 13889
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 22738 13880 22744 13932
rect 22796 13920 22802 13932
rect 23201 13923 23259 13929
rect 23201 13920 23213 13923
rect 22796 13892 23213 13920
rect 22796 13880 22802 13892
rect 23201 13889 23213 13892
rect 23247 13889 23259 13923
rect 23201 13883 23259 13889
rect 23842 13880 23848 13932
rect 23900 13920 23906 13932
rect 23937 13923 23995 13929
rect 23937 13920 23949 13923
rect 23900 13892 23949 13920
rect 23900 13880 23906 13892
rect 23937 13889 23949 13892
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 9769 13855 9827 13861
rect 9769 13852 9781 13855
rect 9548 13824 9781 13852
rect 9548 13812 9554 13824
rect 9769 13821 9781 13824
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 12805 13855 12863 13861
rect 12805 13821 12817 13855
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 11790 13744 11796 13796
rect 11848 13784 11854 13796
rect 12820 13784 12848 13815
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 13725 13855 13783 13861
rect 13725 13852 13737 13855
rect 13688 13824 13737 13852
rect 13688 13812 13694 13824
rect 13725 13821 13737 13824
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 17402 13812 17408 13864
rect 17460 13852 17466 13864
rect 19334 13852 19340 13864
rect 17460 13824 19340 13852
rect 17460 13812 17466 13824
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 20346 13812 20352 13864
rect 20404 13852 20410 13864
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20404 13824 20637 13852
rect 20404 13812 20410 13824
rect 20625 13821 20637 13824
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 21361 13855 21419 13861
rect 21361 13821 21373 13855
rect 21407 13852 21419 13855
rect 22094 13852 22100 13864
rect 21407 13824 22100 13852
rect 21407 13821 21419 13824
rect 21361 13815 21419 13821
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 24670 13812 24676 13864
rect 24728 13812 24734 13864
rect 11848 13756 12848 13784
rect 11848 13744 11854 13756
rect 13538 13744 13544 13796
rect 13596 13784 13602 13796
rect 14274 13784 14280 13796
rect 13596 13756 14280 13784
rect 13596 13744 13602 13756
rect 14274 13744 14280 13756
rect 14332 13744 14338 13796
rect 8284 13719 8342 13725
rect 8284 13685 8296 13719
rect 8330 13716 8342 13719
rect 9858 13716 9864 13728
rect 8330 13688 9864 13716
rect 8330 13685 8342 13688
rect 8284 13679 8342 13685
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 12253 13719 12311 13725
rect 12253 13685 12265 13719
rect 12299 13716 12311 13719
rect 15102 13716 15108 13728
rect 12299 13688 15108 13716
rect 12299 13685 12311 13688
rect 12253 13679 12311 13685
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 17862 13676 17868 13728
rect 17920 13716 17926 13728
rect 19153 13719 19211 13725
rect 19153 13716 19165 13719
rect 17920 13688 19165 13716
rect 17920 13676 17926 13688
rect 19153 13685 19165 13688
rect 19199 13685 19211 13719
rect 19153 13679 19211 13685
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 5868 13484 9996 13512
rect 5868 13472 5874 13484
rect 9033 13447 9091 13453
rect 9033 13413 9045 13447
rect 9079 13444 9091 13447
rect 9582 13444 9588 13456
rect 9079 13416 9588 13444
rect 9079 13413 9091 13416
rect 9033 13407 9091 13413
rect 8478 13376 8484 13388
rect 6840 13348 8484 13376
rect 6840 13320 6868 13348
rect 8478 13336 8484 13348
rect 8536 13376 8542 13388
rect 9125 13379 9183 13385
rect 9125 13376 9137 13379
rect 8536 13348 9137 13376
rect 8536 13336 8542 13348
rect 9125 13345 9137 13348
rect 9171 13345 9183 13379
rect 9125 13339 9183 13345
rect 6822 13268 6828 13320
rect 6880 13268 6886 13320
rect 8386 13308 8392 13320
rect 8234 13280 8392 13308
rect 8386 13268 8392 13280
rect 8444 13308 8450 13320
rect 9232 13308 9260 13416
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 9858 13336 9864 13388
rect 9916 13336 9922 13388
rect 9968 13376 9996 13484
rect 11606 13472 11612 13524
rect 11664 13472 11670 13524
rect 11974 13472 11980 13524
rect 12032 13472 12038 13524
rect 12066 13472 12072 13524
rect 12124 13512 12130 13524
rect 12345 13515 12403 13521
rect 12345 13512 12357 13515
rect 12124 13484 12357 13512
rect 12124 13472 12130 13484
rect 12345 13481 12357 13484
rect 12391 13481 12403 13515
rect 12345 13475 12403 13481
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 13357 13515 13415 13521
rect 13357 13512 13369 13515
rect 12492 13484 13369 13512
rect 12492 13472 12498 13484
rect 13357 13481 13369 13484
rect 13403 13512 13415 13515
rect 13403 13484 15884 13512
rect 13403 13481 13415 13484
rect 13357 13475 13415 13481
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 9968 13348 10149 13376
rect 10137 13345 10149 13348
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 12897 13379 12955 13385
rect 12897 13376 12909 13379
rect 12860 13348 12909 13376
rect 12860 13336 12866 13348
rect 12897 13345 12909 13348
rect 12943 13345 12955 13379
rect 12897 13339 12955 13345
rect 14553 13379 14611 13385
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15378 13376 15384 13388
rect 14599 13348 15384 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 15856 13376 15884 13484
rect 15930 13472 15936 13524
rect 15988 13512 15994 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 15988 13484 16313 13512
rect 15988 13472 15994 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 19242 13472 19248 13524
rect 19300 13512 19306 13524
rect 19300 13484 20024 13512
rect 19300 13472 19306 13484
rect 17773 13447 17831 13453
rect 17773 13413 17785 13447
rect 17819 13444 17831 13447
rect 19334 13444 19340 13456
rect 17819 13416 19340 13444
rect 17819 13413 17831 13416
rect 17773 13407 17831 13413
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 15856 13348 18245 13376
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 18417 13379 18475 13385
rect 18417 13345 18429 13379
rect 18463 13376 18475 13379
rect 18506 13376 18512 13388
rect 18463 13348 18512 13376
rect 18463 13345 18475 13348
rect 18417 13339 18475 13345
rect 8444 13280 9260 13308
rect 12713 13311 12771 13317
rect 8444 13268 8450 13280
rect 12713 13277 12725 13311
rect 12759 13308 12771 13311
rect 14458 13308 14464 13320
rect 12759 13280 14464 13308
rect 12759 13277 12771 13280
rect 12713 13271 12771 13277
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 18248 13308 18276 13339
rect 18506 13336 18512 13348
rect 18564 13376 18570 13388
rect 19996 13385 20024 13484
rect 20714 13472 20720 13524
rect 20772 13472 20778 13524
rect 22278 13512 22284 13524
rect 21560 13484 22284 13512
rect 19981 13379 20039 13385
rect 18564 13348 19932 13376
rect 18564 13336 18570 13348
rect 18785 13311 18843 13317
rect 18785 13308 18797 13311
rect 18248 13280 18797 13308
rect 18785 13277 18797 13280
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19797 13311 19855 13317
rect 19797 13308 19809 13311
rect 19484 13280 19809 13308
rect 19484 13268 19490 13280
rect 19797 13277 19809 13280
rect 19843 13277 19855 13311
rect 19904 13308 19932 13348
rect 19981 13345 19993 13379
rect 20027 13345 20039 13379
rect 19981 13339 20039 13345
rect 20990 13308 20996 13320
rect 19904 13280 20996 13308
rect 19797 13271 19855 13277
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 7098 13200 7104 13252
rect 7156 13200 7162 13252
rect 11514 13240 11520 13252
rect 11362 13212 11520 13240
rect 11514 13200 11520 13212
rect 11572 13240 11578 13252
rect 11974 13240 11980 13252
rect 11572 13212 11980 13240
rect 11572 13200 11578 13212
rect 11974 13200 11980 13212
rect 12032 13200 12038 13252
rect 12805 13243 12863 13249
rect 12805 13209 12817 13243
rect 12851 13240 12863 13243
rect 13998 13240 14004 13252
rect 12851 13212 14004 13240
rect 12851 13209 12863 13212
rect 12805 13203 12863 13209
rect 13998 13200 14004 13212
rect 14056 13200 14062 13252
rect 14550 13200 14556 13252
rect 14608 13240 14614 13252
rect 14826 13240 14832 13252
rect 14608 13212 14832 13240
rect 14608 13200 14614 13212
rect 14826 13200 14832 13212
rect 14884 13200 14890 13252
rect 15286 13200 15292 13252
rect 15344 13200 15350 13252
rect 16114 13200 16120 13252
rect 16172 13240 16178 13252
rect 16172 13212 17540 13240
rect 16172 13200 16178 13212
rect 8573 13175 8631 13181
rect 8573 13141 8585 13175
rect 8619 13172 8631 13175
rect 8754 13172 8760 13184
rect 8619 13144 8760 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 8754 13132 8760 13144
rect 8812 13132 8818 13184
rect 16853 13175 16911 13181
rect 16853 13141 16865 13175
rect 16899 13172 16911 13175
rect 17218 13172 17224 13184
rect 16899 13144 17224 13172
rect 16899 13141 16911 13144
rect 16853 13135 16911 13141
rect 17218 13132 17224 13144
rect 17276 13132 17282 13184
rect 17512 13181 17540 13212
rect 19886 13200 19892 13252
rect 19944 13200 19950 13252
rect 21358 13240 21364 13252
rect 21008 13212 21364 13240
rect 17497 13175 17555 13181
rect 17497 13141 17509 13175
rect 17543 13172 17555 13175
rect 18141 13175 18199 13181
rect 18141 13172 18153 13175
rect 17543 13144 18153 13172
rect 17543 13141 17555 13144
rect 17497 13135 17555 13141
rect 18141 13141 18153 13144
rect 18187 13141 18199 13175
rect 18141 13135 18199 13141
rect 19429 13175 19487 13181
rect 19429 13141 19441 13175
rect 19475 13172 19487 13175
rect 21008 13172 21036 13212
rect 21358 13200 21364 13212
rect 21416 13200 21422 13252
rect 19475 13144 21036 13172
rect 19475 13141 19487 13144
rect 19429 13135 19487 13141
rect 21174 13132 21180 13184
rect 21232 13172 21238 13184
rect 21560 13181 21588 13484
rect 22278 13472 22284 13484
rect 22336 13472 22342 13524
rect 21726 13268 21732 13320
rect 21784 13308 21790 13320
rect 22649 13311 22707 13317
rect 22649 13308 22661 13311
rect 21784 13280 22661 13308
rect 21784 13268 21790 13280
rect 22649 13277 22661 13280
rect 22695 13277 22707 13311
rect 22649 13271 22707 13277
rect 23845 13243 23903 13249
rect 23845 13209 23857 13243
rect 23891 13240 23903 13243
rect 25498 13240 25504 13252
rect 23891 13212 25504 13240
rect 23891 13209 23903 13212
rect 23845 13203 23903 13209
rect 25498 13200 25504 13212
rect 25556 13200 25562 13252
rect 21545 13175 21603 13181
rect 21545 13172 21557 13175
rect 21232 13144 21557 13172
rect 21232 13132 21238 13144
rect 21545 13141 21557 13144
rect 21591 13141 21603 13175
rect 21545 13135 21603 13141
rect 22002 13132 22008 13184
rect 22060 13132 22066 13184
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 8665 12971 8723 12977
rect 8665 12968 8677 12971
rect 7800 12940 8677 12968
rect 7800 12928 7806 12940
rect 8665 12937 8677 12940
rect 8711 12937 8723 12971
rect 8665 12931 8723 12937
rect 11149 12971 11207 12977
rect 11149 12937 11161 12971
rect 11195 12968 11207 12971
rect 11790 12968 11796 12980
rect 11195 12940 11796 12968
rect 11195 12937 11207 12940
rect 11149 12931 11207 12937
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 15286 12968 15292 12980
rect 13280 12940 15292 12968
rect 6638 12860 6644 12912
rect 6696 12900 6702 12912
rect 8386 12900 8392 12912
rect 6696 12872 8392 12900
rect 6696 12860 6702 12872
rect 8386 12860 8392 12872
rect 8444 12860 8450 12912
rect 9674 12900 9680 12912
rect 9416 12872 9680 12900
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 9416 12841 9444 12872
rect 9674 12860 9680 12872
rect 9732 12900 9738 12912
rect 9950 12900 9956 12912
rect 9732 12872 9956 12900
rect 9732 12860 9738 12872
rect 9950 12860 9956 12872
rect 10008 12860 10014 12912
rect 11514 12900 11520 12912
rect 10902 12872 11520 12900
rect 11514 12860 11520 12872
rect 11572 12900 11578 12912
rect 12802 12900 12808 12912
rect 11572 12872 12808 12900
rect 11572 12860 11578 12872
rect 12802 12860 12808 12872
rect 12860 12900 12866 12912
rect 13280 12909 13308 12940
rect 15286 12928 15292 12940
rect 15344 12968 15350 12980
rect 15746 12968 15752 12980
rect 15344 12940 15752 12968
rect 15344 12928 15350 12940
rect 15746 12928 15752 12940
rect 15804 12968 15810 12980
rect 15804 12940 15976 12968
rect 15804 12928 15810 12940
rect 13265 12903 13323 12909
rect 13265 12900 13277 12903
rect 12860 12872 13277 12900
rect 12860 12860 12866 12872
rect 13265 12869 13277 12872
rect 13311 12869 13323 12903
rect 13265 12863 13323 12869
rect 13725 12903 13783 12909
rect 13725 12869 13737 12903
rect 13771 12900 13783 12903
rect 13906 12900 13912 12912
rect 13771 12872 13912 12900
rect 13771 12869 13783 12872
rect 13725 12863 13783 12869
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 14366 12860 14372 12912
rect 14424 12900 14430 12912
rect 14461 12903 14519 12909
rect 14461 12900 14473 12903
rect 14424 12872 14473 12900
rect 14424 12860 14430 12872
rect 14461 12869 14473 12872
rect 14507 12900 14519 12903
rect 14921 12903 14979 12909
rect 14921 12900 14933 12903
rect 14507 12872 14933 12900
rect 14507 12869 14519 12872
rect 14461 12863 14519 12869
rect 14921 12869 14933 12872
rect 14967 12869 14979 12903
rect 14921 12863 14979 12869
rect 15194 12860 15200 12912
rect 15252 12900 15258 12912
rect 15381 12903 15439 12909
rect 15381 12900 15393 12903
rect 15252 12872 15393 12900
rect 15252 12860 15258 12872
rect 15381 12869 15393 12872
rect 15427 12900 15439 12903
rect 15841 12903 15899 12909
rect 15841 12900 15853 12903
rect 15427 12872 15853 12900
rect 15427 12869 15439 12872
rect 15381 12863 15439 12869
rect 15841 12869 15853 12872
rect 15887 12869 15899 12903
rect 15948 12900 15976 12940
rect 16114 12928 16120 12980
rect 16172 12928 16178 12980
rect 17218 12928 17224 12980
rect 17276 12928 17282 12980
rect 17310 12928 17316 12980
rect 17368 12928 17374 12980
rect 18322 12928 18328 12980
rect 18380 12968 18386 12980
rect 18969 12971 19027 12977
rect 18969 12968 18981 12971
rect 18380 12940 18981 12968
rect 18380 12928 18386 12940
rect 18524 12909 18552 12940
rect 18969 12937 18981 12940
rect 19015 12937 19027 12971
rect 20898 12968 20904 12980
rect 18969 12931 19027 12937
rect 19720 12940 20904 12968
rect 16393 12903 16451 12909
rect 16393 12900 16405 12903
rect 15948 12872 16405 12900
rect 15841 12863 15899 12869
rect 16393 12869 16405 12872
rect 16439 12869 16451 12903
rect 16393 12863 16451 12869
rect 18509 12903 18567 12909
rect 18509 12869 18521 12903
rect 18555 12900 18567 12903
rect 18555 12872 18589 12900
rect 18555 12869 18567 12872
rect 18509 12863 18567 12869
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 6604 12804 8585 12832
rect 6604 12792 6610 12804
rect 8573 12801 8585 12804
rect 8619 12801 8631 12835
rect 8573 12795 8631 12801
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 15930 12792 15936 12844
rect 15988 12832 15994 12844
rect 15988 12804 17448 12832
rect 15988 12792 15994 12804
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 9677 12767 9735 12773
rect 9677 12764 9689 12767
rect 8812 12736 9689 12764
rect 8812 12724 8818 12736
rect 9677 12733 9689 12736
rect 9723 12733 9735 12767
rect 14826 12764 14832 12776
rect 9677 12727 9735 12733
rect 10704 12736 14832 12764
rect 8205 12631 8263 12637
rect 8205 12597 8217 12631
rect 8251 12628 8263 12631
rect 10704 12628 10732 12736
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 17420 12773 17448 12804
rect 17405 12767 17463 12773
rect 17405 12733 17417 12767
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 18322 12724 18328 12776
rect 18380 12764 18386 12776
rect 19720 12773 19748 12940
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 20990 12928 20996 12980
rect 21048 12968 21054 12980
rect 21048 12940 21312 12968
rect 21048 12928 21054 12940
rect 21284 12832 21312 12940
rect 21450 12860 21456 12912
rect 21508 12900 21514 12912
rect 21508 12872 23980 12900
rect 21508 12860 21514 12872
rect 22281 12835 22339 12841
rect 19705 12767 19763 12773
rect 19705 12764 19717 12767
rect 18380 12736 19717 12764
rect 18380 12724 18386 12736
rect 19705 12733 19717 12736
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12764 20039 12767
rect 21100 12764 21128 12818
rect 21284 12804 21496 12832
rect 21174 12764 21180 12776
rect 20027 12736 21036 12764
rect 21100 12736 21180 12764
rect 20027 12733 20039 12736
rect 19981 12727 20039 12733
rect 13354 12656 13360 12708
rect 13412 12696 13418 12708
rect 13722 12696 13728 12708
rect 13412 12668 13728 12696
rect 13412 12656 13418 12668
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 13909 12699 13967 12705
rect 13909 12665 13921 12699
rect 13955 12696 13967 12699
rect 14274 12696 14280 12708
rect 13955 12668 14280 12696
rect 13955 12665 13967 12668
rect 13909 12659 13967 12665
rect 14274 12656 14280 12668
rect 14332 12656 14338 12708
rect 14642 12656 14648 12708
rect 14700 12656 14706 12708
rect 15930 12656 15936 12708
rect 15988 12696 15994 12708
rect 16114 12696 16120 12708
rect 15988 12668 16120 12696
rect 15988 12656 15994 12668
rect 16114 12656 16120 12668
rect 16172 12656 16178 12708
rect 16853 12699 16911 12705
rect 16853 12665 16865 12699
rect 16899 12696 16911 12699
rect 21008 12696 21036 12736
rect 21174 12724 21180 12736
rect 21232 12724 21238 12776
rect 21468 12773 21496 12804
rect 22281 12801 22293 12835
rect 22327 12832 22339 12835
rect 22462 12832 22468 12844
rect 22327 12804 22468 12832
rect 22327 12801 22339 12804
rect 22281 12795 22339 12801
rect 22462 12792 22468 12804
rect 22520 12792 22526 12844
rect 23290 12792 23296 12844
rect 23348 12792 23354 12844
rect 23952 12841 23980 12872
rect 23937 12835 23995 12841
rect 23937 12801 23949 12835
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 21453 12767 21511 12773
rect 21453 12733 21465 12767
rect 21499 12733 21511 12767
rect 21453 12727 21511 12733
rect 24762 12724 24768 12776
rect 24820 12724 24826 12776
rect 21818 12696 21824 12708
rect 16899 12668 19840 12696
rect 21008 12668 21824 12696
rect 16899 12665 16911 12668
rect 16853 12659 16911 12665
rect 8251 12600 10732 12628
rect 8251 12597 8263 12600
rect 8205 12591 8263 12597
rect 15470 12588 15476 12640
rect 15528 12588 15534 12640
rect 18598 12588 18604 12640
rect 18656 12588 18662 12640
rect 19812 12628 19840 12668
rect 21818 12656 21824 12668
rect 21876 12656 21882 12708
rect 20530 12628 20536 12640
rect 19812 12600 20536 12628
rect 20530 12588 20536 12600
rect 20588 12588 20594 12640
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 10870 12384 10876 12436
rect 10928 12424 10934 12436
rect 13817 12427 13875 12433
rect 13817 12424 13829 12427
rect 10928 12396 13829 12424
rect 10928 12384 10934 12396
rect 13817 12393 13829 12396
rect 13863 12393 13875 12427
rect 13817 12387 13875 12393
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 10962 12288 10968 12300
rect 9732 12260 10968 12288
rect 9732 12248 9738 12260
rect 10962 12248 10968 12260
rect 11020 12288 11026 12300
rect 11517 12291 11575 12297
rect 11517 12288 11529 12291
rect 11020 12260 11529 12288
rect 11020 12248 11026 12260
rect 11517 12257 11529 12260
rect 11563 12257 11575 12291
rect 11517 12251 11575 12257
rect 11790 12248 11796 12300
rect 11848 12248 11854 12300
rect 13832 12288 13860 12387
rect 13906 12384 13912 12436
rect 13964 12424 13970 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 13964 12396 14105 12424
rect 13964 12384 13970 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 14093 12387 14151 12393
rect 14458 12384 14464 12436
rect 14516 12384 14522 12436
rect 15654 12384 15660 12436
rect 15712 12384 15718 12436
rect 16022 12384 16028 12436
rect 16080 12424 16086 12436
rect 16080 12396 16252 12424
rect 16080 12384 16086 12396
rect 15930 12316 15936 12368
rect 15988 12356 15994 12368
rect 15988 12328 16160 12356
rect 15988 12316 15994 12328
rect 15013 12291 15071 12297
rect 15013 12288 15025 12291
rect 13832 12260 15025 12288
rect 15013 12257 15025 12260
rect 15059 12288 15071 12291
rect 15286 12288 15292 12300
rect 15059 12260 15292 12288
rect 15059 12257 15071 12260
rect 15013 12251 15071 12257
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 16132 12297 16160 12328
rect 16224 12297 16252 12396
rect 17494 12384 17500 12436
rect 17552 12424 17558 12436
rect 18877 12427 18935 12433
rect 18877 12424 18889 12427
rect 17552 12396 18889 12424
rect 17552 12384 17558 12396
rect 18877 12393 18889 12396
rect 18923 12393 18935 12427
rect 18877 12387 18935 12393
rect 22649 12359 22707 12365
rect 22649 12325 22661 12359
rect 22695 12356 22707 12359
rect 24854 12356 24860 12368
rect 22695 12328 24860 12356
rect 22695 12325 22707 12328
rect 22649 12319 22707 12325
rect 24854 12316 24860 12328
rect 24912 12316 24918 12368
rect 16117 12291 16175 12297
rect 16117 12257 16129 12291
rect 16163 12257 16175 12291
rect 16117 12251 16175 12257
rect 16209 12291 16267 12297
rect 16209 12257 16221 12291
rect 16255 12257 16267 12291
rect 16209 12251 16267 12257
rect 17126 12248 17132 12300
rect 17184 12248 17190 12300
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12288 17463 12291
rect 19978 12288 19984 12300
rect 17451 12260 19984 12288
rect 17451 12257 17463 12260
rect 17405 12251 17463 12257
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 21542 12248 21548 12300
rect 21600 12248 21606 12300
rect 21729 12291 21787 12297
rect 21729 12257 21741 12291
rect 21775 12288 21787 12291
rect 21818 12288 21824 12300
rect 21775 12260 21824 12288
rect 21775 12257 21787 12260
rect 21729 12251 21787 12257
rect 21818 12248 21824 12260
rect 21876 12248 21882 12300
rect 22186 12248 22192 12300
rect 22244 12288 22250 12300
rect 22244 12260 23520 12288
rect 22244 12248 22250 12260
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12220 14887 12223
rect 16942 12220 16948 12232
rect 14875 12192 16948 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 18874 12180 18880 12232
rect 18932 12220 18938 12232
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 18932 12192 20637 12220
rect 18932 12180 18938 12192
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 21453 12223 21511 12229
rect 21453 12189 21465 12223
rect 21499 12220 21511 12223
rect 22002 12220 22008 12232
rect 21499 12192 22008 12220
rect 21499 12189 21511 12192
rect 21453 12183 21511 12189
rect 22002 12180 22008 12192
rect 22060 12180 22066 12232
rect 23492 12229 23520 12260
rect 22833 12223 22891 12229
rect 22833 12189 22845 12223
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 23477 12223 23535 12229
rect 23477 12189 23489 12223
rect 23523 12189 23535 12223
rect 23477 12183 23535 12189
rect 12802 12112 12808 12164
rect 12860 12112 12866 12164
rect 16025 12155 16083 12161
rect 16025 12121 16037 12155
rect 16071 12152 16083 12155
rect 16482 12152 16488 12164
rect 16071 12124 16488 12152
rect 16071 12121 16083 12124
rect 16025 12115 16083 12121
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 17862 12152 17868 12164
rect 17788 12124 17868 12152
rect 13262 12044 13268 12096
rect 13320 12044 13326 12096
rect 13722 12044 13728 12096
rect 13780 12084 13786 12096
rect 14921 12087 14979 12093
rect 14921 12084 14933 12087
rect 13780 12056 14933 12084
rect 13780 12044 13786 12056
rect 14921 12053 14933 12056
rect 14967 12084 14979 12087
rect 17402 12084 17408 12096
rect 14967 12056 17408 12084
rect 14967 12053 14979 12056
rect 14921 12047 14979 12053
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 17788 12084 17816 12124
rect 17862 12112 17868 12124
rect 17920 12112 17926 12164
rect 18708 12124 19380 12152
rect 18708 12084 18736 12124
rect 19352 12093 19380 12124
rect 20162 12112 20168 12164
rect 20220 12152 20226 12164
rect 22848 12152 22876 12183
rect 20220 12124 22876 12152
rect 20220 12112 20226 12124
rect 17788 12056 18736 12084
rect 19337 12087 19395 12093
rect 19337 12053 19349 12087
rect 19383 12084 19395 12087
rect 19794 12084 19800 12096
rect 19383 12056 19800 12084
rect 19383 12053 19395 12056
rect 19337 12047 19395 12053
rect 19794 12044 19800 12056
rect 19852 12044 19858 12096
rect 20441 12087 20499 12093
rect 20441 12053 20453 12087
rect 20487 12084 20499 12087
rect 20990 12084 20996 12096
rect 20487 12056 20996 12084
rect 20487 12053 20499 12056
rect 20441 12047 20499 12053
rect 20990 12044 20996 12056
rect 21048 12044 21054 12096
rect 21082 12044 21088 12096
rect 21140 12044 21146 12096
rect 23293 12087 23351 12093
rect 23293 12053 23305 12087
rect 23339 12084 23351 12087
rect 25038 12084 25044 12096
rect 23339 12056 25044 12084
rect 23339 12053 23351 12056
rect 23293 12047 23351 12053
rect 25038 12044 25044 12056
rect 25096 12044 25102 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 13262 11880 13268 11892
rect 13096 11852 13268 11880
rect 13096 11821 13124 11852
rect 13262 11840 13268 11852
rect 13320 11880 13326 11892
rect 13320 11852 14872 11880
rect 13320 11840 13326 11852
rect 13081 11815 13139 11821
rect 13081 11781 13093 11815
rect 13127 11781 13139 11815
rect 13081 11775 13139 11781
rect 13170 11772 13176 11824
rect 13228 11812 13234 11824
rect 14844 11812 14872 11852
rect 15102 11840 15108 11892
rect 15160 11880 15166 11892
rect 15473 11883 15531 11889
rect 15473 11880 15485 11883
rect 15160 11852 15485 11880
rect 15160 11840 15166 11852
rect 15473 11849 15485 11852
rect 15519 11849 15531 11883
rect 15473 11843 15531 11849
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 16025 11883 16083 11889
rect 16025 11880 16037 11883
rect 15804 11852 16037 11880
rect 15804 11840 15810 11852
rect 16025 11849 16037 11852
rect 16071 11880 16083 11883
rect 17862 11880 17868 11892
rect 16071 11852 17868 11880
rect 16071 11849 16083 11852
rect 16025 11843 16083 11849
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 18322 11880 18328 11892
rect 18248 11852 18328 11880
rect 13228 11784 13570 11812
rect 14844 11784 15608 11812
rect 13228 11772 13234 11784
rect 10962 11704 10968 11756
rect 11020 11744 11026 11756
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 11020 11716 12817 11744
rect 11020 11704 11026 11716
rect 12805 11713 12817 11716
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 15102 11704 15108 11756
rect 15160 11744 15166 11756
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 15160 11716 15393 11744
rect 15160 11704 15166 11716
rect 15381 11713 15393 11716
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15580 11685 15608 11784
rect 16758 11772 16764 11824
rect 16816 11812 16822 11824
rect 16945 11815 17003 11821
rect 16945 11812 16957 11815
rect 16816 11784 16957 11812
rect 16816 11772 16822 11784
rect 16945 11781 16957 11784
rect 16991 11812 17003 11815
rect 17405 11815 17463 11821
rect 17405 11812 17417 11815
rect 16991 11784 17417 11812
rect 16991 11781 17003 11784
rect 16945 11775 17003 11781
rect 17405 11781 17417 11784
rect 17451 11781 17463 11815
rect 17405 11775 17463 11781
rect 18248 11753 18276 11852
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 19978 11840 19984 11892
rect 20036 11840 20042 11892
rect 20349 11883 20407 11889
rect 20349 11849 20361 11883
rect 20395 11880 20407 11883
rect 21174 11880 21180 11892
rect 20395 11852 21180 11880
rect 20395 11849 20407 11852
rect 20349 11843 20407 11849
rect 18506 11772 18512 11824
rect 18564 11772 18570 11824
rect 19794 11812 19800 11824
rect 19734 11784 19800 11812
rect 19794 11772 19800 11784
rect 19852 11812 19858 11824
rect 20364 11812 20392 11843
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 19852 11784 20392 11812
rect 19852 11772 19858 11784
rect 20806 11772 20812 11824
rect 20864 11812 20870 11824
rect 20901 11815 20959 11821
rect 20901 11812 20913 11815
rect 20864 11784 20913 11812
rect 20864 11772 20870 11784
rect 20901 11781 20913 11784
rect 20947 11812 20959 11815
rect 21361 11815 21419 11821
rect 21361 11812 21373 11815
rect 20947 11784 21373 11812
rect 20947 11781 20959 11784
rect 20901 11775 20959 11781
rect 21361 11781 21373 11784
rect 21407 11781 21419 11815
rect 21361 11775 21419 11781
rect 18233 11747 18291 11753
rect 18233 11713 18245 11747
rect 18279 11713 18291 11747
rect 18233 11707 18291 11713
rect 22830 11704 22836 11756
rect 22888 11744 22894 11756
rect 23293 11747 23351 11753
rect 23293 11744 23305 11747
rect 22888 11716 23305 11744
rect 22888 11704 22894 11716
rect 23293 11713 23305 11716
rect 23339 11713 23351 11747
rect 23293 11707 23351 11713
rect 15565 11679 15623 11685
rect 15565 11645 15577 11679
rect 15611 11645 15623 11679
rect 15565 11639 15623 11645
rect 16482 11636 16488 11688
rect 16540 11676 16546 11688
rect 19886 11676 19892 11688
rect 16540 11648 19892 11676
rect 16540 11636 16546 11648
rect 19886 11636 19892 11648
rect 19944 11636 19950 11688
rect 24026 11636 24032 11688
rect 24084 11636 24090 11688
rect 14550 11568 14556 11620
rect 14608 11568 14614 11620
rect 15013 11611 15071 11617
rect 15013 11577 15025 11611
rect 15059 11608 15071 11611
rect 21085 11611 21143 11617
rect 15059 11580 18368 11608
rect 15059 11577 15071 11580
rect 15013 11571 15071 11577
rect 18340 11552 18368 11580
rect 21085 11577 21097 11611
rect 21131 11608 21143 11611
rect 22002 11608 22008 11620
rect 21131 11580 22008 11608
rect 21131 11577 21143 11580
rect 21085 11571 21143 11577
rect 22002 11568 22008 11580
rect 22060 11568 22066 11620
rect 17034 11500 17040 11552
rect 17092 11500 17098 11552
rect 18322 11500 18328 11552
rect 18380 11500 18386 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 13998 11296 14004 11348
rect 14056 11336 14062 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 14056 11308 15485 11336
rect 14056 11296 14062 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 15473 11299 15531 11305
rect 14737 11203 14795 11209
rect 14737 11169 14749 11203
rect 14783 11200 14795 11203
rect 15102 11200 15108 11212
rect 14783 11172 15108 11200
rect 14783 11169 14795 11172
rect 14737 11163 14795 11169
rect 15102 11160 15108 11172
rect 15160 11160 15166 11212
rect 15286 11160 15292 11212
rect 15344 11200 15350 11212
rect 16025 11203 16083 11209
rect 16025 11200 16037 11203
rect 15344 11172 16037 11200
rect 15344 11160 15350 11172
rect 16025 11169 16037 11172
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11132 15899 11135
rect 20622 11132 20628 11144
rect 15887 11104 20628 11132
rect 15887 11101 15899 11104
rect 15841 11095 15899 11101
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 15194 11024 15200 11076
rect 15252 11064 15258 11076
rect 15933 11067 15991 11073
rect 15933 11064 15945 11067
rect 15252 11036 15945 11064
rect 15252 11024 15258 11036
rect 15933 11033 15945 11036
rect 15979 11064 15991 11067
rect 16298 11064 16304 11076
rect 15979 11036 16304 11064
rect 15979 11033 15991 11036
rect 15933 11027 15991 11033
rect 16298 11024 16304 11036
rect 16356 11024 16362 11076
rect 20806 11024 20812 11076
rect 20864 11024 20870 11076
rect 20993 11067 21051 11073
rect 20993 11033 21005 11067
rect 21039 11064 21051 11067
rect 23934 11064 23940 11076
rect 21039 11036 23940 11064
rect 21039 11033 21051 11036
rect 20993 11027 21051 11033
rect 23934 11024 23940 11036
rect 23992 11024 23998 11076
rect 19610 10956 19616 11008
rect 19668 10956 19674 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 15286 10752 15292 10804
rect 15344 10752 15350 10804
rect 19521 10795 19579 10801
rect 19521 10761 19533 10795
rect 19567 10792 19579 10795
rect 19610 10792 19616 10804
rect 19567 10764 19616 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 19610 10752 19616 10764
rect 19668 10752 19674 10804
rect 20349 10795 20407 10801
rect 20349 10761 20361 10795
rect 20395 10792 20407 10795
rect 20395 10764 22094 10792
rect 20395 10761 20407 10764
rect 20349 10755 20407 10761
rect 10226 10684 10232 10736
rect 10284 10724 10290 10736
rect 12069 10727 12127 10733
rect 12069 10724 12081 10727
rect 10284 10696 12081 10724
rect 10284 10684 10290 10696
rect 12069 10693 12081 10696
rect 12115 10724 12127 10727
rect 12529 10727 12587 10733
rect 12529 10724 12541 10727
rect 12115 10696 12541 10724
rect 12115 10693 12127 10696
rect 12069 10687 12127 10693
rect 12529 10693 12541 10696
rect 12575 10693 12587 10727
rect 22066 10724 22094 10764
rect 22066 10696 23428 10724
rect 12529 10687 12587 10693
rect 14826 10616 14832 10668
rect 14884 10616 14890 10668
rect 18322 10616 18328 10668
rect 18380 10656 18386 10668
rect 18417 10659 18475 10665
rect 18417 10656 18429 10659
rect 18380 10628 18429 10656
rect 18380 10616 18386 10628
rect 18417 10625 18429 10628
rect 18463 10625 18475 10659
rect 18417 10619 18475 10625
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 19613 10659 19671 10665
rect 19613 10656 19625 10659
rect 19392 10628 19625 10656
rect 19392 10616 19398 10628
rect 19613 10625 19625 10628
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 20530 10616 20536 10668
rect 20588 10616 20594 10668
rect 23400 10665 23428 10696
rect 23385 10659 23443 10665
rect 23385 10625 23397 10659
rect 23431 10625 23443 10659
rect 23385 10619 23443 10625
rect 23658 10616 23664 10668
rect 23716 10656 23722 10668
rect 23937 10659 23995 10665
rect 23937 10656 23949 10659
rect 23716 10628 23949 10656
rect 23716 10616 23722 10628
rect 23937 10625 23949 10628
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 19797 10591 19855 10597
rect 19797 10557 19809 10591
rect 19843 10588 19855 10591
rect 19978 10588 19984 10600
rect 19843 10560 19984 10588
rect 19843 10557 19855 10560
rect 19797 10551 19855 10557
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 12253 10523 12311 10529
rect 12253 10489 12265 10523
rect 12299 10520 12311 10523
rect 12434 10520 12440 10532
rect 12299 10492 12440 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 12434 10480 12440 10492
rect 12492 10480 12498 10532
rect 14645 10523 14703 10529
rect 14645 10489 14657 10523
rect 14691 10520 14703 10523
rect 20806 10520 20812 10532
rect 14691 10492 20812 10520
rect 14691 10489 14703 10492
rect 14645 10483 14703 10489
rect 20806 10480 20812 10492
rect 20864 10480 20870 10532
rect 15194 10412 15200 10464
rect 15252 10412 15258 10464
rect 18230 10412 18236 10464
rect 18288 10412 18294 10464
rect 19153 10455 19211 10461
rect 19153 10421 19165 10455
rect 19199 10452 19211 10455
rect 20622 10452 20628 10464
rect 19199 10424 20628 10452
rect 19199 10421 19211 10424
rect 19153 10415 19211 10421
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 23201 10455 23259 10461
rect 23201 10421 23213 10455
rect 23247 10452 23259 10455
rect 23290 10452 23296 10464
rect 23247 10424 23296 10452
rect 23247 10421 23259 10424
rect 23201 10415 23259 10421
rect 23290 10412 23296 10424
rect 23348 10412 23354 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 20990 10140 20996 10192
rect 21048 10180 21054 10192
rect 21048 10152 22784 10180
rect 21048 10140 21054 10152
rect 18230 10072 18236 10124
rect 18288 10112 18294 10124
rect 18288 10084 22232 10112
rect 18288 10072 18294 10084
rect 13446 10004 13452 10056
rect 13504 10044 13510 10056
rect 14645 10047 14703 10053
rect 14645 10044 14657 10047
rect 13504 10016 14657 10044
rect 13504 10004 13510 10016
rect 14645 10013 14657 10016
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10044 16819 10047
rect 18690 10044 18696 10056
rect 16807 10016 18696 10044
rect 16807 10013 16819 10016
rect 16761 10007 16819 10013
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 21358 10004 21364 10056
rect 21416 10044 21422 10056
rect 22204 10053 22232 10084
rect 21453 10047 21511 10053
rect 21453 10044 21465 10047
rect 21416 10016 21465 10044
rect 21416 10004 21422 10016
rect 21453 10013 21465 10016
rect 21499 10013 21511 10047
rect 21453 10007 21511 10013
rect 22189 10047 22247 10053
rect 22189 10013 22201 10047
rect 22235 10013 22247 10047
rect 22189 10007 22247 10013
rect 22649 10047 22707 10053
rect 22649 10013 22661 10047
rect 22695 10013 22707 10047
rect 22649 10007 22707 10013
rect 14829 9979 14887 9985
rect 14829 9945 14841 9979
rect 14875 9976 14887 9979
rect 19426 9976 19432 9988
rect 14875 9948 19432 9976
rect 14875 9945 14887 9948
rect 14829 9939 14887 9945
rect 19426 9936 19432 9948
rect 19484 9936 19490 9988
rect 22664 9976 22692 10007
rect 22020 9948 22692 9976
rect 22756 9976 22784 10152
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10044 23903 10047
rect 24946 10044 24952 10056
rect 23891 10016 24952 10044
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 24673 9979 24731 9985
rect 24673 9976 24685 9979
rect 22756 9948 24685 9976
rect 16850 9868 16856 9920
rect 16908 9868 16914 9920
rect 21269 9911 21327 9917
rect 21269 9877 21281 9911
rect 21315 9908 21327 9911
rect 21726 9908 21732 9920
rect 21315 9880 21732 9908
rect 21315 9877 21327 9880
rect 21269 9871 21327 9877
rect 21726 9868 21732 9880
rect 21784 9868 21790 9920
rect 22020 9917 22048 9948
rect 24673 9945 24685 9948
rect 24719 9945 24731 9979
rect 24673 9939 24731 9945
rect 22005 9911 22063 9917
rect 22005 9877 22017 9911
rect 22051 9877 22063 9911
rect 22005 9871 22063 9877
rect 24026 9868 24032 9920
rect 24084 9908 24090 9920
rect 24765 9911 24823 9917
rect 24765 9908 24777 9911
rect 24084 9880 24777 9908
rect 24084 9868 24090 9880
rect 24765 9877 24777 9880
rect 24811 9877 24823 9911
rect 24765 9871 24823 9877
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 16206 9596 16212 9648
rect 16264 9636 16270 9648
rect 16945 9639 17003 9645
rect 16945 9636 16957 9639
rect 16264 9608 16957 9636
rect 16264 9596 16270 9608
rect 16945 9605 16957 9608
rect 16991 9605 17003 9639
rect 16945 9599 17003 9605
rect 21910 9596 21916 9648
rect 21968 9636 21974 9648
rect 21968 9608 23980 9636
rect 21968 9596 21974 9608
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 5859 9540 6929 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 19058 9528 19064 9580
rect 19116 9568 19122 9580
rect 19245 9571 19303 9577
rect 19245 9568 19257 9571
rect 19116 9540 19257 9568
rect 19116 9528 19122 9540
rect 19245 9537 19257 9540
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 21082 9528 21088 9580
rect 21140 9568 21146 9580
rect 23952 9577 23980 9608
rect 22925 9571 22983 9577
rect 22925 9568 22937 9571
rect 21140 9540 22937 9568
rect 21140 9528 21146 9540
rect 22925 9537 22937 9540
rect 22971 9537 22983 9571
rect 22925 9531 22983 9537
rect 23937 9571 23995 9577
rect 23937 9537 23949 9571
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 4430 9460 4436 9512
rect 4488 9500 4494 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 4488 9472 7021 9500
rect 4488 9460 4494 9472
rect 7009 9469 7021 9472
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 7098 9460 7104 9512
rect 7156 9460 7162 9512
rect 23382 9460 23388 9512
rect 23440 9500 23446 9512
rect 24397 9503 24455 9509
rect 24397 9500 24409 9503
rect 23440 9472 24409 9500
rect 23440 9460 23446 9472
rect 24397 9469 24409 9472
rect 24443 9469 24455 9503
rect 24397 9463 24455 9469
rect 6546 9392 6552 9444
rect 6604 9392 6610 9444
rect 17129 9435 17187 9441
rect 17129 9401 17141 9435
rect 17175 9432 17187 9435
rect 17586 9432 17592 9444
rect 17175 9404 17592 9432
rect 17175 9401 17187 9404
rect 17129 9395 17187 9401
rect 17586 9392 17592 9404
rect 17644 9392 17650 9444
rect 17678 9324 17684 9376
rect 17736 9364 17742 9376
rect 19061 9367 19119 9373
rect 19061 9364 19073 9367
rect 17736 9336 19073 9364
rect 17736 9324 17742 9336
rect 19061 9333 19073 9336
rect 19107 9333 19119 9367
rect 19061 9327 19119 9333
rect 22738 9324 22744 9376
rect 22796 9324 22802 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 3602 9052 3608 9104
rect 3660 9092 3666 9104
rect 4890 9092 4896 9104
rect 3660 9064 4896 9092
rect 3660 9052 3666 9064
rect 4890 9052 4896 9064
rect 4948 9052 4954 9104
rect 22462 9052 22468 9104
rect 22520 9092 22526 9104
rect 24673 9095 24731 9101
rect 24673 9092 24685 9095
rect 22520 9064 24685 9092
rect 22520 9052 22526 9064
rect 24673 9061 24685 9064
rect 24719 9061 24731 9095
rect 24673 9055 24731 9061
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 21729 8959 21787 8965
rect 21729 8956 21741 8959
rect 20680 8928 21741 8956
rect 20680 8916 20686 8928
rect 21729 8925 21741 8928
rect 21775 8925 21787 8959
rect 21729 8919 21787 8925
rect 22646 8916 22652 8968
rect 22704 8956 22710 8968
rect 23937 8959 23995 8965
rect 23937 8956 23949 8959
rect 22704 8928 23949 8956
rect 22704 8916 22710 8928
rect 23937 8925 23949 8928
rect 23983 8925 23995 8959
rect 23937 8919 23995 8925
rect 24854 8916 24860 8968
rect 24912 8916 24918 8968
rect 21545 8823 21603 8829
rect 21545 8789 21557 8823
rect 21591 8820 21603 8823
rect 22554 8820 22560 8832
rect 21591 8792 22560 8820
rect 21591 8789 21603 8792
rect 21545 8783 21603 8789
rect 22554 8780 22560 8792
rect 22612 8780 22618 8832
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 23753 8823 23811 8829
rect 23753 8820 23765 8823
rect 23532 8792 23765 8820
rect 23532 8780 23538 8792
rect 23753 8789 23765 8792
rect 23799 8789 23811 8823
rect 23753 8783 23811 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 19150 8508 19156 8560
rect 19208 8548 19214 8560
rect 19613 8551 19671 8557
rect 19613 8548 19625 8551
rect 19208 8520 19625 8548
rect 19208 8508 19214 8520
rect 19613 8517 19625 8520
rect 19659 8517 19671 8551
rect 19613 8511 19671 8517
rect 20717 8551 20775 8557
rect 20717 8517 20729 8551
rect 20763 8548 20775 8551
rect 21266 8548 21272 8560
rect 20763 8520 21272 8548
rect 20763 8517 20775 8520
rect 20717 8511 20775 8517
rect 21266 8508 21272 8520
rect 21324 8508 21330 8560
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8480 22339 8483
rect 22646 8480 22652 8492
rect 22327 8452 22652 8480
rect 22327 8449 22339 8452
rect 22281 8443 22339 8449
rect 22646 8440 22652 8452
rect 22704 8440 22710 8492
rect 23934 8440 23940 8492
rect 23992 8440 23998 8492
rect 23290 8372 23296 8424
rect 23348 8372 23354 8424
rect 24670 8372 24676 8424
rect 24728 8372 24734 8424
rect 19337 8347 19395 8353
rect 19337 8313 19349 8347
rect 19383 8344 19395 8347
rect 20714 8344 20720 8356
rect 19383 8316 20720 8344
rect 19383 8313 19395 8316
rect 19337 8307 19395 8313
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 20901 8347 20959 8353
rect 20901 8313 20913 8347
rect 20947 8344 20959 8347
rect 21266 8344 21272 8356
rect 20947 8316 21272 8344
rect 20947 8313 20959 8316
rect 20901 8307 20959 8313
rect 21266 8304 21272 8316
rect 21324 8304 21330 8356
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 6457 8075 6515 8081
rect 6457 8041 6469 8075
rect 6503 8072 6515 8075
rect 6546 8072 6552 8084
rect 6503 8044 6552 8072
rect 6503 8041 6515 8044
rect 6457 8035 6515 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 6641 8075 6699 8081
rect 6641 8041 6653 8075
rect 6687 8072 6699 8075
rect 6822 8072 6828 8084
rect 6687 8044 6828 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 6656 7936 6684 8035
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 22830 8032 22836 8084
rect 22888 8072 22894 8084
rect 24581 8075 24639 8081
rect 24581 8072 24593 8075
rect 22888 8044 24593 8072
rect 22888 8032 22894 8044
rect 24581 8041 24593 8044
rect 24627 8041 24639 8075
rect 24581 8035 24639 8041
rect 4111 7908 6684 7936
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 6546 7868 6552 7880
rect 5474 7840 6552 7868
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 19886 7828 19892 7880
rect 19944 7868 19950 7880
rect 20441 7871 20499 7877
rect 20441 7868 20453 7871
rect 19944 7840 20453 7868
rect 19944 7828 19950 7840
rect 20441 7837 20453 7840
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 21269 7871 21327 7877
rect 21269 7868 21281 7871
rect 20588 7840 21281 7868
rect 20588 7828 20594 7840
rect 21269 7837 21281 7840
rect 21315 7837 21327 7871
rect 21269 7831 21327 7837
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7868 22891 7871
rect 23474 7868 23480 7880
rect 22879 7840 23480 7868
rect 22879 7837 22891 7840
rect 22833 7831 22891 7837
rect 23474 7828 23480 7840
rect 23532 7828 23538 7880
rect 24765 7871 24823 7877
rect 24765 7837 24777 7871
rect 24811 7868 24823 7871
rect 24854 7868 24860 7880
rect 24811 7840 24860 7868
rect 24811 7837 24823 7840
rect 24765 7831 24823 7837
rect 24854 7828 24860 7840
rect 24912 7828 24918 7880
rect 4338 7760 4344 7812
rect 4396 7760 4402 7812
rect 6089 7803 6147 7809
rect 6089 7769 6101 7803
rect 6135 7800 6147 7803
rect 9214 7800 9220 7812
rect 6135 7772 9220 7800
rect 6135 7769 6147 7772
rect 6089 7763 6147 7769
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 23845 7803 23903 7809
rect 23845 7769 23857 7803
rect 23891 7800 23903 7803
rect 24486 7800 24492 7812
rect 23891 7772 24492 7800
rect 23891 7769 23903 7772
rect 23845 7763 23903 7769
rect 24486 7760 24492 7772
rect 24544 7760 24550 7812
rect 20257 7735 20315 7741
rect 20257 7701 20269 7735
rect 20303 7732 20315 7735
rect 20806 7732 20812 7744
rect 20303 7704 20812 7732
rect 20303 7701 20315 7704
rect 20257 7695 20315 7701
rect 20806 7692 20812 7704
rect 20864 7692 20870 7744
rect 21082 7692 21088 7744
rect 21140 7692 21146 7744
rect 22462 7692 22468 7744
rect 22520 7732 22526 7744
rect 22830 7732 22836 7744
rect 22520 7704 22836 7732
rect 22520 7692 22526 7704
rect 22830 7692 22836 7704
rect 22888 7692 22894 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 16942 7420 16948 7472
rect 17000 7460 17006 7472
rect 18785 7463 18843 7469
rect 18785 7460 18797 7463
rect 17000 7432 18797 7460
rect 17000 7420 17006 7432
rect 18785 7429 18797 7432
rect 18831 7429 18843 7463
rect 18785 7423 18843 7429
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 20272 7324 20300 7355
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 20772 7364 22109 7392
rect 20772 7352 20778 7364
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 23382 7352 23388 7404
rect 23440 7392 23446 7404
rect 23937 7395 23995 7401
rect 23937 7392 23949 7395
rect 23440 7364 23949 7392
rect 23440 7352 23446 7364
rect 23937 7361 23949 7364
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 20898 7324 20904 7336
rect 20272 7296 20904 7324
rect 20898 7284 20904 7296
rect 20956 7284 20962 7336
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 21358 7324 21364 7336
rect 21315 7296 21364 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 21358 7284 21364 7296
rect 21416 7284 21422 7336
rect 22278 7284 22284 7336
rect 22336 7324 22342 7336
rect 22557 7327 22615 7333
rect 22557 7324 22569 7327
rect 22336 7296 22569 7324
rect 22336 7284 22342 7296
rect 22557 7293 22569 7296
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 18969 7259 19027 7265
rect 18969 7225 18981 7259
rect 19015 7256 19027 7259
rect 20622 7256 20628 7268
rect 19015 7228 20628 7256
rect 19015 7225 19027 7228
rect 18969 7219 19027 7225
rect 20622 7216 20628 7228
rect 20680 7216 20686 7268
rect 22554 7148 22560 7200
rect 22612 7188 22618 7200
rect 23382 7188 23388 7200
rect 22612 7160 23388 7188
rect 22612 7148 22618 7160
rect 23382 7148 23388 7160
rect 23440 7148 23446 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 15896 6752 19717 6780
rect 15896 6740 15902 6752
rect 19705 6749 19717 6752
rect 19751 6780 19763 6783
rect 19981 6783 20039 6789
rect 19981 6780 19993 6783
rect 19751 6752 19993 6780
rect 19751 6749 19763 6752
rect 19705 6743 19763 6749
rect 19981 6749 19993 6752
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 20806 6740 20812 6792
rect 20864 6740 20870 6792
rect 22830 6740 22836 6792
rect 22888 6740 22894 6792
rect 24857 6783 24915 6789
rect 24857 6749 24869 6783
rect 24903 6780 24915 6783
rect 24946 6780 24952 6792
rect 24903 6752 24952 6780
rect 24903 6749 24915 6752
rect 24857 6743 24915 6749
rect 24946 6740 24952 6752
rect 25004 6740 25010 6792
rect 21818 6672 21824 6724
rect 21876 6672 21882 6724
rect 23845 6715 23903 6721
rect 23845 6681 23857 6715
rect 23891 6712 23903 6715
rect 25038 6712 25044 6724
rect 23891 6684 25044 6712
rect 23891 6681 23903 6684
rect 23845 6675 23903 6681
rect 25038 6672 25044 6684
rect 25096 6672 25102 6724
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 19521 6647 19579 6653
rect 19521 6644 19533 6647
rect 18380 6616 19533 6644
rect 18380 6604 18386 6616
rect 19521 6613 19533 6616
rect 19567 6613 19579 6647
rect 19521 6607 19579 6613
rect 24670 6604 24676 6656
rect 24728 6604 24734 6656
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 1854 6400 1860 6452
rect 1912 6400 1918 6452
rect 3697 6443 3755 6449
rect 3697 6409 3709 6443
rect 3743 6440 3755 6443
rect 4338 6440 4344 6452
rect 3743 6412 4344 6440
rect 3743 6409 3755 6412
rect 3697 6403 3755 6409
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 17957 6443 18015 6449
rect 17957 6440 17969 6443
rect 11664 6412 17969 6440
rect 11664 6400 11670 6412
rect 17957 6409 17969 6412
rect 18003 6409 18015 6443
rect 17957 6403 18015 6409
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1688 6236 1716 6267
rect 2406 6264 2412 6316
rect 2464 6304 2470 6316
rect 2593 6307 2651 6313
rect 2593 6304 2605 6307
rect 2464 6276 2605 6304
rect 2464 6264 2470 6276
rect 2593 6273 2605 6276
rect 2639 6273 2651 6307
rect 2593 6267 2651 6273
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 3326 6304 3332 6316
rect 3099 6276 3332 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 17972 6304 18000 6403
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 17972 6276 18245 6304
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6304 20315 6307
rect 21082 6304 21088 6316
rect 20303 6276 21088 6304
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 22002 6264 22008 6316
rect 22060 6264 22066 6316
rect 22554 6264 22560 6316
rect 22612 6304 22618 6316
rect 23937 6307 23995 6313
rect 23937 6304 23949 6307
rect 22612 6276 23949 6304
rect 22612 6264 22618 6276
rect 23937 6273 23949 6276
rect 23983 6273 23995 6307
rect 23937 6267 23995 6273
rect 2774 6236 2780 6248
rect 1688 6208 2780 6236
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 19429 6239 19487 6245
rect 19429 6205 19441 6239
rect 19475 6236 19487 6239
rect 20714 6236 20720 6248
rect 19475 6208 20720 6236
rect 19475 6205 19487 6208
rect 19429 6199 19487 6205
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 21269 6239 21327 6245
rect 21269 6205 21281 6239
rect 21315 6236 21327 6239
rect 21450 6236 21456 6248
rect 21315 6208 21456 6236
rect 21315 6205 21327 6208
rect 21269 6199 21327 6205
rect 21450 6196 21456 6208
rect 21508 6196 21514 6248
rect 21910 6196 21916 6248
rect 21968 6236 21974 6248
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 21968 6208 22477 6236
rect 21968 6196 21974 6208
rect 22465 6205 22477 6208
rect 22511 6205 22523 6239
rect 22465 6199 22523 6205
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 2409 6103 2467 6109
rect 2409 6069 2421 6103
rect 2455 6100 2467 6103
rect 2498 6100 2504 6112
rect 2455 6072 2504 6100
rect 2455 6069 2467 6072
rect 2409 6063 2467 6069
rect 2498 6060 2504 6072
rect 2556 6060 2562 6112
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 3145 5899 3203 5905
rect 3145 5865 3157 5899
rect 3191 5896 3203 5899
rect 3326 5896 3332 5908
rect 3191 5868 3332 5896
rect 3191 5865 3203 5868
rect 3145 5859 3203 5865
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 9306 5896 9312 5908
rect 4212 5868 9312 5896
rect 4212 5856 4218 5868
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 20898 5856 20904 5908
rect 20956 5896 20962 5908
rect 24765 5899 24823 5905
rect 24765 5896 24777 5899
rect 20956 5868 24777 5896
rect 20956 5856 20962 5868
rect 24765 5865 24777 5868
rect 24811 5865 24823 5899
rect 24765 5859 24823 5865
rect 2041 5831 2099 5837
rect 2041 5797 2053 5831
rect 2087 5828 2099 5831
rect 4982 5828 4988 5840
rect 2087 5800 4988 5828
rect 2087 5797 2099 5800
rect 2041 5791 2099 5797
rect 4982 5788 4988 5800
rect 5040 5788 5046 5840
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 10778 5760 10784 5772
rect 5960 5732 10784 5760
rect 5960 5720 5966 5732
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 20993 5763 21051 5769
rect 20993 5760 21005 5763
rect 20496 5732 21005 5760
rect 20496 5720 20502 5732
rect 20993 5729 21005 5732
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 21542 5720 21548 5772
rect 21600 5760 21606 5772
rect 22833 5763 22891 5769
rect 22833 5760 22845 5763
rect 21600 5732 22845 5760
rect 21600 5720 21606 5732
rect 22833 5729 22845 5732
rect 22879 5729 22891 5763
rect 22833 5723 22891 5729
rect 2498 5652 2504 5704
rect 2556 5652 2562 5704
rect 3050 5652 3056 5704
rect 3108 5692 3114 5704
rect 8662 5692 8668 5704
rect 3108 5664 8668 5692
rect 3108 5652 3114 5664
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 17678 5652 17684 5704
rect 17736 5652 17742 5704
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20533 5695 20591 5701
rect 20533 5692 20545 5695
rect 20404 5664 20545 5692
rect 20404 5652 20410 5664
rect 20533 5661 20545 5664
rect 20579 5661 20591 5695
rect 20533 5655 20591 5661
rect 20622 5652 20628 5704
rect 20680 5692 20686 5704
rect 22373 5695 22431 5701
rect 22373 5692 22385 5695
rect 20680 5664 22385 5692
rect 20680 5652 20686 5664
rect 22373 5661 22385 5664
rect 22419 5661 22431 5695
rect 22373 5655 22431 5661
rect 1854 5584 1860 5636
rect 1912 5584 1918 5636
rect 2130 5584 2136 5636
rect 2188 5624 2194 5636
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 2188 5596 3801 5624
rect 2188 5584 2194 5596
rect 3789 5593 3801 5596
rect 3835 5593 3847 5627
rect 3789 5587 3847 5593
rect 9306 5584 9312 5636
rect 9364 5624 9370 5636
rect 18693 5627 18751 5633
rect 9364 5596 12434 5624
rect 9364 5584 9370 5596
rect 3602 5516 3608 5568
rect 3660 5516 3666 5568
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 3973 5559 4031 5565
rect 3973 5556 3985 5559
rect 3936 5528 3985 5556
rect 3936 5516 3942 5528
rect 3973 5525 3985 5528
rect 4019 5525 4031 5559
rect 3973 5519 4031 5525
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 6362 5556 6368 5568
rect 4856 5528 6368 5556
rect 4856 5516 4862 5528
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 8846 5516 8852 5568
rect 8904 5556 8910 5568
rect 10318 5556 10324 5568
rect 8904 5528 10324 5556
rect 8904 5516 8910 5528
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 12406 5556 12434 5596
rect 18693 5593 18705 5627
rect 18739 5624 18751 5627
rect 21174 5624 21180 5636
rect 18739 5596 21180 5624
rect 18739 5593 18751 5596
rect 18693 5587 18751 5593
rect 21174 5584 21180 5596
rect 21232 5584 21238 5636
rect 24673 5627 24731 5633
rect 24673 5593 24685 5627
rect 24719 5593 24731 5627
rect 24673 5587 24731 5593
rect 14090 5556 14096 5568
rect 12406 5528 14096 5556
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 21726 5516 21732 5568
rect 21784 5556 21790 5568
rect 24688 5556 24716 5587
rect 21784 5528 24716 5556
rect 21784 5516 21790 5528
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 3050 5312 3056 5364
rect 3108 5312 3114 5364
rect 3786 5312 3792 5364
rect 3844 5312 3850 5364
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 4430 5352 4436 5364
rect 4387 5324 4436 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 5166 5312 5172 5364
rect 5224 5312 5230 5364
rect 2409 5287 2467 5293
rect 2409 5253 2421 5287
rect 2455 5284 2467 5287
rect 2455 5256 4568 5284
rect 2455 5253 2467 5256
rect 2409 5247 2467 5253
rect 1670 5176 1676 5228
rect 1728 5216 1734 5228
rect 1765 5219 1823 5225
rect 1765 5216 1777 5219
rect 1728 5188 1777 5216
rect 1728 5176 1734 5188
rect 1765 5185 1777 5188
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 2866 5176 2872 5228
rect 2924 5176 2930 5228
rect 4540 5225 4568 5256
rect 19334 5244 19340 5296
rect 19392 5284 19398 5296
rect 20349 5287 20407 5293
rect 20349 5284 20361 5287
rect 19392 5256 20361 5284
rect 19392 5244 19398 5256
rect 20349 5253 20361 5256
rect 20395 5253 20407 5287
rect 20349 5247 20407 5253
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5994 5216 6000 5228
rect 5031 5188 6000 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 2314 5108 2320 5160
rect 2372 5148 2378 5160
rect 3620 5148 3648 5179
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 17770 5176 17776 5228
rect 17828 5176 17834 5228
rect 19518 5176 19524 5228
rect 19576 5176 19582 5228
rect 22186 5176 22192 5228
rect 22244 5176 22250 5228
rect 24026 5176 24032 5228
rect 24084 5176 24090 5228
rect 2372 5120 3648 5148
rect 18785 5151 18843 5157
rect 2372 5108 2378 5120
rect 18785 5117 18797 5151
rect 18831 5148 18843 5151
rect 20254 5148 20260 5160
rect 18831 5120 20260 5148
rect 18831 5117 18843 5120
rect 18785 5111 18843 5117
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 22462 5108 22468 5160
rect 22520 5108 22526 5160
rect 24578 5108 24584 5160
rect 24636 5108 24642 5160
rect 1489 5015 1547 5021
rect 1489 4981 1501 5015
rect 1535 5012 1547 5015
rect 1670 5012 1676 5024
rect 1535 4984 1676 5012
rect 1535 4981 1547 4984
rect 1489 4975 1547 4981
rect 1670 4972 1676 4984
rect 1728 4972 1734 5024
rect 5350 4972 5356 5024
rect 5408 5012 5414 5024
rect 6089 5015 6147 5021
rect 6089 5012 6101 5015
rect 5408 4984 6101 5012
rect 5408 4972 5414 4984
rect 6089 4981 6101 4984
rect 6135 4981 6147 5015
rect 6089 4975 6147 4981
rect 7374 4972 7380 5024
rect 7432 4972 7438 5024
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 4154 4768 4160 4820
rect 4212 4768 4218 4820
rect 5902 4768 5908 4820
rect 5960 4768 5966 4820
rect 6730 4768 6736 4820
rect 6788 4768 6794 4820
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7745 4811 7803 4817
rect 7745 4808 7757 4811
rect 7064 4780 7757 4808
rect 7064 4768 7070 4780
rect 7745 4777 7757 4780
rect 7791 4777 7803 4811
rect 7745 4771 7803 4777
rect 8478 4768 8484 4820
rect 8536 4768 8542 4820
rect 9769 4811 9827 4817
rect 9769 4777 9781 4811
rect 9815 4808 9827 4811
rect 12342 4808 12348 4820
rect 9815 4780 12348 4808
rect 9815 4777 9827 4780
rect 9769 4771 9827 4777
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 17770 4768 17776 4820
rect 17828 4808 17834 4820
rect 23845 4811 23903 4817
rect 23845 4808 23857 4811
rect 17828 4780 23857 4808
rect 17828 4768 17834 4780
rect 23845 4777 23857 4780
rect 23891 4777 23903 4811
rect 23845 4771 23903 4777
rect 5169 4743 5227 4749
rect 5169 4709 5181 4743
rect 5215 4740 5227 4743
rect 10042 4740 10048 4752
rect 5215 4712 10048 4740
rect 5215 4709 5227 4712
rect 5169 4703 5227 4709
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 11701 4743 11759 4749
rect 11701 4709 11713 4743
rect 11747 4740 11759 4743
rect 15194 4740 15200 4752
rect 11747 4712 15200 4740
rect 11747 4709 11759 4712
rect 11701 4703 11759 4709
rect 15194 4700 15200 4712
rect 15252 4700 15258 4752
rect 22646 4700 22652 4752
rect 22704 4740 22710 4752
rect 24857 4743 24915 4749
rect 24857 4740 24869 4743
rect 22704 4712 24869 4740
rect 22704 4700 22710 4712
rect 24857 4709 24869 4712
rect 24903 4709 24915 4743
rect 24857 4703 24915 4709
rect 3329 4675 3387 4681
rect 3329 4672 3341 4675
rect 1596 4644 3341 4672
rect 1596 4613 1624 4644
rect 3329 4641 3341 4644
rect 3375 4641 3387 4675
rect 4525 4675 4583 4681
rect 4525 4672 4537 4675
rect 3329 4635 3387 4641
rect 3436 4644 4537 4672
rect 3436 4616 3464 4644
rect 4525 4641 4537 4644
rect 4571 4641 4583 4675
rect 4525 4635 4583 4641
rect 19886 4632 19892 4684
rect 19944 4632 19950 4684
rect 21726 4632 21732 4684
rect 21784 4632 21790 4684
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4573 1639 4607
rect 1581 4567 1639 4573
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 3418 4604 3424 4616
rect 2731 4576 3424 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 4982 4564 4988 4616
rect 5040 4564 5046 4616
rect 5718 4564 5724 4616
rect 5776 4564 5782 4616
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4604 6607 4607
rect 7190 4604 7196 4616
rect 6595 4576 7196 4604
rect 6595 4573 6607 4576
rect 6549 4567 6607 4573
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 8294 4564 8300 4616
rect 8352 4564 8358 4616
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4604 9643 4607
rect 9858 4604 9864 4616
rect 9631 4576 9864 4604
rect 9631 4573 9643 4576
rect 9585 4567 9643 4573
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 11606 4564 11612 4616
rect 11664 4604 11670 4616
rect 11885 4607 11943 4613
rect 11885 4604 11897 4607
rect 11664 4576 11897 4604
rect 11664 4564 11670 4576
rect 11885 4573 11897 4576
rect 11931 4604 11943 4607
rect 12161 4607 12219 4613
rect 12161 4604 12173 4607
rect 11931 4576 12173 4604
rect 11931 4573 11943 4576
rect 11885 4567 11943 4573
rect 12161 4573 12173 4576
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4604 17739 4607
rect 18322 4604 18328 4616
rect 17727 4576 18328 4604
rect 17727 4573 17739 4576
rect 17681 4567 17739 4573
rect 18322 4564 18328 4576
rect 18380 4564 18386 4616
rect 18598 4564 18604 4616
rect 18656 4604 18662 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 18656 4576 19441 4604
rect 18656 4564 18662 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 21266 4564 21272 4616
rect 21324 4564 21330 4616
rect 22738 4564 22744 4616
rect 22796 4604 22802 4616
rect 24029 4607 24087 4613
rect 24029 4604 24041 4607
rect 22796 4576 24041 4604
rect 22796 4564 22802 4576
rect 24029 4573 24041 4576
rect 24075 4573 24087 4607
rect 24029 4567 24087 4573
rect 7650 4496 7656 4548
rect 7708 4496 7714 4548
rect 7834 4496 7840 4548
rect 7892 4536 7898 4548
rect 8941 4539 8999 4545
rect 8941 4536 8953 4539
rect 7892 4508 8953 4536
rect 7892 4496 7898 4508
rect 8941 4505 8953 4508
rect 8987 4505 8999 4539
rect 8941 4499 8999 4505
rect 9030 4496 9036 4548
rect 9088 4536 9094 4548
rect 10137 4539 10195 4545
rect 10137 4536 10149 4539
rect 9088 4508 10149 4536
rect 9088 4496 9094 4508
rect 10137 4505 10149 4508
rect 10183 4505 10195 4539
rect 10137 4499 10195 4505
rect 18693 4539 18751 4545
rect 18693 4505 18705 4539
rect 18739 4536 18751 4539
rect 20162 4536 20168 4548
rect 18739 4508 20168 4536
rect 18739 4505 18751 4508
rect 18693 4499 18751 4505
rect 20162 4496 20168 4508
rect 20220 4496 20226 4548
rect 23382 4496 23388 4548
rect 23440 4536 23446 4548
rect 24673 4539 24731 4545
rect 24673 4536 24685 4539
rect 23440 4508 24685 4536
rect 23440 4496 23446 4508
rect 24673 4505 24685 4508
rect 24719 4505 24731 4539
rect 24673 4499 24731 4505
rect 1762 4428 1768 4480
rect 1820 4468 1826 4480
rect 2225 4471 2283 4477
rect 2225 4468 2237 4471
rect 1820 4440 2237 4468
rect 1820 4428 1826 4440
rect 2225 4437 2237 4440
rect 2271 4437 2283 4471
rect 2225 4431 2283 4437
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 6604 4440 7113 4468
rect 6604 4428 6610 4440
rect 7101 4437 7113 4440
rect 7147 4437 7159 4471
rect 7101 4431 7159 4437
rect 8478 4428 8484 4480
rect 8536 4468 8542 4480
rect 9125 4471 9183 4477
rect 9125 4468 9137 4471
rect 8536 4440 9137 4468
rect 8536 4428 8542 4440
rect 9125 4437 9137 4440
rect 9171 4437 9183 4471
rect 9125 4431 9183 4437
rect 10226 4428 10232 4480
rect 10284 4468 10290 4480
rect 10321 4471 10379 4477
rect 10321 4468 10333 4471
rect 10284 4440 10333 4468
rect 10284 4428 10290 4440
rect 10321 4437 10333 4440
rect 10367 4437 10379 4471
rect 10321 4431 10379 4437
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 1762 4088 1768 4140
rect 1820 4088 1826 4140
rect 2406 4088 2412 4140
rect 2464 4088 2470 4140
rect 2961 4131 3019 4137
rect 2961 4097 2973 4131
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 4617 4131 4675 4137
rect 4617 4128 4629 4131
rect 3743 4100 4629 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 2976 4060 3004 4091
rect 4341 4063 4399 4069
rect 4341 4060 4353 4063
rect 2976 4032 4353 4060
rect 4341 4029 4353 4032
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 3878 3952 3884 4004
rect 3936 3992 3942 4004
rect 4448 3992 4476 4100
rect 4617 4097 4629 4100
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 5350 4088 5356 4140
rect 5408 4088 5414 4140
rect 5994 4088 6000 4140
rect 6052 4088 6058 4140
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 7190 4088 7196 4140
rect 7248 4088 7254 4140
rect 7929 4131 7987 4137
rect 7929 4097 7941 4131
rect 7975 4128 7987 4131
rect 8570 4128 8576 4140
rect 7975 4100 8576 4128
rect 7975 4097 7987 4100
rect 7929 4091 7987 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 8680 4060 8708 4091
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 10321 4131 10379 4137
rect 10321 4128 10333 4131
rect 9456 4100 10333 4128
rect 9456 4088 9462 4100
rect 10321 4097 10333 4100
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11296 4100 11713 4128
rect 11296 4088 11302 4100
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 13630 4088 13636 4140
rect 13688 4088 13694 4140
rect 16114 4088 16120 4140
rect 16172 4088 16178 4140
rect 16666 4088 16672 4140
rect 16724 4128 16730 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16724 4100 16865 4128
rect 16724 4088 16730 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 18690 4088 18696 4140
rect 18748 4088 18754 4140
rect 20254 4088 20260 4140
rect 20312 4128 20318 4140
rect 22094 4128 22100 4140
rect 20312 4100 22100 4128
rect 20312 4088 20318 4100
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 22189 4131 22247 4137
rect 22189 4097 22201 4131
rect 22235 4128 22247 4131
rect 22370 4128 22376 4140
rect 22235 4100 22376 4128
rect 22235 4097 22247 4100
rect 22189 4091 22247 4097
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 24121 4131 24179 4137
rect 24121 4097 24133 4131
rect 24167 4128 24179 4131
rect 24670 4128 24676 4140
rect 24167 4100 24676 4128
rect 24167 4097 24179 4100
rect 24121 4091 24179 4097
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 8680 4032 10057 4060
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 13504 4032 14013 4060
rect 13504 4020 13510 4032
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16448 4032 17325 4060
rect 16448 4020 16454 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 17552 4032 19165 4060
rect 17552 4020 17558 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 20070 4020 20076 4072
rect 20128 4060 20134 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 20128 4032 22477 4060
rect 20128 4020 20134 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 24762 4020 24768 4072
rect 24820 4020 24826 4072
rect 5442 3992 5448 4004
rect 3936 3964 4476 3992
rect 4540 3964 5448 3992
rect 3936 3952 3942 3964
rect 1486 3884 1492 3936
rect 1544 3884 1550 3936
rect 3145 3927 3203 3933
rect 3145 3893 3157 3927
rect 3191 3924 3203 3927
rect 4540 3924 4568 3964
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 6914 3952 6920 4004
rect 6972 3992 6978 4004
rect 8113 3995 8171 4001
rect 8113 3992 8125 3995
rect 6972 3964 8125 3992
rect 6972 3952 6978 3964
rect 8113 3961 8125 3964
rect 8159 3961 8171 3995
rect 8113 3955 8171 3961
rect 8846 3952 8852 4004
rect 8904 3952 8910 4004
rect 10318 3952 10324 4004
rect 10376 3992 10382 4004
rect 11057 3995 11115 4001
rect 11057 3992 11069 3995
rect 10376 3964 11069 3992
rect 10376 3952 10382 3964
rect 11057 3961 11069 3964
rect 11103 3961 11115 3995
rect 11057 3955 11115 3961
rect 20714 3952 20720 4004
rect 20772 3992 20778 4004
rect 24946 3992 24952 4004
rect 20772 3964 24952 3992
rect 20772 3952 20778 3964
rect 24946 3952 24952 3964
rect 25004 3952 25010 4004
rect 3191 3896 4568 3924
rect 3191 3893 3203 3896
rect 3145 3887 3203 3893
rect 4890 3884 4896 3936
rect 4948 3884 4954 3936
rect 5077 3927 5135 3933
rect 5077 3893 5089 3927
rect 5123 3924 5135 3927
rect 5534 3924 5540 3936
rect 5123 3896 5540 3924
rect 5123 3893 5135 3896
rect 5077 3887 5135 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 6822 3884 6828 3936
rect 6880 3924 6886 3936
rect 7561 3927 7619 3933
rect 7561 3924 7573 3927
rect 6880 3896 7573 3924
rect 6880 3884 6886 3896
rect 7561 3893 7573 3896
rect 7607 3893 7619 3927
rect 7561 3887 7619 3893
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 10100 3896 10517 3924
rect 10100 3884 10106 3896
rect 10505 3893 10517 3896
rect 10551 3893 10563 3927
rect 10505 3887 10563 3893
rect 10870 3884 10876 3936
rect 10928 3884 10934 3936
rect 11238 3884 11244 3936
rect 11296 3884 11302 3936
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 11756 3896 12357 3924
rect 11756 3884 11762 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12345 3887 12403 3893
rect 16209 3927 16267 3933
rect 16209 3893 16221 3927
rect 16255 3924 16267 3927
rect 22554 3924 22560 3936
rect 16255 3896 22560 3924
rect 16255 3893 16267 3896
rect 16209 3887 16267 3893
rect 22554 3884 22560 3896
rect 22612 3884 22618 3936
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 1854 3680 1860 3732
rect 1912 3720 1918 3732
rect 2317 3723 2375 3729
rect 2317 3720 2329 3723
rect 1912 3692 2329 3720
rect 1912 3680 1918 3692
rect 2317 3689 2329 3692
rect 2363 3689 2375 3723
rect 2317 3683 2375 3689
rect 2866 3680 2872 3732
rect 2924 3720 2930 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 2924 3692 3433 3720
rect 2924 3680 2930 3692
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 3421 3683 3479 3689
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 5261 3723 5319 3729
rect 5261 3720 5273 3723
rect 5040 3692 5273 3720
rect 5040 3680 5046 3692
rect 5261 3689 5273 3692
rect 5307 3689 5319 3723
rect 5261 3683 5319 3689
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 6365 3723 6423 3729
rect 6365 3720 6377 3723
rect 5776 3692 6377 3720
rect 5776 3680 5782 3692
rect 6365 3689 6377 3692
rect 6411 3689 6423 3723
rect 6365 3683 6423 3689
rect 8570 3680 8576 3732
rect 8628 3680 8634 3732
rect 9306 3680 9312 3732
rect 9364 3680 9370 3732
rect 12526 3680 12532 3732
rect 12584 3720 12590 3732
rect 12710 3720 12716 3732
rect 12584 3692 12716 3720
rect 12584 3680 12590 3692
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 18601 3723 18659 3729
rect 18601 3689 18613 3723
rect 18647 3720 18659 3723
rect 18690 3720 18696 3732
rect 18647 3692 18696 3720
rect 18647 3689 18659 3692
rect 18601 3683 18659 3689
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 3973 3655 4031 3661
rect 3973 3621 3985 3655
rect 4019 3652 4031 3655
rect 16114 3652 16120 3664
rect 4019 3624 16120 3652
rect 4019 3621 4031 3624
rect 3973 3615 4031 3621
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 18966 3612 18972 3664
rect 19024 3652 19030 3664
rect 19024 3624 21772 3652
rect 19024 3612 19030 3624
rect 10870 3544 10876 3596
rect 10928 3584 10934 3596
rect 10965 3587 11023 3593
rect 10965 3584 10977 3587
rect 10928 3556 10977 3584
rect 10928 3544 10934 3556
rect 10965 3553 10977 3556
rect 11011 3553 11023 3587
rect 10965 3547 11023 3553
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3584 11299 3587
rect 11287 3556 12664 3584
rect 11287 3553 11299 3556
rect 11241 3547 11299 3553
rect 1486 3476 1492 3528
rect 1544 3516 1550 3528
rect 1673 3519 1731 3525
rect 1673 3516 1685 3519
rect 1544 3488 1685 3516
rect 1544 3476 1550 3488
rect 1673 3485 1685 3488
rect 1719 3516 1731 3519
rect 2038 3516 2044 3528
rect 1719 3488 2044 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 2038 3476 2044 3488
rect 2096 3476 2102 3528
rect 2774 3476 2780 3528
rect 2832 3476 2838 3528
rect 4154 3476 4160 3528
rect 4212 3476 4218 3528
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 4982 3516 4988 3528
rect 4663 3488 4988 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 5718 3476 5724 3528
rect 5776 3476 5782 3528
rect 6822 3476 6828 3528
rect 6880 3476 6886 3528
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 7892 3488 7941 3516
rect 7892 3476 7898 3488
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9140 3448 9168 3479
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9824 3488 9873 3516
rect 9824 3476 9830 3488
rect 9861 3485 9873 3488
rect 9907 3516 9919 3519
rect 10042 3516 10048 3528
rect 9907 3488 10048 3516
rect 9907 3485 9919 3488
rect 9861 3479 9919 3485
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 12526 3476 12532 3528
rect 12584 3476 12590 3528
rect 12636 3516 12664 3556
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 12805 3587 12863 3593
rect 12805 3584 12817 3587
rect 12768 3556 12817 3584
rect 12768 3544 12774 3556
rect 12805 3553 12817 3556
rect 12851 3553 12863 3587
rect 12805 3547 12863 3553
rect 14918 3544 14924 3596
rect 14976 3584 14982 3596
rect 15473 3587 15531 3593
rect 15473 3584 15485 3587
rect 14976 3556 15485 3584
rect 14976 3544 14982 3556
rect 15473 3553 15485 3556
rect 15519 3553 15531 3587
rect 15473 3547 15531 3553
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 16080 3556 17325 3584
rect 16080 3544 16086 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 17862 3544 17868 3596
rect 17920 3584 17926 3596
rect 21744 3593 21772 3624
rect 19889 3587 19947 3593
rect 19889 3584 19901 3587
rect 17920 3556 19901 3584
rect 17920 3544 17926 3556
rect 19889 3553 19901 3556
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 14826 3516 14832 3528
rect 12636 3488 14832 3516
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3516 15163 3519
rect 15562 3516 15568 3528
rect 15151 3488 15568 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 10505 3451 10563 3457
rect 10505 3448 10517 3451
rect 9140 3420 10517 3448
rect 10505 3417 10517 3420
rect 10551 3417 10563 3451
rect 10505 3411 10563 3417
rect 15470 3408 15476 3460
rect 15528 3448 15534 3460
rect 16868 3448 16896 3479
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 17460 3488 19441 3516
rect 17460 3476 17466 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3516 21511 3519
rect 21634 3516 21640 3528
rect 21499 3488 21640 3516
rect 21499 3485 21511 3488
rect 21453 3479 21511 3485
rect 21634 3476 21640 3488
rect 21692 3476 21698 3528
rect 23106 3476 23112 3528
rect 23164 3516 23170 3528
rect 23385 3519 23443 3525
rect 23385 3516 23397 3519
rect 23164 3488 23397 3516
rect 23164 3476 23170 3488
rect 23385 3485 23397 3488
rect 23431 3485 23443 3519
rect 23385 3479 23443 3485
rect 24029 3519 24087 3525
rect 24029 3485 24041 3519
rect 24075 3516 24087 3519
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 24075 3488 24593 3516
rect 24075 3485 24087 3488
rect 24029 3479 24087 3485
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 15528 3420 16896 3448
rect 15528 3408 15534 3420
rect 19702 3408 19708 3460
rect 19760 3448 19766 3460
rect 21726 3448 21732 3460
rect 19760 3420 21732 3448
rect 19760 3408 19766 3420
rect 21726 3408 21732 3420
rect 21784 3408 21790 3460
rect 4614 3340 4620 3392
rect 4672 3380 4678 3392
rect 7469 3383 7527 3389
rect 7469 3380 7481 3383
rect 4672 3352 7481 3380
rect 4672 3340 4678 3352
rect 7469 3349 7481 3352
rect 7515 3349 7527 3383
rect 7469 3343 7527 3349
rect 18598 3340 18604 3392
rect 18656 3380 18662 3392
rect 19886 3380 19892 3392
rect 18656 3352 19892 3380
rect 18656 3340 18662 3352
rect 19886 3340 19892 3352
rect 19944 3340 19950 3392
rect 21818 3340 21824 3392
rect 21876 3380 21882 3392
rect 22830 3380 22836 3392
rect 21876 3352 22836 3380
rect 21876 3340 21882 3352
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 24578 3340 24584 3392
rect 24636 3380 24642 3392
rect 25225 3383 25283 3389
rect 25225 3380 25237 3383
rect 24636 3352 25237 3380
rect 24636 3340 24642 3352
rect 25225 3349 25237 3352
rect 25271 3349 25283 3383
rect 25225 3343 25283 3349
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 2866 3176 2872 3188
rect 2823 3148 2872 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 5997 3179 6055 3185
rect 5997 3176 6009 3179
rect 4212 3148 6009 3176
rect 4212 3136 4218 3148
rect 5997 3145 6009 3148
rect 6043 3145 6055 3179
rect 5997 3139 6055 3145
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 8573 3179 8631 3185
rect 8573 3176 8585 3179
rect 8352 3148 8585 3176
rect 8352 3136 8358 3148
rect 8573 3145 8585 3148
rect 8619 3145 8631 3179
rect 8573 3139 8631 3145
rect 11885 3179 11943 3185
rect 11885 3145 11897 3179
rect 11931 3176 11943 3179
rect 13354 3176 13360 3188
rect 11931 3148 13360 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 21450 3136 21456 3188
rect 21508 3176 21514 3188
rect 22646 3176 22652 3188
rect 21508 3148 22652 3176
rect 21508 3136 21514 3148
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 23106 3136 23112 3188
rect 23164 3136 23170 3188
rect 24854 3136 24860 3188
rect 24912 3176 24918 3188
rect 25133 3179 25191 3185
rect 25133 3176 25145 3179
rect 24912 3148 25145 3176
rect 24912 3136 24918 3148
rect 25133 3145 25145 3148
rect 25179 3145 25191 3179
rect 25133 3139 25191 3145
rect 13722 3108 13728 3120
rect 10612 3080 13728 3108
rect 2130 3000 2136 3052
rect 2188 3040 2194 3052
rect 2406 3040 2412 3052
rect 2188 3012 2412 3040
rect 2188 3000 2194 3012
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 4614 3000 4620 3052
rect 4672 3000 4678 3052
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 5534 3040 5540 3052
rect 5399 3012 5540 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 5534 3000 5540 3012
rect 5592 3040 5598 3052
rect 6086 3040 6092 3052
rect 5592 3012 6092 3040
rect 5592 3000 5598 3012
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6595 3012 6837 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 6825 3009 6837 3012
rect 6871 3040 6883 3043
rect 7190 3040 7196 3052
rect 6871 3012 7196 3040
rect 6871 3009 6883 3012
rect 6825 3003 6883 3009
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3040 7987 3043
rect 8478 3040 8484 3052
rect 7975 3012 8484 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3040 9367 3043
rect 9582 3040 9588 3052
rect 9355 3012 9588 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10502 3040 10508 3052
rect 10376 3012 10508 3040
rect 10376 3000 10382 3012
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 10612 3049 10640 3080
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 11698 3000 11704 3052
rect 11756 3000 11762 3052
rect 12621 3043 12679 3049
rect 12621 3009 12633 3043
rect 12667 3040 12679 3043
rect 13538 3040 13544 3052
rect 12667 3012 13544 3040
rect 12667 3009 12679 3012
rect 12621 3003 12679 3009
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 14274 3000 14280 3052
rect 14332 3000 14338 3052
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 18782 3000 18788 3052
rect 18840 3000 18846 3052
rect 22465 3043 22523 3049
rect 22465 3009 22477 3043
rect 22511 3040 22523 3043
rect 22511 3012 23520 3040
rect 22511 3009 22523 3012
rect 22465 3003 22523 3009
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 2774 2972 2780 2984
rect 1903 2944 2780 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2972 3295 2975
rect 3326 2972 3332 2984
rect 3283 2944 3332 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 1489 2907 1547 2913
rect 1489 2873 1501 2907
rect 1535 2904 1547 2907
rect 3252 2904 3280 2935
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 10134 2972 10140 2984
rect 3559 2944 10140 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 13354 2932 13360 2984
rect 13412 2932 13418 2984
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14240 2944 14749 2972
rect 14240 2932 14246 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15712 2944 17325 2972
rect 15712 2932 15718 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 1535 2876 3280 2904
rect 1535 2873 1547 2876
rect 1489 2867 1547 2873
rect 4798 2864 4804 2916
rect 4856 2864 4862 2916
rect 17126 2864 17132 2916
rect 17184 2904 17190 2916
rect 19168 2904 19196 2935
rect 20162 2932 20168 2984
rect 20220 2972 20226 2984
rect 23382 2972 23388 2984
rect 20220 2944 23388 2972
rect 20220 2932 20226 2944
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 17184 2876 19196 2904
rect 17184 2864 17190 2876
rect 1673 2839 1731 2845
rect 1673 2805 1685 2839
rect 1719 2836 1731 2839
rect 4706 2836 4712 2848
rect 1719 2808 4712 2836
rect 1719 2805 1731 2808
rect 1673 2799 1731 2805
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 7466 2796 7472 2848
rect 7524 2796 7530 2848
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 17954 2836 17960 2848
rect 16816 2808 17960 2836
rect 16816 2796 16822 2808
rect 17954 2796 17960 2808
rect 18012 2796 18018 2848
rect 20806 2796 20812 2848
rect 20864 2836 20870 2848
rect 22462 2836 22468 2848
rect 20864 2808 22468 2836
rect 20864 2796 20870 2808
rect 22462 2796 22468 2808
rect 22520 2796 22526 2848
rect 23492 2845 23520 3012
rect 25314 3000 25320 3052
rect 25372 3000 25378 3052
rect 23477 2839 23535 2845
rect 23477 2805 23489 2839
rect 23523 2836 23535 2839
rect 24118 2836 24124 2848
rect 23523 2808 24124 2836
rect 23523 2805 23535 2808
rect 23477 2799 23535 2805
rect 24118 2796 24124 2808
rect 24176 2796 24182 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 2314 2592 2320 2644
rect 2372 2592 2378 2644
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 3970 2632 3976 2644
rect 3467 2604 3976 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 7466 2632 7472 2644
rect 4908 2604 7472 2632
rect 3510 2496 3516 2508
rect 1688 2468 3516 2496
rect 1688 2437 1716 2468
rect 3510 2456 3516 2468
rect 3568 2496 3574 2508
rect 3786 2496 3792 2508
rect 3568 2468 3792 2496
rect 3568 2456 3574 2468
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 4908 2496 4936 2604
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 9858 2592 9864 2644
rect 9916 2592 9922 2644
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 15930 2632 15936 2644
rect 11747 2604 15936 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 18601 2635 18659 2641
rect 18601 2601 18613 2635
rect 18647 2632 18659 2635
rect 18782 2632 18788 2644
rect 18647 2604 18788 2632
rect 18647 2601 18659 2604
rect 18601 2595 18659 2601
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 25225 2635 25283 2641
rect 25225 2601 25237 2635
rect 25271 2632 25283 2635
rect 25314 2632 25320 2644
rect 25271 2604 25320 2632
rect 25271 2601 25283 2604
rect 25225 2595 25283 2601
rect 25314 2592 25320 2604
rect 25372 2592 25378 2644
rect 7098 2564 7104 2576
rect 5000 2536 7104 2564
rect 5000 2505 5028 2536
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 7193 2567 7251 2573
rect 7193 2533 7205 2567
rect 7239 2564 7251 2567
rect 7650 2564 7656 2576
rect 7239 2536 7656 2564
rect 7239 2533 7251 2536
rect 7193 2527 7251 2533
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 12342 2564 12348 2576
rect 10336 2536 12348 2564
rect 10336 2505 10364 2536
rect 12342 2524 12348 2536
rect 12400 2564 12406 2576
rect 14277 2567 14335 2573
rect 14277 2564 14289 2567
rect 12400 2536 14289 2564
rect 12400 2524 12406 2536
rect 14277 2533 14289 2536
rect 14323 2533 14335 2567
rect 14277 2527 14335 2533
rect 17678 2524 17684 2576
rect 17736 2564 17742 2576
rect 17736 2536 22048 2564
rect 17736 2524 17742 2536
rect 3988 2468 4936 2496
rect 4985 2499 5043 2505
rect 3988 2437 4016 2468
rect 4985 2465 4997 2499
rect 5031 2465 5043 2499
rect 4985 2459 5043 2465
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2496 6055 2499
rect 10321 2499 10379 2505
rect 6043 2468 7604 2496
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 7576 2440 7604 2468
rect 10321 2465 10333 2499
rect 10367 2465 10379 2499
rect 11974 2496 11980 2508
rect 10321 2459 10379 2465
rect 11900 2468 11980 2496
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2397 1731 2431
rect 1673 2391 1731 2397
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2397 2835 2431
rect 2777 2391 2835 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 2792 2360 2820 2391
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 7374 2428 7380 2440
rect 6595 2400 7380 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 7374 2388 7380 2400
rect 7432 2428 7438 2440
rect 7432 2400 7512 2428
rect 7432 2388 7438 2400
rect 3602 2360 3608 2372
rect 2792 2332 3608 2360
rect 3602 2320 3608 2332
rect 3660 2360 3666 2372
rect 4062 2360 4068 2372
rect 3660 2332 4068 2360
rect 3660 2320 3666 2332
rect 4062 2320 4068 2332
rect 4120 2320 4126 2372
rect 7282 2360 7288 2372
rect 4172 2332 7288 2360
rect 4172 2301 4200 2332
rect 7282 2320 7288 2332
rect 7340 2320 7346 2372
rect 7484 2360 7512 2400
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7616 2400 7665 2428
rect 7616 2388 7622 2400
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2428 7987 2431
rect 9217 2431 9275 2437
rect 7975 2400 9168 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8202 2360 8208 2372
rect 7484 2332 8208 2360
rect 8202 2320 8208 2332
rect 8260 2320 8266 2372
rect 9140 2360 9168 2400
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 10226 2428 10232 2440
rect 9263 2400 10232 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 10226 2388 10232 2400
rect 10284 2388 10290 2440
rect 11900 2437 11928 2468
rect 11974 2456 11980 2468
rect 12032 2496 12038 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 12032 2468 14105 2496
rect 12032 2456 12038 2468
rect 14093 2465 14105 2468
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 14608 2468 15209 2496
rect 14608 2456 14614 2468
rect 15197 2465 15209 2468
rect 15243 2465 15255 2499
rect 15197 2459 15255 2465
rect 15286 2456 15292 2508
rect 15344 2496 15350 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 15344 2468 17325 2496
rect 15344 2456 15350 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 18012 2468 19901 2496
rect 18012 2456 18018 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 10612 2360 10640 2391
rect 12434 2388 12440 2440
rect 12492 2388 12498 2440
rect 14642 2388 14648 2440
rect 14700 2388 14706 2440
rect 16850 2388 16856 2440
rect 16908 2388 16914 2440
rect 19518 2388 19524 2440
rect 19576 2388 19582 2440
rect 22020 2437 22048 2536
rect 22465 2499 22523 2505
rect 22465 2465 22477 2499
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 24029 2499 24087 2505
rect 24029 2465 24041 2499
rect 24075 2496 24087 2499
rect 24854 2496 24860 2508
rect 24075 2468 24860 2496
rect 24075 2465 24087 2468
rect 24029 2459 24087 2465
rect 22005 2431 22063 2437
rect 22005 2397 22017 2431
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 12618 2360 12624 2372
rect 9140 2332 10548 2360
rect 10612 2332 12624 2360
rect 4157 2295 4215 2301
rect 4157 2261 4169 2295
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 5718 2252 5724 2304
rect 5776 2292 5782 2304
rect 6089 2295 6147 2301
rect 6089 2292 6101 2295
rect 5776 2264 6101 2292
rect 5776 2252 5782 2264
rect 6089 2261 6101 2264
rect 6135 2261 6147 2295
rect 6089 2255 6147 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 10410 2292 10416 2304
rect 7156 2264 10416 2292
rect 7156 2252 7162 2264
rect 10410 2252 10416 2264
rect 10468 2252 10474 2304
rect 10520 2292 10548 2332
rect 12618 2320 12624 2332
rect 12676 2320 12682 2372
rect 13541 2363 13599 2369
rect 13541 2329 13553 2363
rect 13587 2360 13599 2363
rect 13814 2360 13820 2372
rect 13587 2332 13820 2360
rect 13587 2329 13599 2332
rect 13541 2323 13599 2329
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 18322 2320 18328 2372
rect 18380 2360 18386 2372
rect 22480 2360 22508 2459
rect 24854 2456 24860 2468
rect 24912 2456 24918 2508
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 18380 2332 22508 2360
rect 18380 2320 18386 2332
rect 15010 2292 15016 2304
rect 10520 2264 15016 2292
rect 15010 2252 15016 2264
rect 15068 2252 15074 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 7282 2048 7288 2100
rect 7340 2088 7346 2100
rect 11790 2088 11796 2100
rect 7340 2060 11796 2088
rect 7340 2048 7346 2060
rect 11790 2048 11796 2060
rect 11848 2048 11854 2100
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 3976 54315 4028 54324
rect 3976 54281 3985 54315
rect 3985 54281 4019 54315
rect 4019 54281 4028 54315
rect 3976 54272 4028 54281
rect 9956 54272 10008 54324
rect 14004 54272 14056 54324
rect 14740 54272 14792 54324
rect 7840 54204 7892 54256
rect 11428 54204 11480 54256
rect 2320 54136 2372 54188
rect 4620 54179 4672 54188
rect 4620 54145 4629 54179
rect 4629 54145 4663 54179
rect 4663 54145 4672 54179
rect 4620 54136 4672 54145
rect 5908 54068 5960 54120
rect 9956 54179 10008 54188
rect 9956 54145 9965 54179
rect 9965 54145 9999 54179
rect 9999 54145 10008 54179
rect 9956 54136 10008 54145
rect 11612 54136 11664 54188
rect 12900 54204 12952 54256
rect 13636 54204 13688 54256
rect 12348 54179 12400 54188
rect 12348 54145 12357 54179
rect 12357 54145 12391 54179
rect 12391 54145 12400 54179
rect 12348 54136 12400 54145
rect 15568 54204 15620 54256
rect 17408 54136 17460 54188
rect 17960 54179 18012 54188
rect 17960 54145 17969 54179
rect 17969 54145 18003 54179
rect 18003 54145 18012 54179
rect 17960 54136 18012 54145
rect 19432 54179 19484 54188
rect 19432 54145 19441 54179
rect 19441 54145 19475 54179
rect 19475 54145 19484 54179
rect 19432 54136 19484 54145
rect 11244 54068 11296 54120
rect 12532 54068 12584 54120
rect 18696 54068 18748 54120
rect 19156 54068 19208 54120
rect 20720 54136 20772 54188
rect 21364 54068 21416 54120
rect 24032 54136 24084 54188
rect 24676 54136 24728 54188
rect 20536 54000 20588 54052
rect 25044 54000 25096 54052
rect 3792 53975 3844 53984
rect 3792 53941 3801 53975
rect 3801 53941 3835 53975
rect 3835 53941 3844 53975
rect 3792 53932 3844 53941
rect 12716 53932 12768 53984
rect 15292 53932 15344 53984
rect 17500 53975 17552 53984
rect 17500 53941 17509 53975
rect 17509 53941 17543 53975
rect 17543 53941 17552 53975
rect 17500 53932 17552 53941
rect 18604 53975 18656 53984
rect 18604 53941 18613 53975
rect 18613 53941 18647 53975
rect 18647 53941 18656 53975
rect 18604 53932 18656 53941
rect 19340 53932 19392 53984
rect 21180 53975 21232 53984
rect 21180 53941 21189 53975
rect 21189 53941 21223 53975
rect 21223 53941 21232 53975
rect 21180 53932 21232 53941
rect 22100 53932 22152 53984
rect 23756 53975 23808 53984
rect 23756 53941 23765 53975
rect 23765 53941 23799 53975
rect 23799 53941 23808 53975
rect 23756 53932 23808 53941
rect 23848 53932 23900 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 16580 53728 16632 53780
rect 17960 53728 18012 53780
rect 18420 53728 18472 53780
rect 2228 53660 2280 53712
rect 3424 53660 3476 53712
rect 5540 53660 5592 53712
rect 17684 53660 17736 53712
rect 7380 53592 7432 53644
rect 8852 53592 8904 53644
rect 11060 53635 11112 53644
rect 11060 53601 11069 53635
rect 11069 53601 11103 53635
rect 11103 53601 11112 53635
rect 11060 53592 11112 53601
rect 12164 53592 12216 53644
rect 18696 53635 18748 53644
rect 18696 53601 18705 53635
rect 18705 53601 18739 53635
rect 18739 53601 18748 53635
rect 18696 53592 18748 53601
rect 2228 53567 2280 53576
rect 2228 53533 2237 53567
rect 2237 53533 2271 53567
rect 2271 53533 2280 53567
rect 2228 53524 2280 53533
rect 3976 53567 4028 53576
rect 3976 53533 3985 53567
rect 3985 53533 4019 53567
rect 4019 53533 4028 53567
rect 3976 53524 4028 53533
rect 6828 53524 6880 53576
rect 8668 53524 8720 53576
rect 12072 53524 12124 53576
rect 12624 53524 12676 53576
rect 14004 53524 14056 53576
rect 15108 53524 15160 53576
rect 16212 53524 16264 53576
rect 16948 53524 17000 53576
rect 17684 53567 17736 53576
rect 17684 53533 17693 53567
rect 17693 53533 17727 53567
rect 17727 53533 17736 53567
rect 17684 53524 17736 53533
rect 6552 53388 6604 53440
rect 14280 53388 14332 53440
rect 15568 53388 15620 53440
rect 16856 53388 16908 53440
rect 17592 53388 17644 53440
rect 22652 53660 22704 53712
rect 22468 53592 22520 53644
rect 19524 53524 19576 53576
rect 20536 53567 20588 53576
rect 20536 53533 20545 53567
rect 20545 53533 20579 53567
rect 20579 53533 20588 53567
rect 20536 53524 20588 53533
rect 20996 53524 21048 53576
rect 21456 53524 21508 53576
rect 22192 53456 22244 53508
rect 24584 53524 24636 53576
rect 25964 53524 26016 53576
rect 19432 53388 19484 53440
rect 20168 53388 20220 53440
rect 20904 53388 20956 53440
rect 22008 53388 22060 53440
rect 23480 53388 23532 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 11612 53227 11664 53236
rect 11612 53193 11621 53227
rect 11621 53193 11655 53227
rect 11655 53193 11664 53227
rect 11612 53184 11664 53193
rect 17408 53227 17460 53236
rect 17408 53193 17417 53227
rect 17417 53193 17451 53227
rect 17451 53193 17460 53227
rect 17408 53184 17460 53193
rect 17684 53227 17736 53236
rect 17684 53193 17693 53227
rect 17693 53193 17727 53227
rect 17727 53193 17736 53227
rect 17684 53184 17736 53193
rect 4436 53116 4488 53168
rect 6276 53116 6328 53168
rect 9220 53116 9272 53168
rect 13360 53116 13412 53168
rect 17500 53116 17552 53168
rect 4528 53048 4580 53100
rect 4712 53091 4764 53100
rect 4712 53057 4721 53091
rect 4721 53057 4755 53091
rect 4755 53057 4764 53091
rect 4712 53048 4764 53057
rect 6552 53091 6604 53100
rect 6552 53057 6561 53091
rect 6561 53057 6595 53091
rect 6595 53057 6604 53091
rect 6552 53048 6604 53057
rect 7564 53048 7616 53100
rect 9312 53048 9364 53100
rect 11888 53091 11940 53100
rect 11888 53057 11897 53091
rect 11897 53057 11931 53091
rect 11931 53057 11940 53091
rect 11888 53048 11940 53057
rect 13636 53048 13688 53100
rect 14832 53091 14884 53100
rect 14832 53057 14841 53091
rect 14841 53057 14875 53091
rect 14875 53057 14884 53091
rect 14832 53048 14884 53057
rect 18604 53116 18656 53168
rect 19340 53159 19392 53168
rect 19340 53125 19349 53159
rect 19349 53125 19383 53159
rect 19383 53125 19392 53159
rect 19340 53116 19392 53125
rect 18328 53048 18380 53100
rect 19892 53048 19944 53100
rect 22008 53091 22060 53100
rect 22008 53057 22017 53091
rect 22017 53057 22051 53091
rect 22051 53057 22060 53091
rect 22008 53048 22060 53057
rect 23756 53116 23808 53168
rect 23480 53091 23532 53100
rect 23480 53057 23489 53091
rect 23489 53057 23523 53091
rect 23523 53057 23532 53091
rect 23480 53048 23532 53057
rect 24768 53048 24820 53100
rect 25044 53091 25096 53100
rect 25044 53057 25053 53091
rect 25053 53057 25087 53091
rect 25087 53057 25096 53091
rect 25044 53048 25096 53057
rect 10324 53023 10376 53032
rect 10324 52989 10333 53023
rect 10333 52989 10367 53023
rect 10367 52989 10376 53023
rect 10324 52980 10376 52989
rect 11796 52980 11848 53032
rect 16396 52912 16448 52964
rect 21640 52912 21692 52964
rect 22744 52912 22796 52964
rect 1768 52844 1820 52896
rect 14372 52887 14424 52896
rect 14372 52853 14381 52887
rect 14381 52853 14415 52887
rect 14415 52853 14424 52887
rect 14372 52844 14424 52853
rect 14556 52844 14608 52896
rect 17040 52887 17092 52896
rect 17040 52853 17049 52887
rect 17049 52853 17083 52887
rect 17083 52853 17092 52887
rect 17040 52844 17092 52853
rect 18788 52887 18840 52896
rect 18788 52853 18797 52887
rect 18797 52853 18831 52887
rect 18831 52853 18840 52887
rect 18788 52844 18840 52853
rect 19432 52887 19484 52896
rect 19432 52853 19441 52887
rect 19441 52853 19475 52887
rect 19475 52853 19484 52887
rect 19432 52844 19484 52853
rect 22560 52844 22612 52896
rect 23664 52887 23716 52896
rect 23664 52853 23673 52887
rect 23673 52853 23707 52887
rect 23707 52853 23716 52887
rect 23664 52844 23716 52853
rect 23940 52844 23992 52896
rect 24952 52844 25004 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 1860 52640 1912 52692
rect 3516 52640 3568 52692
rect 12624 52683 12676 52692
rect 12624 52649 12633 52683
rect 12633 52649 12667 52683
rect 12667 52649 12676 52683
rect 12624 52640 12676 52649
rect 14832 52683 14884 52692
rect 14832 52649 14841 52683
rect 14841 52649 14875 52683
rect 14875 52649 14884 52683
rect 14832 52640 14884 52649
rect 15108 52640 15160 52692
rect 16212 52640 16264 52692
rect 17132 52640 17184 52692
rect 21364 52640 21416 52692
rect 24032 52683 24084 52692
rect 24032 52649 24041 52683
rect 24041 52649 24075 52683
rect 24075 52649 24084 52683
rect 24032 52640 24084 52649
rect 24584 52640 24636 52692
rect 24768 52683 24820 52692
rect 24768 52649 24777 52683
rect 24777 52649 24811 52683
rect 24811 52649 24820 52683
rect 24768 52640 24820 52649
rect 1308 52572 1360 52624
rect 3792 52572 3844 52624
rect 3700 52504 3752 52556
rect 15660 52572 15712 52624
rect 21548 52572 21600 52624
rect 22468 52572 22520 52624
rect 25136 52572 25188 52624
rect 5172 52436 5224 52488
rect 5908 52436 5960 52488
rect 6644 52436 6696 52488
rect 7288 52479 7340 52488
rect 7288 52445 7297 52479
rect 7297 52445 7331 52479
rect 7331 52445 7340 52479
rect 7288 52436 7340 52445
rect 7748 52547 7800 52556
rect 7748 52513 7757 52547
rect 7757 52513 7791 52547
rect 7791 52513 7800 52547
rect 7748 52504 7800 52513
rect 10692 52504 10744 52556
rect 8576 52436 8628 52488
rect 9588 52436 9640 52488
rect 12808 52479 12860 52488
rect 12808 52445 12817 52479
rect 12817 52445 12851 52479
rect 12851 52445 12860 52479
rect 12808 52436 12860 52445
rect 13544 52436 13596 52488
rect 14280 52479 14332 52488
rect 14280 52445 14289 52479
rect 14289 52445 14323 52479
rect 14323 52445 14332 52479
rect 14280 52436 14332 52445
rect 15568 52479 15620 52488
rect 15568 52445 15577 52479
rect 15577 52445 15611 52479
rect 15611 52445 15620 52479
rect 15568 52436 15620 52445
rect 16856 52479 16908 52488
rect 16856 52445 16865 52479
rect 16865 52445 16899 52479
rect 16899 52445 16908 52479
rect 16856 52436 16908 52445
rect 17592 52479 17644 52488
rect 17592 52445 17601 52479
rect 17601 52445 17635 52479
rect 17635 52445 17644 52479
rect 17592 52436 17644 52445
rect 18788 52436 18840 52488
rect 21180 52504 21232 52556
rect 21732 52504 21784 52556
rect 20168 52479 20220 52488
rect 20168 52445 20177 52479
rect 20177 52445 20211 52479
rect 20211 52445 20220 52479
rect 20168 52436 20220 52445
rect 20904 52479 20956 52488
rect 20904 52445 20913 52479
rect 20913 52445 20947 52479
rect 20947 52445 20956 52479
rect 20904 52436 20956 52445
rect 22100 52436 22152 52488
rect 22744 52436 22796 52488
rect 22928 52436 22980 52488
rect 23296 52436 23348 52488
rect 24768 52436 24820 52488
rect 14556 52368 14608 52420
rect 14464 52343 14516 52352
rect 14464 52309 14473 52343
rect 14473 52309 14507 52343
rect 14507 52309 14516 52343
rect 14464 52300 14516 52309
rect 15752 52343 15804 52352
rect 15752 52309 15761 52343
rect 15761 52309 15795 52343
rect 15795 52309 15804 52343
rect 15752 52300 15804 52309
rect 18512 52343 18564 52352
rect 18512 52309 18521 52343
rect 18521 52309 18555 52343
rect 18555 52309 18564 52343
rect 18512 52300 18564 52309
rect 19616 52343 19668 52352
rect 19616 52309 19625 52343
rect 19625 52309 19659 52343
rect 19659 52309 19668 52343
rect 19616 52300 19668 52309
rect 20352 52343 20404 52352
rect 20352 52309 20361 52343
rect 20361 52309 20395 52343
rect 20395 52309 20404 52343
rect 20352 52300 20404 52309
rect 21088 52343 21140 52352
rect 21088 52309 21097 52343
rect 21097 52309 21131 52343
rect 21131 52309 21140 52343
rect 21088 52300 21140 52309
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 4528 52096 4580 52148
rect 11888 52096 11940 52148
rect 12348 52139 12400 52148
rect 12348 52105 12357 52139
rect 12357 52105 12391 52139
rect 12391 52105 12400 52139
rect 12348 52096 12400 52105
rect 19892 52139 19944 52148
rect 19892 52105 19901 52139
rect 19901 52105 19935 52139
rect 19935 52105 19944 52139
rect 19892 52096 19944 52105
rect 21456 52139 21508 52148
rect 21456 52105 21465 52139
rect 21465 52105 21499 52139
rect 21499 52105 21508 52139
rect 21456 52096 21508 52105
rect 9128 52028 9180 52080
rect 14372 52028 14424 52080
rect 1676 52003 1728 52012
rect 1676 51969 1685 52003
rect 1685 51969 1719 52003
rect 1719 51969 1728 52003
rect 1676 51960 1728 51969
rect 3332 51935 3384 51944
rect 3332 51901 3341 51935
rect 3341 51901 3375 51935
rect 3375 51901 3384 51935
rect 3332 51892 3384 51901
rect 7196 51960 7248 52012
rect 4896 51892 4948 51944
rect 9680 52003 9732 52012
rect 9680 51969 9689 52003
rect 9689 51969 9723 52003
rect 9723 51969 9732 52003
rect 9680 51960 9732 51969
rect 10876 51960 10928 52012
rect 11980 51960 12032 52012
rect 14648 52003 14700 52012
rect 14648 51969 14657 52003
rect 14657 51969 14691 52003
rect 14691 51969 14700 52003
rect 14648 51960 14700 51969
rect 15844 51960 15896 52012
rect 17316 51960 17368 52012
rect 18880 51960 18932 52012
rect 20260 51960 20312 52012
rect 22836 51960 22888 52012
rect 23664 51960 23716 52012
rect 24676 52003 24728 52012
rect 24676 51969 24685 52003
rect 24685 51969 24719 52003
rect 24719 51969 24728 52003
rect 24676 51960 24728 51969
rect 8484 51935 8536 51944
rect 8484 51901 8493 51935
rect 8493 51901 8527 51935
rect 8527 51901 8536 51935
rect 8484 51892 8536 51901
rect 9772 51892 9824 51944
rect 10416 51824 10468 51876
rect 14096 51824 14148 51876
rect 15016 51824 15068 51876
rect 17224 51824 17276 51876
rect 18420 51824 18472 51876
rect 22744 51824 22796 51876
rect 3976 51756 4028 51808
rect 4896 51756 4948 51808
rect 18604 51756 18656 51808
rect 20168 51756 20220 51808
rect 22376 51756 22428 51808
rect 25780 51756 25832 51808
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 9956 51552 10008 51604
rect 2872 51459 2924 51468
rect 2872 51425 2881 51459
rect 2881 51425 2915 51459
rect 2915 51425 2924 51459
rect 2872 51416 2924 51425
rect 6920 51416 6972 51468
rect 7012 51416 7064 51468
rect 3976 51391 4028 51400
rect 3976 51357 3985 51391
rect 3985 51357 4019 51391
rect 4019 51357 4028 51391
rect 3976 51348 4028 51357
rect 5540 51348 5592 51400
rect 7104 51391 7156 51400
rect 7104 51357 7113 51391
rect 7113 51357 7147 51391
rect 7147 51357 7156 51391
rect 7104 51348 7156 51357
rect 9220 51348 9272 51400
rect 25044 51391 25096 51400
rect 25044 51357 25053 51391
rect 25053 51357 25087 51391
rect 25087 51357 25096 51391
rect 25044 51348 25096 51357
rect 6736 51280 6788 51332
rect 7012 51280 7064 51332
rect 7196 51280 7248 51332
rect 4252 51212 4304 51264
rect 25872 51212 25924 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 1676 51008 1728 51060
rect 6920 51051 6972 51060
rect 6920 51017 6929 51051
rect 6929 51017 6963 51051
rect 6963 51017 6972 51051
rect 6920 51008 6972 51017
rect 2320 50940 2372 50992
rect 1768 50915 1820 50924
rect 1768 50881 1777 50915
rect 1777 50881 1811 50915
rect 1811 50881 1820 50915
rect 1768 50872 1820 50881
rect 2780 50847 2832 50856
rect 2780 50813 2789 50847
rect 2789 50813 2823 50847
rect 2823 50813 2832 50847
rect 2780 50804 2832 50813
rect 5448 50872 5500 50924
rect 7656 50872 7708 50924
rect 9588 50983 9640 50992
rect 9588 50949 9597 50983
rect 9597 50949 9631 50983
rect 9631 50949 9640 50983
rect 9588 50940 9640 50949
rect 7840 50872 7892 50924
rect 25044 50915 25096 50924
rect 25044 50881 25053 50915
rect 25053 50881 25087 50915
rect 25087 50881 25096 50915
rect 25044 50872 25096 50881
rect 4344 50804 4396 50856
rect 7472 50847 7524 50856
rect 7472 50813 7481 50847
rect 7481 50813 7515 50847
rect 7515 50813 7524 50847
rect 7472 50804 7524 50813
rect 4160 50736 4212 50788
rect 25688 50668 25740 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 6828 50507 6880 50516
rect 6828 50473 6837 50507
rect 6837 50473 6871 50507
rect 6871 50473 6880 50507
rect 6828 50464 6880 50473
rect 8668 50464 8720 50516
rect 1308 50328 1360 50380
rect 3424 50328 3476 50380
rect 4436 50260 4488 50312
rect 5816 50260 5868 50312
rect 9404 50303 9456 50312
rect 9404 50269 9413 50303
rect 9413 50269 9447 50303
rect 9447 50269 9456 50303
rect 9404 50260 9456 50269
rect 5080 50192 5132 50244
rect 25320 50124 25372 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 3516 49852 3568 49904
rect 1952 49827 2004 49836
rect 1952 49793 1961 49827
rect 1961 49793 1995 49827
rect 1995 49793 2004 49827
rect 1952 49784 2004 49793
rect 9864 49920 9916 49972
rect 20996 49920 21048 49972
rect 4252 49895 4304 49904
rect 4252 49861 4261 49895
rect 4261 49861 4295 49895
rect 4295 49861 4304 49895
rect 4252 49852 4304 49861
rect 9036 49852 9088 49904
rect 9312 49895 9364 49904
rect 9312 49861 9321 49895
rect 9321 49861 9355 49895
rect 9355 49861 9364 49895
rect 9312 49852 9364 49861
rect 7748 49784 7800 49836
rect 25320 49827 25372 49836
rect 25320 49793 25329 49827
rect 25329 49793 25363 49827
rect 25363 49793 25372 49827
rect 25320 49784 25372 49793
rect 8852 49716 8904 49768
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 11980 49376 12032 49428
rect 1492 49240 1544 49292
rect 10692 49172 10744 49224
rect 25320 49215 25372 49224
rect 25320 49181 25329 49215
rect 25329 49181 25363 49215
rect 25363 49181 25372 49215
rect 25320 49172 25372 49181
rect 10784 49036 10836 49088
rect 18328 49036 18380 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 12808 48832 12860 48884
rect 12532 48696 12584 48748
rect 25504 48535 25556 48544
rect 25504 48501 25513 48535
rect 25513 48501 25547 48535
rect 25547 48501 25556 48535
rect 25504 48492 25556 48501
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 17316 48220 17368 48272
rect 19432 48220 19484 48272
rect 25320 48127 25372 48136
rect 25320 48093 25329 48127
rect 25329 48093 25363 48127
rect 25363 48093 25372 48127
rect 25320 48084 25372 48093
rect 1308 48016 1360 48068
rect 4068 47948 4120 48000
rect 7564 47948 7616 48000
rect 11336 47948 11388 48000
rect 20260 47948 20312 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 9128 47787 9180 47796
rect 9128 47753 9137 47787
rect 9137 47753 9171 47787
rect 9171 47753 9180 47787
rect 9128 47744 9180 47753
rect 17224 47787 17276 47796
rect 17224 47753 17233 47787
rect 17233 47753 17267 47787
rect 17267 47753 17276 47787
rect 17224 47744 17276 47753
rect 17316 47787 17368 47796
rect 17316 47753 17325 47787
rect 17325 47753 17359 47787
rect 17359 47753 17368 47787
rect 17316 47744 17368 47753
rect 18420 47787 18472 47796
rect 18420 47753 18429 47787
rect 18429 47753 18463 47787
rect 18463 47753 18472 47787
rect 18420 47744 18472 47753
rect 18512 47787 18564 47796
rect 18512 47753 18521 47787
rect 18521 47753 18555 47787
rect 18555 47753 18564 47787
rect 18512 47744 18564 47753
rect 11428 47608 11480 47660
rect 24400 47608 24452 47660
rect 16304 47472 16356 47524
rect 18420 47540 18472 47592
rect 25504 47540 25556 47592
rect 16580 47404 16632 47456
rect 17500 47404 17552 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 9864 47243 9916 47252
rect 9864 47209 9873 47243
rect 9873 47209 9907 47243
rect 9907 47209 9916 47243
rect 9864 47200 9916 47209
rect 18420 47200 18472 47252
rect 18512 47132 18564 47184
rect 20352 47200 20404 47252
rect 21640 47243 21692 47252
rect 21640 47209 21649 47243
rect 21649 47209 21683 47243
rect 21683 47209 21692 47243
rect 21640 47200 21692 47209
rect 16672 47064 16724 47116
rect 16948 47064 17000 47116
rect 17316 47064 17368 47116
rect 18604 47107 18656 47116
rect 18604 47073 18613 47107
rect 18613 47073 18647 47107
rect 18647 47073 18656 47107
rect 18604 47064 18656 47073
rect 21824 47132 21876 47184
rect 19340 47064 19392 47116
rect 21640 46996 21692 47048
rect 22652 46996 22704 47048
rect 9036 46928 9088 46980
rect 10508 46971 10560 46980
rect 10508 46937 10517 46971
rect 10517 46937 10551 46971
rect 10551 46937 10560 46971
rect 10508 46928 10560 46937
rect 10048 46860 10100 46912
rect 12624 46928 12676 46980
rect 13084 46928 13136 46980
rect 16396 46928 16448 46980
rect 12164 46860 12216 46912
rect 17592 46860 17644 46912
rect 22008 46903 22060 46912
rect 22008 46869 22017 46903
rect 22017 46869 22051 46903
rect 22051 46869 22060 46903
rect 22008 46860 22060 46869
rect 22652 46860 22704 46912
rect 24768 46928 24820 46980
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 7472 46656 7524 46708
rect 10876 46699 10928 46708
rect 10876 46665 10885 46699
rect 10885 46665 10919 46699
rect 10919 46665 10928 46699
rect 10876 46656 10928 46665
rect 14188 46656 14240 46708
rect 18420 46656 18472 46708
rect 18972 46656 19024 46708
rect 22560 46656 22612 46708
rect 13084 46588 13136 46640
rect 15108 46588 15160 46640
rect 16396 46588 16448 46640
rect 17592 46588 17644 46640
rect 20904 46588 20956 46640
rect 22744 46699 22796 46708
rect 22744 46665 22753 46699
rect 22753 46665 22787 46699
rect 22787 46665 22796 46699
rect 22744 46656 22796 46665
rect 7564 46520 7616 46572
rect 11060 46563 11112 46572
rect 11060 46529 11069 46563
rect 11069 46529 11103 46563
rect 11103 46529 11112 46563
rect 11060 46520 11112 46529
rect 24216 46520 24268 46572
rect 11888 46452 11940 46504
rect 13360 46452 13412 46504
rect 13728 46316 13780 46368
rect 16304 46359 16356 46368
rect 16304 46325 16313 46359
rect 16313 46325 16347 46359
rect 16347 46325 16356 46359
rect 16304 46316 16356 46325
rect 16856 46495 16908 46504
rect 16856 46461 16865 46495
rect 16865 46461 16899 46495
rect 16899 46461 16908 46495
rect 16856 46452 16908 46461
rect 18604 46452 18656 46504
rect 17224 46316 17276 46368
rect 19340 46495 19392 46504
rect 19340 46461 19349 46495
rect 19349 46461 19383 46495
rect 19383 46461 19392 46495
rect 19340 46452 19392 46461
rect 22192 46452 22244 46504
rect 24492 46495 24544 46504
rect 24492 46461 24501 46495
rect 24501 46461 24535 46495
rect 24535 46461 24544 46495
rect 24492 46452 24544 46461
rect 19432 46316 19484 46368
rect 22744 46316 22796 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 5908 46112 5960 46164
rect 9220 46112 9272 46164
rect 10692 46155 10744 46164
rect 10692 46121 10701 46155
rect 10701 46121 10735 46155
rect 10735 46121 10744 46155
rect 10692 46112 10744 46121
rect 17592 46112 17644 46164
rect 19616 46112 19668 46164
rect 24492 46112 24544 46164
rect 25504 46112 25556 46164
rect 7656 46044 7708 46096
rect 9496 45976 9548 46028
rect 11888 46019 11940 46028
rect 11888 45985 11897 46019
rect 11897 45985 11931 46019
rect 11931 45985 11940 46019
rect 11888 45976 11940 45985
rect 12164 46019 12216 46028
rect 12164 45985 12173 46019
rect 12173 45985 12207 46019
rect 12207 45985 12216 46019
rect 12164 45976 12216 45985
rect 12624 45976 12676 46028
rect 14004 45976 14056 46028
rect 20168 46019 20220 46028
rect 20168 45985 20177 46019
rect 20177 45985 20211 46019
rect 20211 45985 20220 46019
rect 20168 45976 20220 45985
rect 20444 45976 20496 46028
rect 21364 46019 21416 46028
rect 21364 45985 21373 46019
rect 21373 45985 21407 46019
rect 21407 45985 21416 46019
rect 21364 45976 21416 45985
rect 21732 45976 21784 46028
rect 1308 45908 1360 45960
rect 7196 45908 7248 45960
rect 6920 45840 6972 45892
rect 11796 45908 11848 45960
rect 19616 45908 19668 45960
rect 20076 45951 20128 45960
rect 20076 45917 20085 45951
rect 20085 45917 20119 45951
rect 20119 45917 20128 45951
rect 20076 45908 20128 45917
rect 21088 45908 21140 45960
rect 21916 45951 21968 45960
rect 21916 45917 21925 45951
rect 21925 45917 21959 45951
rect 21959 45917 21968 45951
rect 21916 45908 21968 45917
rect 11152 45815 11204 45824
rect 11152 45781 11161 45815
rect 11161 45781 11195 45815
rect 11195 45781 11204 45815
rect 11152 45772 11204 45781
rect 12624 45840 12676 45892
rect 14740 45840 14792 45892
rect 13636 45815 13688 45824
rect 13636 45781 13645 45815
rect 13645 45781 13679 45815
rect 13679 45781 13688 45815
rect 13636 45772 13688 45781
rect 16396 45815 16448 45824
rect 16396 45781 16405 45815
rect 16405 45781 16439 45815
rect 16439 45781 16448 45815
rect 16396 45772 16448 45781
rect 19892 45772 19944 45824
rect 20720 45772 20772 45824
rect 24032 45908 24084 45960
rect 24860 45772 24912 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 1308 45568 1360 45620
rect 19340 45568 19392 45620
rect 8852 45543 8904 45552
rect 8852 45509 8861 45543
rect 8861 45509 8895 45543
rect 8895 45509 8904 45543
rect 8852 45500 8904 45509
rect 9772 45500 9824 45552
rect 10048 45500 10100 45552
rect 14004 45500 14056 45552
rect 15108 45500 15160 45552
rect 21732 45500 21784 45552
rect 9220 45475 9272 45484
rect 9220 45441 9229 45475
rect 9229 45441 9263 45475
rect 9263 45441 9272 45475
rect 9220 45432 9272 45441
rect 9864 45364 9916 45416
rect 10508 45296 10560 45348
rect 12256 45296 12308 45348
rect 10048 45228 10100 45280
rect 12440 45228 12492 45280
rect 16304 45364 16356 45416
rect 18328 45364 18380 45416
rect 20076 45364 20128 45416
rect 15844 45296 15896 45348
rect 16396 45339 16448 45348
rect 16396 45305 16405 45339
rect 16405 45305 16439 45339
rect 16439 45305 16448 45339
rect 16396 45296 16448 45305
rect 14832 45228 14884 45280
rect 16120 45271 16172 45280
rect 16120 45237 16129 45271
rect 16129 45237 16163 45271
rect 16163 45237 16172 45271
rect 16120 45228 16172 45237
rect 18880 45228 18932 45280
rect 20904 45228 20956 45280
rect 23388 45296 23440 45348
rect 22284 45228 22336 45280
rect 24492 45407 24544 45416
rect 24492 45373 24501 45407
rect 24501 45373 24535 45407
rect 24535 45373 24544 45407
rect 24492 45364 24544 45373
rect 24676 45364 24728 45416
rect 24308 45228 24360 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 7288 45024 7340 45076
rect 11244 45024 11296 45076
rect 12072 45024 12124 45076
rect 12532 45024 12584 45076
rect 16396 45024 16448 45076
rect 4712 44956 4764 45008
rect 12624 44888 12676 44940
rect 13728 44888 13780 44940
rect 13452 44820 13504 44872
rect 14832 44820 14884 44872
rect 16856 44888 16908 44940
rect 21640 44931 21692 44940
rect 21640 44897 21649 44931
rect 21649 44897 21683 44931
rect 21683 44897 21692 44931
rect 21640 44888 21692 44897
rect 16764 44820 16816 44872
rect 16948 44820 17000 44872
rect 19524 44863 19576 44872
rect 19524 44829 19533 44863
rect 19533 44829 19567 44863
rect 19567 44829 19576 44863
rect 19524 44820 19576 44829
rect 20904 44820 20956 44872
rect 22284 44863 22336 44872
rect 22284 44829 22293 44863
rect 22293 44829 22327 44863
rect 22327 44829 22336 44863
rect 22284 44820 22336 44829
rect 6644 44684 6696 44736
rect 7288 44684 7340 44736
rect 8668 44684 8720 44736
rect 9772 44727 9824 44736
rect 9772 44693 9781 44727
rect 9781 44693 9815 44727
rect 9815 44693 9824 44727
rect 9772 44684 9824 44693
rect 12440 44752 12492 44804
rect 15660 44752 15712 44804
rect 15844 44752 15896 44804
rect 19800 44795 19852 44804
rect 19800 44761 19809 44795
rect 19809 44761 19843 44795
rect 19843 44761 19852 44795
rect 19800 44752 19852 44761
rect 22560 44795 22612 44804
rect 22560 44761 22569 44795
rect 22569 44761 22603 44795
rect 22603 44761 22612 44795
rect 22560 44752 22612 44761
rect 12532 44684 12584 44736
rect 15200 44684 15252 44736
rect 17224 44684 17276 44736
rect 19984 44684 20036 44736
rect 23388 44684 23440 44736
rect 24308 44684 24360 44736
rect 24492 44684 24544 44736
rect 25504 44727 25556 44736
rect 25504 44693 25513 44727
rect 25513 44693 25547 44727
rect 25547 44693 25556 44727
rect 25504 44684 25556 44693
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 5816 44523 5868 44532
rect 5816 44489 5825 44523
rect 5825 44489 5859 44523
rect 5859 44489 5868 44523
rect 5816 44480 5868 44489
rect 6736 44523 6788 44532
rect 6736 44489 6745 44523
rect 6745 44489 6779 44523
rect 6779 44489 6788 44523
rect 6736 44480 6788 44489
rect 7380 44480 7432 44532
rect 7840 44480 7892 44532
rect 9680 44480 9732 44532
rect 11152 44480 11204 44532
rect 16396 44480 16448 44532
rect 18880 44523 18932 44532
rect 7104 44412 7156 44464
rect 12348 44412 12400 44464
rect 5264 44344 5316 44396
rect 6736 44344 6788 44396
rect 7380 44387 7432 44396
rect 7380 44353 7389 44387
rect 7389 44353 7423 44387
rect 7423 44353 7432 44387
rect 7380 44344 7432 44353
rect 7472 44344 7524 44396
rect 8944 44387 8996 44396
rect 8944 44353 8953 44387
rect 8953 44353 8987 44387
rect 8987 44353 8996 44387
rect 13360 44412 13412 44464
rect 14004 44412 14056 44464
rect 15108 44412 15160 44464
rect 15844 44412 15896 44464
rect 18880 44489 18889 44523
rect 18889 44489 18923 44523
rect 18923 44489 18932 44523
rect 18880 44480 18932 44489
rect 19800 44480 19852 44532
rect 20444 44480 20496 44532
rect 21640 44523 21692 44532
rect 21640 44489 21649 44523
rect 21649 44489 21683 44523
rect 21683 44489 21692 44523
rect 21640 44480 21692 44489
rect 22560 44480 22612 44532
rect 24308 44412 24360 44464
rect 8944 44344 8996 44353
rect 25320 44344 25372 44396
rect 11704 44276 11756 44328
rect 11612 44251 11664 44260
rect 11612 44217 11621 44251
rect 11621 44217 11655 44251
rect 11655 44217 11664 44251
rect 11612 44208 11664 44217
rect 12256 44208 12308 44260
rect 14188 44276 14240 44328
rect 16856 44319 16908 44328
rect 16856 44285 16865 44319
rect 16865 44285 16899 44319
rect 16899 44285 16908 44319
rect 16856 44276 16908 44285
rect 18972 44276 19024 44328
rect 19524 44319 19576 44328
rect 19524 44285 19533 44319
rect 19533 44285 19567 44319
rect 19567 44285 19576 44319
rect 19524 44276 19576 44285
rect 13636 44140 13688 44192
rect 16488 44140 16540 44192
rect 18328 44140 18380 44192
rect 18604 44183 18656 44192
rect 18604 44149 18613 44183
rect 18613 44149 18647 44183
rect 18647 44149 18656 44183
rect 18604 44140 18656 44149
rect 18788 44140 18840 44192
rect 20812 44276 20864 44328
rect 22284 44319 22336 44328
rect 22284 44285 22293 44319
rect 22293 44285 22327 44319
rect 22327 44285 22336 44319
rect 22284 44276 22336 44285
rect 22652 44276 22704 44328
rect 24768 44319 24820 44328
rect 24768 44285 24777 44319
rect 24777 44285 24811 44319
rect 24811 44285 24820 44319
rect 24768 44276 24820 44285
rect 23296 44140 23348 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 9404 43936 9456 43988
rect 11336 43936 11388 43988
rect 23296 43936 23348 43988
rect 23480 43936 23532 43988
rect 7012 43868 7064 43920
rect 9404 43800 9456 43852
rect 22468 43843 22520 43852
rect 22468 43809 22477 43843
rect 22477 43809 22511 43843
rect 22511 43809 22520 43843
rect 22468 43800 22520 43809
rect 23296 43800 23348 43852
rect 8484 43732 8536 43784
rect 1216 43596 1268 43648
rect 7104 43596 7156 43648
rect 10048 43664 10100 43716
rect 15476 43732 15528 43784
rect 10968 43596 11020 43648
rect 12072 43639 12124 43648
rect 12072 43605 12081 43639
rect 12081 43605 12115 43639
rect 12115 43605 12124 43639
rect 12072 43596 12124 43605
rect 17408 43596 17460 43648
rect 20260 43596 20312 43648
rect 21916 43596 21968 43648
rect 22468 43596 22520 43648
rect 22836 43596 22888 43648
rect 24308 43596 24360 43648
rect 25320 43639 25372 43648
rect 25320 43605 25329 43639
rect 25329 43605 25363 43639
rect 25363 43605 25372 43639
rect 25320 43596 25372 43605
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 7748 43435 7800 43444
rect 7748 43401 7757 43435
rect 7757 43401 7791 43435
rect 7791 43401 7800 43435
rect 7748 43392 7800 43401
rect 8576 43392 8628 43444
rect 9588 43392 9640 43444
rect 10416 43392 10468 43444
rect 15016 43435 15068 43444
rect 15016 43401 15025 43435
rect 15025 43401 15059 43435
rect 15059 43401 15068 43435
rect 15016 43392 15068 43401
rect 17408 43435 17460 43444
rect 17408 43401 17417 43435
rect 17417 43401 17451 43435
rect 17451 43401 17460 43435
rect 17408 43392 17460 43401
rect 17500 43435 17552 43444
rect 17500 43401 17509 43435
rect 17509 43401 17543 43435
rect 17543 43401 17552 43435
rect 17500 43392 17552 43401
rect 20076 43435 20128 43444
rect 20076 43401 20085 43435
rect 20085 43401 20119 43435
rect 20119 43401 20128 43435
rect 20076 43392 20128 43401
rect 4620 43324 4672 43376
rect 10048 43324 10100 43376
rect 12624 43367 12676 43376
rect 12624 43333 12633 43367
rect 12633 43333 12667 43367
rect 12667 43333 12676 43367
rect 12624 43324 12676 43333
rect 14004 43324 14056 43376
rect 21364 43392 21416 43444
rect 21640 43392 21692 43444
rect 22376 43392 22428 43444
rect 1216 43256 1268 43308
rect 7656 43256 7708 43308
rect 8392 43256 8444 43308
rect 9496 43256 9548 43308
rect 10324 43256 10376 43308
rect 12348 43299 12400 43308
rect 12348 43265 12357 43299
rect 12357 43265 12391 43299
rect 12391 43265 12400 43299
rect 12348 43256 12400 43265
rect 8852 43188 8904 43240
rect 11704 43120 11756 43172
rect 14924 43120 14976 43172
rect 2228 43095 2280 43104
rect 2228 43061 2237 43095
rect 2237 43061 2271 43095
rect 2271 43061 2280 43095
rect 2228 43052 2280 43061
rect 14004 43052 14056 43104
rect 14188 43052 14240 43104
rect 24308 43324 24360 43376
rect 21640 43256 21692 43308
rect 15660 43188 15712 43240
rect 17316 43188 17368 43240
rect 18328 43231 18380 43240
rect 18328 43197 18337 43231
rect 18337 43197 18371 43231
rect 18371 43197 18380 43231
rect 18328 43188 18380 43197
rect 19984 43188 20036 43240
rect 22652 43231 22704 43240
rect 22652 43197 22661 43231
rect 22661 43197 22695 43231
rect 22695 43197 22704 43231
rect 22652 43188 22704 43197
rect 23480 43188 23532 43240
rect 23848 43231 23900 43240
rect 23848 43197 23857 43231
rect 23857 43197 23891 43231
rect 23891 43197 23900 43231
rect 23848 43188 23900 43197
rect 18144 43120 18196 43172
rect 15568 43052 15620 43104
rect 15844 43052 15896 43104
rect 16672 43095 16724 43104
rect 16672 43061 16681 43095
rect 16681 43061 16715 43095
rect 16715 43061 16724 43095
rect 16672 43052 16724 43061
rect 17040 43095 17092 43104
rect 17040 43061 17049 43095
rect 17049 43061 17083 43095
rect 17083 43061 17092 43095
rect 17040 43052 17092 43061
rect 19248 43052 19300 43104
rect 21640 43095 21692 43104
rect 21640 43061 21649 43095
rect 21649 43061 21683 43095
rect 21683 43061 21692 43095
rect 21640 43052 21692 43061
rect 24952 43052 25004 43104
rect 25228 43052 25280 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 8576 42891 8628 42900
rect 8576 42857 8585 42891
rect 8585 42857 8619 42891
rect 8619 42857 8628 42891
rect 8576 42848 8628 42857
rect 4896 42712 4948 42764
rect 8576 42712 8628 42764
rect 8852 42848 8904 42900
rect 9312 42848 9364 42900
rect 9496 42848 9548 42900
rect 12164 42848 12216 42900
rect 13912 42848 13964 42900
rect 15568 42848 15620 42900
rect 15844 42848 15896 42900
rect 16672 42848 16724 42900
rect 20352 42848 20404 42900
rect 21732 42848 21784 42900
rect 9220 42712 9272 42764
rect 9404 42712 9456 42764
rect 12348 42712 12400 42764
rect 14832 42755 14884 42764
rect 14832 42721 14841 42755
rect 14841 42721 14875 42755
rect 14875 42721 14884 42755
rect 14832 42712 14884 42721
rect 18144 42755 18196 42764
rect 18144 42721 18153 42755
rect 18153 42721 18187 42755
rect 18187 42721 18196 42755
rect 18144 42712 18196 42721
rect 18420 42755 18472 42764
rect 18420 42721 18429 42755
rect 18429 42721 18463 42755
rect 18463 42721 18472 42755
rect 18420 42712 18472 42721
rect 2228 42644 2280 42696
rect 12164 42644 12216 42696
rect 12440 42644 12492 42696
rect 14372 42644 14424 42696
rect 21364 42644 21416 42696
rect 22008 42712 22060 42764
rect 22560 42712 22612 42764
rect 24308 42712 24360 42764
rect 22836 42644 22888 42696
rect 3976 42576 4028 42628
rect 4804 42619 4856 42628
rect 4804 42585 4813 42619
rect 4813 42585 4847 42619
rect 4847 42585 4856 42619
rect 4804 42576 4856 42585
rect 7564 42576 7616 42628
rect 9680 42576 9732 42628
rect 8392 42508 8444 42560
rect 8852 42508 8904 42560
rect 10324 42551 10376 42560
rect 10324 42517 10333 42551
rect 10333 42517 10367 42551
rect 10367 42517 10376 42551
rect 10324 42508 10376 42517
rect 10876 42508 10928 42560
rect 12440 42508 12492 42560
rect 15568 42576 15620 42628
rect 16396 42576 16448 42628
rect 16672 42508 16724 42560
rect 21180 42576 21232 42628
rect 23664 42644 23716 42696
rect 23756 42644 23808 42696
rect 24860 42644 24912 42696
rect 19340 42508 19392 42560
rect 20536 42508 20588 42560
rect 22100 42508 22152 42560
rect 24860 42508 24912 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 4160 42304 4212 42356
rect 5080 42347 5132 42356
rect 5080 42313 5089 42347
rect 5089 42313 5123 42347
rect 5123 42313 5132 42347
rect 5080 42304 5132 42313
rect 5448 42304 5500 42356
rect 8116 42304 8168 42356
rect 9220 42304 9272 42356
rect 9680 42347 9732 42356
rect 9680 42313 9689 42347
rect 9689 42313 9723 42347
rect 9723 42313 9732 42347
rect 9680 42304 9732 42313
rect 11428 42304 11480 42356
rect 13452 42304 13504 42356
rect 15200 42304 15252 42356
rect 19800 42304 19852 42356
rect 20168 42304 20220 42356
rect 4252 42211 4304 42220
rect 4252 42177 4261 42211
rect 4261 42177 4295 42211
rect 4295 42177 4304 42211
rect 4252 42168 4304 42177
rect 7012 42168 7064 42220
rect 15568 42236 15620 42288
rect 17868 42236 17920 42288
rect 20720 42347 20772 42356
rect 20720 42313 20729 42347
rect 20729 42313 20763 42347
rect 20763 42313 20772 42347
rect 20720 42304 20772 42313
rect 21364 42347 21416 42356
rect 21364 42313 21373 42347
rect 21373 42313 21407 42347
rect 21407 42313 21416 42347
rect 21364 42304 21416 42313
rect 23296 42304 23348 42356
rect 21088 42236 21140 42288
rect 24308 42236 24360 42288
rect 8852 42168 8904 42220
rect 9128 42168 9180 42220
rect 7748 42143 7800 42152
rect 7748 42109 7757 42143
rect 7757 42109 7791 42143
rect 7791 42109 7800 42143
rect 11152 42168 11204 42220
rect 7748 42100 7800 42109
rect 10140 42143 10192 42152
rect 10140 42109 10149 42143
rect 10149 42109 10183 42143
rect 10183 42109 10192 42143
rect 10140 42100 10192 42109
rect 12440 42143 12492 42152
rect 12440 42109 12449 42143
rect 12449 42109 12483 42143
rect 12483 42109 12492 42143
rect 12440 42100 12492 42109
rect 13360 42032 13412 42084
rect 14280 42100 14332 42152
rect 6092 41964 6144 42016
rect 7012 41964 7064 42016
rect 9588 41964 9640 42016
rect 10508 41964 10560 42016
rect 15108 41964 15160 42016
rect 16488 42032 16540 42084
rect 19524 42168 19576 42220
rect 19248 42100 19300 42152
rect 19708 42100 19760 42152
rect 20536 42100 20588 42152
rect 22836 42143 22888 42152
rect 22836 42109 22845 42143
rect 22845 42109 22879 42143
rect 22879 42109 22888 42143
rect 23480 42143 23532 42152
rect 22836 42100 22888 42109
rect 23480 42109 23489 42143
rect 23489 42109 23523 42143
rect 23523 42109 23532 42143
rect 23480 42100 23532 42109
rect 25228 42100 25280 42152
rect 20720 41964 20772 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 5172 41803 5224 41812
rect 5172 41769 5181 41803
rect 5181 41769 5215 41803
rect 5215 41769 5224 41803
rect 5172 41760 5224 41769
rect 7748 41760 7800 41812
rect 7840 41760 7892 41812
rect 8116 41803 8168 41812
rect 8116 41769 8125 41803
rect 8125 41769 8159 41803
rect 8159 41769 8168 41803
rect 8116 41760 8168 41769
rect 11060 41760 11112 41812
rect 20812 41760 20864 41812
rect 21272 41760 21324 41812
rect 21732 41760 21784 41812
rect 25872 41760 25924 41812
rect 6184 41624 6236 41676
rect 8300 41692 8352 41744
rect 8760 41692 8812 41744
rect 9680 41692 9732 41744
rect 10876 41692 10928 41744
rect 9220 41624 9272 41676
rect 10600 41624 10652 41676
rect 10784 41624 10836 41676
rect 12348 41624 12400 41676
rect 12808 41624 12860 41676
rect 13636 41624 13688 41676
rect 13912 41624 13964 41676
rect 16120 41624 16172 41676
rect 10508 41556 10560 41608
rect 1400 41463 1452 41472
rect 1400 41429 1409 41463
rect 1409 41429 1443 41463
rect 1443 41429 1452 41463
rect 1400 41420 1452 41429
rect 5724 41420 5776 41472
rect 7748 41488 7800 41540
rect 9128 41488 9180 41540
rect 16580 41556 16632 41608
rect 7564 41420 7616 41472
rect 8576 41420 8628 41472
rect 9312 41420 9364 41472
rect 10784 41420 10836 41472
rect 10968 41420 11020 41472
rect 11060 41463 11112 41472
rect 11060 41429 11069 41463
rect 11069 41429 11103 41463
rect 11103 41429 11112 41463
rect 11060 41420 11112 41429
rect 12348 41420 12400 41472
rect 16212 41463 16264 41472
rect 16212 41429 16221 41463
rect 16221 41429 16255 41463
rect 16255 41429 16264 41463
rect 16212 41420 16264 41429
rect 18512 41624 18564 41676
rect 18972 41624 19024 41676
rect 19248 41624 19300 41676
rect 25044 41692 25096 41744
rect 22560 41624 22612 41676
rect 22744 41624 22796 41676
rect 23480 41624 23532 41676
rect 23848 41624 23900 41676
rect 23756 41556 23808 41608
rect 25320 41599 25372 41608
rect 25320 41565 25329 41599
rect 25329 41565 25363 41599
rect 25363 41565 25372 41599
rect 25320 41556 25372 41565
rect 19708 41531 19760 41540
rect 19708 41497 19717 41531
rect 19717 41497 19751 41531
rect 19751 41497 19760 41531
rect 19708 41488 19760 41497
rect 21364 41488 21416 41540
rect 21548 41488 21600 41540
rect 22284 41488 22336 41540
rect 18420 41420 18472 41472
rect 19156 41420 19208 41472
rect 21640 41463 21692 41472
rect 21640 41429 21649 41463
rect 21649 41429 21683 41463
rect 21683 41429 21692 41463
rect 21640 41420 21692 41429
rect 22008 41463 22060 41472
rect 22008 41429 22017 41463
rect 22017 41429 22051 41463
rect 22051 41429 22060 41463
rect 22008 41420 22060 41429
rect 23848 41420 23900 41472
rect 24308 41420 24360 41472
rect 24860 41463 24912 41472
rect 24860 41429 24869 41463
rect 24869 41429 24903 41463
rect 24903 41429 24912 41463
rect 24860 41420 24912 41429
rect 25136 41463 25188 41472
rect 25136 41429 25145 41463
rect 25145 41429 25179 41463
rect 25179 41429 25188 41463
rect 25136 41420 25188 41429
rect 25320 41420 25372 41472
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 1952 41216 2004 41268
rect 6184 41216 6236 41268
rect 7840 41216 7892 41268
rect 1308 41080 1360 41132
rect 4620 41080 4672 41132
rect 9404 41216 9456 41268
rect 9128 41148 9180 41200
rect 10048 41216 10100 41268
rect 11520 41216 11572 41268
rect 11704 41259 11756 41268
rect 11704 41225 11713 41259
rect 11713 41225 11747 41259
rect 11747 41225 11756 41259
rect 11704 41216 11756 41225
rect 14924 41216 14976 41268
rect 15844 41216 15896 41268
rect 10508 41080 10560 41132
rect 13636 41123 13688 41132
rect 13636 41089 13645 41123
rect 13645 41089 13679 41123
rect 13679 41089 13688 41123
rect 13636 41080 13688 41089
rect 15016 41080 15068 41132
rect 19248 41216 19300 41268
rect 19892 41259 19944 41268
rect 19892 41225 19901 41259
rect 19901 41225 19935 41259
rect 19935 41225 19944 41259
rect 19892 41216 19944 41225
rect 22008 41259 22060 41268
rect 22008 41225 22017 41259
rect 22017 41225 22051 41259
rect 22051 41225 22060 41259
rect 22008 41216 22060 41225
rect 23480 41216 23532 41268
rect 18880 41191 18932 41200
rect 18880 41157 18889 41191
rect 18889 41157 18923 41191
rect 18923 41157 18932 41191
rect 18880 41148 18932 41157
rect 24492 41148 24544 41200
rect 20444 41080 20496 41132
rect 20904 41080 20956 41132
rect 25320 41123 25372 41132
rect 25320 41089 25329 41123
rect 25329 41089 25363 41123
rect 25363 41089 25372 41123
rect 25320 41080 25372 41089
rect 10232 41012 10284 41064
rect 12256 41055 12308 41064
rect 12256 41021 12265 41055
rect 12265 41021 12299 41055
rect 12299 41021 12308 41055
rect 12256 41012 12308 41021
rect 13912 41055 13964 41064
rect 13912 41021 13921 41055
rect 13921 41021 13955 41055
rect 13955 41021 13964 41055
rect 13912 41012 13964 41021
rect 16672 41012 16724 41064
rect 15384 40987 15436 40996
rect 15384 40953 15393 40987
rect 15393 40953 15427 40987
rect 15427 40953 15436 40987
rect 15384 40944 15436 40953
rect 16396 40944 16448 40996
rect 19984 41055 20036 41064
rect 19984 41021 19993 41055
rect 19993 41021 20027 41055
rect 20027 41021 20036 41055
rect 19984 41012 20036 41021
rect 20996 41012 21048 41064
rect 22468 41012 22520 41064
rect 22652 41012 22704 41064
rect 22836 41012 22888 41064
rect 22192 40944 22244 40996
rect 24860 41012 24912 41064
rect 1768 40876 1820 40928
rect 8484 40876 8536 40928
rect 9036 40876 9088 40928
rect 10324 40876 10376 40928
rect 10692 40919 10744 40928
rect 10692 40885 10701 40919
rect 10701 40885 10735 40919
rect 10735 40885 10744 40919
rect 10692 40876 10744 40885
rect 18328 40876 18380 40928
rect 19156 40919 19208 40928
rect 19156 40885 19165 40919
rect 19165 40885 19199 40919
rect 19199 40885 19208 40919
rect 19156 40876 19208 40885
rect 19432 40919 19484 40928
rect 19432 40885 19441 40919
rect 19441 40885 19475 40919
rect 19475 40885 19484 40919
rect 19432 40876 19484 40885
rect 20812 40876 20864 40928
rect 20904 40876 20956 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 7564 40672 7616 40724
rect 8484 40715 8536 40724
rect 8484 40681 8493 40715
rect 8493 40681 8527 40715
rect 8527 40681 8536 40715
rect 8484 40672 8536 40681
rect 9588 40672 9640 40724
rect 10600 40715 10652 40724
rect 10600 40681 10609 40715
rect 10609 40681 10643 40715
rect 10643 40681 10652 40715
rect 10600 40672 10652 40681
rect 17684 40672 17736 40724
rect 19984 40672 20036 40724
rect 21180 40672 21232 40724
rect 6552 40536 6604 40588
rect 9404 40536 9456 40588
rect 14648 40604 14700 40656
rect 18696 40604 18748 40656
rect 13636 40536 13688 40588
rect 13820 40536 13872 40588
rect 14004 40536 14056 40588
rect 16948 40536 17000 40588
rect 17040 40536 17092 40588
rect 17224 40579 17276 40588
rect 17224 40545 17233 40579
rect 17233 40545 17267 40579
rect 17267 40545 17276 40579
rect 17224 40536 17276 40545
rect 1768 40511 1820 40520
rect 1768 40477 1777 40511
rect 1777 40477 1811 40511
rect 1811 40477 1820 40511
rect 1768 40468 1820 40477
rect 6184 40511 6236 40520
rect 6184 40477 6193 40511
rect 6193 40477 6227 40511
rect 6227 40477 6236 40511
rect 6184 40468 6236 40477
rect 1860 40332 1912 40384
rect 7288 40332 7340 40384
rect 9220 40468 9272 40520
rect 11888 40468 11940 40520
rect 11980 40468 12032 40520
rect 9496 40400 9548 40452
rect 8300 40375 8352 40384
rect 8300 40341 8309 40375
rect 8309 40341 8343 40375
rect 8343 40341 8352 40375
rect 8300 40332 8352 40341
rect 9128 40332 9180 40384
rect 9220 40375 9272 40384
rect 9220 40341 9229 40375
rect 9229 40341 9263 40375
rect 9263 40341 9272 40375
rect 9220 40332 9272 40341
rect 9588 40375 9640 40384
rect 9588 40341 9597 40375
rect 9597 40341 9631 40375
rect 9631 40341 9640 40375
rect 9588 40332 9640 40341
rect 12256 40400 12308 40452
rect 12716 40468 12768 40520
rect 16856 40468 16908 40520
rect 19340 40468 19392 40520
rect 19984 40468 20036 40520
rect 21180 40468 21232 40520
rect 22744 40672 22796 40724
rect 25780 40672 25832 40724
rect 21548 40579 21600 40588
rect 21548 40545 21557 40579
rect 21557 40545 21591 40579
rect 21591 40545 21600 40579
rect 21548 40536 21600 40545
rect 21732 40536 21784 40588
rect 22100 40536 22152 40588
rect 23388 40536 23440 40588
rect 21640 40468 21692 40520
rect 23020 40468 23072 40520
rect 24400 40468 24452 40520
rect 24768 40468 24820 40520
rect 15844 40400 15896 40452
rect 19156 40400 19208 40452
rect 12164 40375 12216 40384
rect 12164 40341 12173 40375
rect 12173 40341 12207 40375
rect 12207 40341 12216 40375
rect 12164 40332 12216 40341
rect 12624 40375 12676 40384
rect 12624 40341 12633 40375
rect 12633 40341 12667 40375
rect 12667 40341 12676 40375
rect 12624 40332 12676 40341
rect 15200 40375 15252 40384
rect 15200 40341 15209 40375
rect 15209 40341 15243 40375
rect 15243 40341 15252 40375
rect 15200 40332 15252 40341
rect 16304 40375 16356 40384
rect 16304 40341 16313 40375
rect 16313 40341 16347 40375
rect 16347 40341 16356 40375
rect 16304 40332 16356 40341
rect 17500 40332 17552 40384
rect 20444 40332 20496 40384
rect 21548 40400 21600 40452
rect 22376 40400 22428 40452
rect 23756 40400 23808 40452
rect 21732 40332 21784 40384
rect 23388 40332 23440 40384
rect 24216 40375 24268 40384
rect 24216 40341 24225 40375
rect 24225 40341 24259 40375
rect 24259 40341 24268 40375
rect 24216 40332 24268 40341
rect 24492 40375 24544 40384
rect 24492 40341 24501 40375
rect 24501 40341 24535 40375
rect 24535 40341 24544 40375
rect 24492 40332 24544 40341
rect 24584 40332 24636 40384
rect 25320 40332 25372 40384
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 7196 40128 7248 40180
rect 9128 40128 9180 40180
rect 9404 40128 9456 40180
rect 8760 40060 8812 40112
rect 11520 40171 11572 40180
rect 11520 40137 11529 40171
rect 11529 40137 11563 40171
rect 11563 40137 11572 40171
rect 11520 40128 11572 40137
rect 12256 40171 12308 40180
rect 12256 40137 12265 40171
rect 12265 40137 12299 40171
rect 12299 40137 12308 40171
rect 12256 40128 12308 40137
rect 14648 40128 14700 40180
rect 15016 40171 15068 40180
rect 15016 40137 15025 40171
rect 15025 40137 15059 40171
rect 15059 40137 15068 40171
rect 15016 40128 15068 40137
rect 15568 40171 15620 40180
rect 15568 40137 15577 40171
rect 15577 40137 15611 40171
rect 15611 40137 15620 40171
rect 15568 40128 15620 40137
rect 16304 40128 16356 40180
rect 22100 40128 22152 40180
rect 22652 40128 22704 40180
rect 14556 40060 14608 40112
rect 7932 39992 7984 40044
rect 12440 39992 12492 40044
rect 12808 39992 12860 40044
rect 18604 40103 18656 40112
rect 18604 40069 18613 40103
rect 18613 40069 18647 40103
rect 18647 40069 18656 40103
rect 18604 40060 18656 40069
rect 16304 39992 16356 40044
rect 7840 39967 7892 39976
rect 7840 39933 7849 39967
rect 7849 39933 7883 39967
rect 7883 39933 7892 39967
rect 7840 39924 7892 39933
rect 10324 39924 10376 39976
rect 10968 39967 11020 39976
rect 10968 39933 10977 39967
rect 10977 39933 11011 39967
rect 11011 39933 11020 39967
rect 10968 39924 11020 39933
rect 15384 39924 15436 39976
rect 16028 39967 16080 39976
rect 16028 39933 16037 39967
rect 16037 39933 16071 39967
rect 16071 39933 16080 39967
rect 16028 39924 16080 39933
rect 8484 39856 8536 39908
rect 18420 39924 18472 39976
rect 18788 39967 18840 39976
rect 18788 39933 18797 39967
rect 18797 39933 18831 39967
rect 18831 39933 18840 39967
rect 18788 39924 18840 39933
rect 20260 40035 20312 40044
rect 20260 40001 20269 40035
rect 20269 40001 20303 40035
rect 20303 40001 20312 40035
rect 20260 39992 20312 40001
rect 21180 40060 21232 40112
rect 23664 40128 23716 40180
rect 23756 40128 23808 40180
rect 22836 40060 22888 40112
rect 21364 39992 21416 40044
rect 21732 39992 21784 40044
rect 22744 39992 22796 40044
rect 24492 40060 24544 40112
rect 13728 39788 13780 39840
rect 18236 39899 18288 39908
rect 18236 39865 18245 39899
rect 18245 39865 18279 39899
rect 18279 39865 18288 39899
rect 18236 39856 18288 39865
rect 14648 39831 14700 39840
rect 14648 39797 14657 39831
rect 14657 39797 14691 39831
rect 14691 39797 14700 39831
rect 14648 39788 14700 39797
rect 14832 39788 14884 39840
rect 16304 39788 16356 39840
rect 17132 39788 17184 39840
rect 20444 39967 20496 39976
rect 20444 39933 20453 39967
rect 20453 39933 20487 39967
rect 20487 39933 20496 39967
rect 20444 39924 20496 39933
rect 20536 39924 20588 39976
rect 21548 39924 21600 39976
rect 22652 39924 22704 39976
rect 23020 39924 23072 39976
rect 24492 39924 24544 39976
rect 19524 39856 19576 39908
rect 19064 39788 19116 39840
rect 21824 39856 21876 39908
rect 20260 39788 20312 39840
rect 23756 39788 23808 39840
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 6552 39584 6604 39636
rect 8484 39584 8536 39636
rect 12256 39584 12308 39636
rect 13084 39627 13136 39636
rect 13084 39593 13093 39627
rect 13093 39593 13127 39627
rect 13127 39593 13136 39627
rect 13084 39584 13136 39593
rect 14280 39584 14332 39636
rect 14556 39584 14608 39636
rect 14740 39584 14792 39636
rect 18512 39584 18564 39636
rect 19064 39627 19116 39636
rect 19064 39593 19073 39627
rect 19073 39593 19107 39627
rect 19107 39593 19116 39627
rect 19064 39584 19116 39593
rect 19616 39584 19668 39636
rect 20444 39627 20496 39636
rect 20444 39593 20453 39627
rect 20453 39593 20487 39627
rect 20487 39593 20496 39627
rect 20444 39584 20496 39593
rect 22284 39584 22336 39636
rect 6184 39448 6236 39500
rect 9220 39448 9272 39500
rect 10324 39491 10376 39500
rect 10324 39457 10333 39491
rect 10333 39457 10367 39491
rect 10367 39457 10376 39491
rect 10324 39448 10376 39457
rect 12440 39448 12492 39500
rect 13820 39516 13872 39568
rect 15844 39516 15896 39568
rect 16028 39516 16080 39568
rect 25136 39516 25188 39568
rect 13452 39448 13504 39500
rect 15660 39448 15712 39500
rect 17776 39448 17828 39500
rect 19432 39448 19484 39500
rect 20076 39491 20128 39500
rect 20076 39457 20085 39491
rect 20085 39457 20119 39491
rect 20119 39457 20128 39491
rect 20076 39448 20128 39457
rect 21548 39448 21600 39500
rect 22192 39448 22244 39500
rect 23480 39448 23532 39500
rect 25044 39491 25096 39500
rect 25044 39457 25053 39491
rect 25053 39457 25087 39491
rect 25087 39457 25096 39491
rect 25044 39448 25096 39457
rect 25228 39491 25280 39500
rect 25228 39457 25237 39491
rect 25237 39457 25271 39491
rect 25271 39457 25280 39491
rect 25228 39448 25280 39457
rect 7288 39312 7340 39364
rect 5816 39244 5868 39296
rect 8300 39244 8352 39296
rect 11520 39312 11572 39364
rect 15844 39380 15896 39432
rect 15016 39312 15068 39364
rect 17040 39312 17092 39364
rect 20260 39380 20312 39432
rect 13820 39287 13872 39296
rect 13820 39253 13829 39287
rect 13829 39253 13863 39287
rect 13863 39253 13872 39287
rect 13820 39244 13872 39253
rect 14740 39287 14792 39296
rect 14740 39253 14749 39287
rect 14749 39253 14783 39287
rect 14783 39253 14792 39287
rect 14740 39244 14792 39253
rect 15384 39244 15436 39296
rect 16028 39287 16080 39296
rect 16028 39253 16037 39287
rect 16037 39253 16071 39287
rect 16071 39253 16080 39287
rect 16028 39244 16080 39253
rect 18420 39244 18472 39296
rect 19892 39244 19944 39296
rect 21732 39355 21784 39364
rect 21732 39321 21741 39355
rect 21741 39321 21775 39355
rect 21775 39321 21784 39355
rect 21732 39312 21784 39321
rect 22744 39312 22796 39364
rect 24768 39244 24820 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 7288 39083 7340 39092
rect 7288 39049 7297 39083
rect 7297 39049 7331 39083
rect 7331 39049 7340 39083
rect 7288 39040 7340 39049
rect 9496 39083 9548 39092
rect 9496 39049 9505 39083
rect 9505 39049 9539 39083
rect 9539 39049 9548 39083
rect 9496 39040 9548 39049
rect 10968 39040 11020 39092
rect 11520 38972 11572 39024
rect 4068 38904 4120 38956
rect 9496 38768 9548 38820
rect 1400 38743 1452 38752
rect 1400 38709 1409 38743
rect 1409 38709 1443 38743
rect 1443 38709 1452 38743
rect 1400 38700 1452 38709
rect 9128 38743 9180 38752
rect 9128 38709 9137 38743
rect 9137 38709 9171 38743
rect 9171 38709 9180 38743
rect 9128 38700 9180 38709
rect 9680 38879 9732 38888
rect 9680 38845 9689 38879
rect 9689 38845 9723 38879
rect 9723 38845 9732 38879
rect 9680 38836 9732 38845
rect 10968 38836 11020 38888
rect 13728 39040 13780 39092
rect 14740 39040 14792 39092
rect 14832 39040 14884 39092
rect 15016 39040 15068 39092
rect 15936 39040 15988 39092
rect 16028 39040 16080 39092
rect 20996 39040 21048 39092
rect 22100 39040 22152 39092
rect 12440 38972 12492 39024
rect 13084 38972 13136 39024
rect 18512 38972 18564 39024
rect 20812 38972 20864 39024
rect 23664 38972 23716 39024
rect 25412 38972 25464 39024
rect 21364 38904 21416 38956
rect 14648 38836 14700 38888
rect 11152 38768 11204 38820
rect 11980 38768 12032 38820
rect 11520 38743 11572 38752
rect 11520 38709 11529 38743
rect 11529 38709 11563 38743
rect 11563 38709 11572 38743
rect 11520 38700 11572 38709
rect 11704 38700 11756 38752
rect 15568 38879 15620 38888
rect 15568 38845 15577 38879
rect 15577 38845 15611 38879
rect 15611 38845 15620 38879
rect 15568 38836 15620 38845
rect 16856 38879 16908 38888
rect 16856 38845 16865 38879
rect 16865 38845 16899 38879
rect 16899 38845 16908 38879
rect 16856 38836 16908 38845
rect 18420 38879 18472 38888
rect 18420 38845 18429 38879
rect 18429 38845 18463 38879
rect 18463 38845 18472 38879
rect 18420 38836 18472 38845
rect 19156 38836 19208 38888
rect 18328 38768 18380 38820
rect 20444 38836 20496 38888
rect 20996 38879 21048 38888
rect 20996 38845 21005 38879
rect 21005 38845 21039 38879
rect 21039 38845 21048 38879
rect 20996 38836 21048 38845
rect 14004 38700 14056 38752
rect 16028 38743 16080 38752
rect 16028 38709 16037 38743
rect 16037 38709 16071 38743
rect 16071 38709 16080 38743
rect 16028 38700 16080 38709
rect 16580 38700 16632 38752
rect 18512 38700 18564 38752
rect 18696 38700 18748 38752
rect 20352 38743 20404 38752
rect 20352 38709 20361 38743
rect 20361 38709 20395 38743
rect 20395 38709 20404 38743
rect 20352 38700 20404 38709
rect 20444 38700 20496 38752
rect 22100 38700 22152 38752
rect 23112 38836 23164 38888
rect 23756 38836 23808 38888
rect 24216 38904 24268 38956
rect 24860 38904 24912 38956
rect 25320 38947 25372 38956
rect 25320 38913 25329 38947
rect 25329 38913 25363 38947
rect 25363 38913 25372 38947
rect 25320 38904 25372 38913
rect 24584 38836 24636 38888
rect 22836 38700 22888 38752
rect 23664 38700 23716 38752
rect 25136 38743 25188 38752
rect 25136 38709 25145 38743
rect 25145 38709 25179 38743
rect 25179 38709 25188 38743
rect 25136 38700 25188 38709
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 6920 38496 6972 38548
rect 7196 38496 7248 38548
rect 7748 38496 7800 38548
rect 9864 38496 9916 38548
rect 10324 38496 10376 38548
rect 11060 38496 11112 38548
rect 12348 38496 12400 38548
rect 15844 38496 15896 38548
rect 8576 38428 8628 38480
rect 10140 38428 10192 38480
rect 6920 38360 6972 38412
rect 7840 38360 7892 38412
rect 1308 38292 1360 38344
rect 1768 38156 1820 38208
rect 8300 38292 8352 38344
rect 7380 38224 7432 38276
rect 7564 38224 7616 38276
rect 9128 38360 9180 38412
rect 9220 38292 9272 38344
rect 10232 38360 10284 38412
rect 13452 38428 13504 38480
rect 17868 38496 17920 38548
rect 12164 38360 12216 38412
rect 13268 38403 13320 38412
rect 13268 38369 13277 38403
rect 13277 38369 13311 38403
rect 13311 38369 13320 38403
rect 13268 38360 13320 38369
rect 14280 38360 14332 38412
rect 12716 38292 12768 38344
rect 15200 38292 15252 38344
rect 11980 38224 12032 38276
rect 15108 38224 15160 38276
rect 15660 38224 15712 38276
rect 18328 38360 18380 38412
rect 15936 38335 15988 38344
rect 15936 38301 15945 38335
rect 15945 38301 15979 38335
rect 15979 38301 15988 38335
rect 15936 38292 15988 38301
rect 17316 38292 17368 38344
rect 20812 38428 20864 38480
rect 18696 38403 18748 38412
rect 18696 38369 18705 38403
rect 18705 38369 18739 38403
rect 18739 38369 18748 38403
rect 18696 38360 18748 38369
rect 18880 38360 18932 38412
rect 21088 38403 21140 38412
rect 21088 38369 21097 38403
rect 21097 38369 21131 38403
rect 21131 38369 21140 38403
rect 21088 38360 21140 38369
rect 21272 38403 21324 38412
rect 21272 38369 21281 38403
rect 21281 38369 21315 38403
rect 21315 38369 21324 38403
rect 21272 38360 21324 38369
rect 19064 38292 19116 38344
rect 20444 38292 20496 38344
rect 20628 38292 20680 38344
rect 25964 38496 26016 38548
rect 22284 38428 22336 38480
rect 24676 38428 24728 38480
rect 21916 38360 21968 38412
rect 22652 38403 22704 38412
rect 22652 38369 22661 38403
rect 22661 38369 22695 38403
rect 22695 38369 22704 38403
rect 22652 38360 22704 38369
rect 23664 38360 23716 38412
rect 23756 38403 23808 38412
rect 23756 38369 23765 38403
rect 23765 38369 23799 38403
rect 23799 38369 23808 38403
rect 23756 38360 23808 38369
rect 24952 38360 25004 38412
rect 23848 38292 23900 38344
rect 6552 38156 6604 38208
rect 7196 38156 7248 38208
rect 8208 38156 8260 38208
rect 8484 38156 8536 38208
rect 10692 38156 10744 38208
rect 10784 38199 10836 38208
rect 10784 38165 10793 38199
rect 10793 38165 10827 38199
rect 10827 38165 10836 38199
rect 10784 38156 10836 38165
rect 11060 38156 11112 38208
rect 14556 38156 14608 38208
rect 19248 38224 19300 38276
rect 19340 38224 19392 38276
rect 17776 38156 17828 38208
rect 18788 38156 18840 38208
rect 21088 38156 21140 38208
rect 21916 38156 21968 38208
rect 23940 38224 23992 38276
rect 23572 38199 23624 38208
rect 23572 38165 23581 38199
rect 23581 38165 23615 38199
rect 23615 38165 23624 38199
rect 23572 38156 23624 38165
rect 23664 38199 23716 38208
rect 23664 38165 23673 38199
rect 23673 38165 23707 38199
rect 23707 38165 23716 38199
rect 23664 38156 23716 38165
rect 23756 38156 23808 38208
rect 24676 38156 24728 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 5264 37995 5316 38004
rect 5264 37961 5273 37995
rect 5273 37961 5307 37995
rect 5307 37961 5316 37995
rect 5264 37952 5316 37961
rect 9128 37952 9180 38004
rect 10508 37952 10560 38004
rect 10784 37952 10836 38004
rect 12440 37952 12492 38004
rect 6920 37884 6972 37936
rect 7564 37884 7616 37936
rect 1768 37859 1820 37868
rect 1768 37825 1777 37859
rect 1777 37825 1811 37859
rect 1811 37825 1820 37859
rect 1768 37816 1820 37825
rect 4988 37816 5040 37868
rect 5816 37791 5868 37800
rect 5816 37757 5825 37791
rect 5825 37757 5859 37791
rect 5859 37757 5868 37791
rect 5816 37748 5868 37757
rect 6552 37791 6604 37800
rect 6552 37757 6561 37791
rect 6561 37757 6595 37791
rect 6595 37757 6604 37791
rect 6552 37748 6604 37757
rect 7380 37748 7432 37800
rect 7564 37748 7616 37800
rect 7840 37748 7892 37800
rect 9588 37884 9640 37936
rect 9312 37816 9364 37868
rect 10508 37859 10560 37868
rect 10508 37825 10517 37859
rect 10517 37825 10551 37859
rect 10551 37825 10560 37859
rect 10508 37816 10560 37825
rect 2688 37612 2740 37664
rect 6644 37612 6696 37664
rect 10048 37612 10100 37664
rect 10232 37612 10284 37664
rect 11244 37927 11296 37936
rect 11244 37893 11253 37927
rect 11253 37893 11287 37927
rect 11287 37893 11296 37927
rect 11244 37884 11296 37893
rect 13544 37952 13596 38004
rect 13728 37952 13780 38004
rect 14372 37952 14424 38004
rect 15476 37952 15528 38004
rect 16120 37952 16172 38004
rect 16672 37952 16724 38004
rect 16856 37952 16908 38004
rect 17316 37952 17368 38004
rect 18236 37952 18288 38004
rect 18696 37952 18748 38004
rect 12716 37859 12768 37868
rect 12716 37825 12725 37859
rect 12725 37825 12759 37859
rect 12759 37825 12768 37859
rect 12716 37816 12768 37825
rect 16304 37816 16356 37868
rect 16488 37816 16540 37868
rect 17408 37816 17460 37868
rect 18880 37884 18932 37936
rect 20628 37952 20680 38004
rect 21548 37995 21600 38004
rect 21548 37961 21557 37995
rect 21557 37961 21591 37995
rect 21591 37961 21600 37995
rect 21548 37952 21600 37961
rect 24676 37952 24728 38004
rect 21456 37884 21508 37936
rect 22468 37927 22520 37936
rect 18696 37816 18748 37868
rect 20260 37816 20312 37868
rect 13452 37748 13504 37800
rect 13544 37791 13596 37800
rect 13544 37757 13553 37791
rect 13553 37757 13587 37791
rect 13587 37757 13596 37791
rect 13544 37748 13596 37757
rect 15568 37748 15620 37800
rect 16120 37748 16172 37800
rect 16672 37748 16724 37800
rect 18972 37748 19024 37800
rect 20536 37748 20588 37800
rect 21548 37748 21600 37800
rect 17868 37723 17920 37732
rect 17868 37689 17877 37723
rect 17877 37689 17911 37723
rect 17911 37689 17920 37723
rect 17868 37680 17920 37689
rect 12072 37612 12124 37664
rect 12348 37655 12400 37664
rect 12348 37621 12357 37655
rect 12357 37621 12391 37655
rect 12391 37621 12400 37655
rect 12348 37612 12400 37621
rect 15016 37655 15068 37664
rect 15016 37621 15025 37655
rect 15025 37621 15059 37655
rect 15059 37621 15068 37655
rect 15016 37612 15068 37621
rect 16304 37612 16356 37664
rect 18604 37680 18656 37732
rect 19064 37680 19116 37732
rect 21640 37680 21692 37732
rect 18696 37655 18748 37664
rect 18696 37621 18705 37655
rect 18705 37621 18739 37655
rect 18739 37621 18748 37655
rect 18696 37612 18748 37621
rect 18972 37612 19024 37664
rect 19432 37612 19484 37664
rect 20168 37612 20220 37664
rect 22008 37612 22060 37664
rect 22468 37893 22477 37927
rect 22477 37893 22511 37927
rect 22511 37893 22520 37927
rect 22468 37884 22520 37893
rect 24584 37884 24636 37936
rect 22744 37816 22796 37868
rect 23296 37816 23348 37868
rect 22468 37748 22520 37800
rect 22836 37748 22888 37800
rect 23848 37791 23900 37800
rect 23848 37757 23857 37791
rect 23857 37757 23891 37791
rect 23891 37757 23900 37791
rect 23848 37748 23900 37757
rect 24492 37748 24544 37800
rect 23480 37612 23532 37664
rect 23664 37612 23716 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 8576 37451 8628 37460
rect 8576 37417 8585 37451
rect 8585 37417 8619 37451
rect 8619 37417 8628 37451
rect 8576 37408 8628 37417
rect 8668 37408 8720 37460
rect 10416 37451 10468 37460
rect 10416 37417 10425 37451
rect 10425 37417 10459 37451
rect 10459 37417 10468 37451
rect 10416 37408 10468 37417
rect 10876 37451 10928 37460
rect 10876 37417 10885 37451
rect 10885 37417 10919 37451
rect 10919 37417 10928 37451
rect 10876 37408 10928 37417
rect 15108 37408 15160 37460
rect 16304 37408 16356 37460
rect 23480 37408 23532 37460
rect 23572 37408 23624 37460
rect 24676 37451 24728 37460
rect 24676 37417 24685 37451
rect 24685 37417 24719 37451
rect 24719 37417 24728 37451
rect 24676 37408 24728 37417
rect 8852 37340 8904 37392
rect 11520 37340 11572 37392
rect 8668 37272 8720 37324
rect 9404 37272 9456 37324
rect 10876 37272 10928 37324
rect 13820 37340 13872 37392
rect 14832 37340 14884 37392
rect 16396 37340 16448 37392
rect 13912 37272 13964 37324
rect 6552 37204 6604 37256
rect 7564 37136 7616 37188
rect 10416 37136 10468 37188
rect 10692 37136 10744 37188
rect 10784 37068 10836 37120
rect 11244 37111 11296 37120
rect 11244 37077 11253 37111
rect 11253 37077 11287 37111
rect 11287 37077 11296 37111
rect 11244 37068 11296 37077
rect 11704 37179 11756 37188
rect 11704 37145 11713 37179
rect 11713 37145 11747 37179
rect 11747 37145 11756 37179
rect 11704 37136 11756 37145
rect 13084 37136 13136 37188
rect 13544 37204 13596 37256
rect 15016 37272 15068 37324
rect 15200 37272 15252 37324
rect 16212 37272 16264 37324
rect 20536 37340 20588 37392
rect 21548 37340 21600 37392
rect 25044 37340 25096 37392
rect 17868 37315 17920 37324
rect 17868 37281 17877 37315
rect 17877 37281 17911 37315
rect 17911 37281 17920 37315
rect 17868 37272 17920 37281
rect 12716 37068 12768 37120
rect 20260 37272 20312 37324
rect 24032 37272 24084 37324
rect 20720 37204 20772 37256
rect 17592 37136 17644 37188
rect 14556 37068 14608 37120
rect 14924 37111 14976 37120
rect 14924 37077 14933 37111
rect 14933 37077 14967 37111
rect 14967 37077 14976 37111
rect 14924 37068 14976 37077
rect 15476 37068 15528 37120
rect 16396 37068 16448 37120
rect 17316 37111 17368 37120
rect 17316 37077 17325 37111
rect 17325 37077 17359 37111
rect 17359 37077 17368 37111
rect 17316 37068 17368 37077
rect 18512 37111 18564 37120
rect 18512 37077 18521 37111
rect 18521 37077 18555 37111
rect 18555 37077 18564 37111
rect 18512 37068 18564 37077
rect 19432 37179 19484 37188
rect 19432 37145 19441 37179
rect 19441 37145 19475 37179
rect 19475 37145 19484 37179
rect 19432 37136 19484 37145
rect 20168 37179 20220 37188
rect 20168 37145 20177 37179
rect 20177 37145 20211 37179
rect 20211 37145 20220 37179
rect 20168 37136 20220 37145
rect 20812 37136 20864 37188
rect 21180 37136 21232 37188
rect 22836 37136 22888 37188
rect 20076 37068 20128 37120
rect 23940 37068 23992 37120
rect 25320 37247 25372 37256
rect 25320 37213 25329 37247
rect 25329 37213 25363 37247
rect 25363 37213 25372 37247
rect 25320 37204 25372 37213
rect 25320 37068 25372 37120
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 5540 36864 5592 36916
rect 6552 36864 6604 36916
rect 7472 36907 7524 36916
rect 7472 36873 7481 36907
rect 7481 36873 7515 36907
rect 7515 36873 7524 36907
rect 7472 36864 7524 36873
rect 8484 36864 8536 36916
rect 9036 36907 9088 36916
rect 9036 36873 9045 36907
rect 9045 36873 9079 36907
rect 9079 36873 9088 36907
rect 9036 36864 9088 36873
rect 12716 36864 12768 36916
rect 13544 36864 13596 36916
rect 14188 36864 14240 36916
rect 15108 36864 15160 36916
rect 15200 36864 15252 36916
rect 17040 36907 17092 36916
rect 17040 36873 17049 36907
rect 17049 36873 17083 36907
rect 17083 36873 17092 36907
rect 17040 36864 17092 36873
rect 18512 36864 18564 36916
rect 20444 36864 20496 36916
rect 23940 36864 23992 36916
rect 5632 36796 5684 36848
rect 7564 36796 7616 36848
rect 10416 36796 10468 36848
rect 7840 36771 7892 36780
rect 7840 36737 7849 36771
rect 7849 36737 7883 36771
rect 7883 36737 7892 36771
rect 7840 36728 7892 36737
rect 9312 36728 9364 36780
rect 5264 36660 5316 36712
rect 5816 36660 5868 36712
rect 6000 36660 6052 36712
rect 7380 36592 7432 36644
rect 9404 36592 9456 36644
rect 9588 36703 9640 36712
rect 9588 36669 9597 36703
rect 9597 36669 9631 36703
rect 9631 36669 9640 36703
rect 9588 36660 9640 36669
rect 10968 36703 11020 36712
rect 10968 36669 10977 36703
rect 10977 36669 11011 36703
rect 11011 36669 11020 36703
rect 10968 36660 11020 36669
rect 13084 36796 13136 36848
rect 17316 36796 17368 36848
rect 24676 36796 24728 36848
rect 12072 36728 12124 36780
rect 11888 36703 11940 36712
rect 11888 36669 11897 36703
rect 11897 36669 11931 36703
rect 11931 36669 11940 36703
rect 11888 36660 11940 36669
rect 12808 36703 12860 36712
rect 12808 36669 12817 36703
rect 12817 36669 12851 36703
rect 12851 36669 12860 36703
rect 12808 36660 12860 36669
rect 13912 36728 13964 36780
rect 16672 36771 16724 36780
rect 16672 36737 16681 36771
rect 16681 36737 16715 36771
rect 16715 36737 16724 36771
rect 16672 36728 16724 36737
rect 19800 36728 19852 36780
rect 25320 36771 25372 36780
rect 25320 36737 25329 36771
rect 25329 36737 25363 36771
rect 25363 36737 25372 36771
rect 25320 36728 25372 36737
rect 14004 36703 14056 36712
rect 14004 36669 14013 36703
rect 14013 36669 14047 36703
rect 14047 36669 14056 36703
rect 14004 36660 14056 36669
rect 14556 36660 14608 36712
rect 15200 36703 15252 36712
rect 15200 36669 15209 36703
rect 15209 36669 15243 36703
rect 15243 36669 15252 36703
rect 15200 36660 15252 36669
rect 15844 36703 15896 36712
rect 15844 36669 15853 36703
rect 15853 36669 15887 36703
rect 15887 36669 15896 36703
rect 15844 36660 15896 36669
rect 17684 36703 17736 36712
rect 17684 36669 17693 36703
rect 17693 36669 17727 36703
rect 17727 36669 17736 36703
rect 17684 36660 17736 36669
rect 18512 36660 18564 36712
rect 22836 36703 22888 36712
rect 22836 36669 22845 36703
rect 22845 36669 22879 36703
rect 22879 36669 22888 36703
rect 22836 36660 22888 36669
rect 16028 36592 16080 36644
rect 19432 36592 19484 36644
rect 20444 36592 20496 36644
rect 22468 36592 22520 36644
rect 23572 36660 23624 36712
rect 23848 36660 23900 36712
rect 1584 36524 1636 36576
rect 8668 36567 8720 36576
rect 8668 36533 8677 36567
rect 8677 36533 8711 36567
rect 8711 36533 8720 36567
rect 8668 36524 8720 36533
rect 10876 36524 10928 36576
rect 14280 36524 14332 36576
rect 14556 36567 14608 36576
rect 14556 36533 14565 36567
rect 14565 36533 14599 36567
rect 14599 36533 14608 36567
rect 14556 36524 14608 36533
rect 17224 36524 17276 36576
rect 20076 36524 20128 36576
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 7656 36363 7708 36372
rect 7656 36329 7665 36363
rect 7665 36329 7699 36363
rect 7699 36329 7708 36363
rect 7656 36320 7708 36329
rect 9128 36363 9180 36372
rect 9128 36329 9137 36363
rect 9137 36329 9171 36363
rect 9171 36329 9180 36363
rect 9128 36320 9180 36329
rect 12532 36320 12584 36372
rect 13360 36320 13412 36372
rect 13544 36320 13596 36372
rect 7104 36252 7156 36304
rect 7564 36184 7616 36236
rect 1584 36159 1636 36168
rect 1584 36125 1593 36159
rect 1593 36125 1627 36159
rect 1627 36125 1636 36159
rect 1584 36116 1636 36125
rect 7380 36116 7432 36168
rect 12716 36184 12768 36236
rect 13544 36184 13596 36236
rect 12348 36116 12400 36168
rect 15384 36320 15436 36372
rect 18788 36320 18840 36372
rect 19248 36320 19300 36372
rect 13820 36295 13872 36304
rect 13820 36261 13829 36295
rect 13829 36261 13863 36295
rect 13863 36261 13872 36295
rect 13820 36252 13872 36261
rect 16948 36252 17000 36304
rect 15660 36184 15712 36236
rect 19708 36184 19760 36236
rect 10416 36048 10468 36100
rect 1768 35980 1820 36032
rect 7472 35980 7524 36032
rect 11336 35980 11388 36032
rect 12716 35980 12768 36032
rect 14648 36023 14700 36032
rect 14648 35989 14657 36023
rect 14657 35989 14691 36023
rect 14691 35989 14700 36023
rect 14648 35980 14700 35989
rect 15660 36048 15712 36100
rect 21732 36320 21784 36372
rect 20352 36184 20404 36236
rect 21364 36227 21416 36236
rect 21364 36193 21373 36227
rect 21373 36193 21407 36227
rect 21407 36193 21416 36227
rect 21364 36184 21416 36193
rect 20904 36116 20956 36168
rect 23204 36320 23256 36372
rect 25136 36320 25188 36372
rect 24400 36252 24452 36304
rect 23756 36227 23808 36236
rect 23756 36193 23765 36227
rect 23765 36193 23799 36227
rect 23799 36193 23808 36227
rect 23756 36184 23808 36193
rect 24492 36184 24544 36236
rect 24124 36116 24176 36168
rect 25320 36159 25372 36168
rect 25320 36125 25329 36159
rect 25329 36125 25363 36159
rect 25363 36125 25372 36159
rect 25320 36116 25372 36125
rect 19616 35980 19668 36032
rect 20904 35980 20956 36032
rect 21824 36048 21876 36100
rect 22284 35980 22336 36032
rect 23204 35980 23256 36032
rect 23664 36023 23716 36032
rect 23664 35989 23673 36023
rect 23673 35989 23707 36023
rect 23707 35989 23716 36023
rect 23664 35980 23716 35989
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 1768 35683 1820 35692
rect 1768 35649 1777 35683
rect 1777 35649 1811 35683
rect 1811 35649 1820 35683
rect 1768 35640 1820 35649
rect 5540 35776 5592 35828
rect 6000 35819 6052 35828
rect 6000 35785 6009 35819
rect 6009 35785 6043 35819
rect 6043 35785 6052 35819
rect 6000 35776 6052 35785
rect 7288 35776 7340 35828
rect 8576 35776 8628 35828
rect 10232 35776 10284 35828
rect 5632 35640 5684 35692
rect 6920 35640 6972 35692
rect 13452 35776 13504 35828
rect 13544 35776 13596 35828
rect 14648 35776 14700 35828
rect 17592 35776 17644 35828
rect 17408 35708 17460 35760
rect 17776 35708 17828 35760
rect 18328 35708 18380 35760
rect 19984 35708 20036 35760
rect 5816 35572 5868 35624
rect 4068 35436 4120 35488
rect 9588 35572 9640 35624
rect 8576 35436 8628 35488
rect 9772 35436 9824 35488
rect 10968 35572 11020 35624
rect 11980 35615 12032 35624
rect 11980 35581 11989 35615
rect 11989 35581 12023 35615
rect 12023 35581 12032 35615
rect 11980 35572 12032 35581
rect 10232 35479 10284 35488
rect 10232 35445 10241 35479
rect 10241 35445 10275 35479
rect 10275 35445 10284 35479
rect 10232 35436 10284 35445
rect 10784 35436 10836 35488
rect 11704 35436 11756 35488
rect 13636 35436 13688 35488
rect 15200 35572 15252 35624
rect 17408 35572 17460 35624
rect 21548 35640 21600 35692
rect 13912 35436 13964 35488
rect 15936 35436 15988 35488
rect 19156 35504 19208 35556
rect 17960 35436 18012 35488
rect 19800 35479 19852 35488
rect 19800 35445 19809 35479
rect 19809 35445 19843 35479
rect 19843 35445 19852 35479
rect 19800 35436 19852 35445
rect 22192 35776 22244 35828
rect 23572 35776 23624 35828
rect 24676 35708 24728 35760
rect 25228 35708 25280 35760
rect 22100 35640 22152 35692
rect 22192 35640 22244 35692
rect 22836 35640 22888 35692
rect 22468 35615 22520 35624
rect 22468 35581 22477 35615
rect 22477 35581 22511 35615
rect 22511 35581 22520 35615
rect 22468 35572 22520 35581
rect 23388 35615 23440 35624
rect 23388 35581 23397 35615
rect 23397 35581 23431 35615
rect 23431 35581 23440 35615
rect 23388 35572 23440 35581
rect 22376 35504 22428 35556
rect 22560 35504 22612 35556
rect 22836 35504 22888 35556
rect 20720 35436 20772 35488
rect 25228 35479 25280 35488
rect 25228 35445 25237 35479
rect 25237 35445 25271 35479
rect 25271 35445 25280 35479
rect 25228 35436 25280 35445
rect 25320 35436 25372 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 7380 35232 7432 35284
rect 8760 35232 8812 35284
rect 9404 35232 9456 35284
rect 16120 35232 16172 35284
rect 11980 35164 12032 35216
rect 13820 35164 13872 35216
rect 5540 35096 5592 35148
rect 6092 35139 6144 35148
rect 6092 35105 6101 35139
rect 6101 35105 6135 35139
rect 6135 35105 6144 35139
rect 6092 35096 6144 35105
rect 9772 35096 9824 35148
rect 9864 35139 9916 35148
rect 9864 35105 9873 35139
rect 9873 35105 9907 35139
rect 9907 35105 9916 35139
rect 9864 35096 9916 35105
rect 11152 35096 11204 35148
rect 15752 35096 15804 35148
rect 14556 35028 14608 35080
rect 18328 35232 18380 35284
rect 19708 35232 19760 35284
rect 20352 35232 20404 35284
rect 21640 35275 21692 35284
rect 21640 35241 21649 35275
rect 21649 35241 21683 35275
rect 21683 35241 21692 35275
rect 21640 35232 21692 35241
rect 20720 35164 20772 35216
rect 17960 35096 18012 35148
rect 18328 35096 18380 35148
rect 20168 35096 20220 35148
rect 22192 35028 22244 35080
rect 6920 34960 6972 35012
rect 8668 34960 8720 35012
rect 14188 34960 14240 35012
rect 7012 34892 7064 34944
rect 8300 34892 8352 34944
rect 10692 34892 10744 34944
rect 13360 34935 13412 34944
rect 13360 34901 13369 34935
rect 13369 34901 13403 34935
rect 13403 34901 13412 34935
rect 13360 34892 13412 34901
rect 19708 35003 19760 35012
rect 19708 34969 19717 35003
rect 19717 34969 19751 35003
rect 19751 34969 19760 35003
rect 19708 34960 19760 34969
rect 19892 34892 19944 34944
rect 20720 34960 20772 35012
rect 21272 34960 21324 35012
rect 22652 34960 22704 35012
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 25228 34960 25280 35012
rect 20996 34892 21048 34944
rect 21364 34892 21416 34944
rect 22376 34892 22428 34944
rect 23204 34892 23256 34944
rect 23388 34892 23440 34944
rect 24308 34892 24360 34944
rect 24492 34892 24544 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 7196 34688 7248 34740
rect 8300 34731 8352 34740
rect 8300 34697 8309 34731
rect 8309 34697 8343 34731
rect 8343 34697 8352 34731
rect 8300 34688 8352 34697
rect 9496 34688 9548 34740
rect 10692 34688 10744 34740
rect 12808 34688 12860 34740
rect 13728 34688 13780 34740
rect 19800 34688 19852 34740
rect 20260 34731 20312 34740
rect 20260 34697 20269 34731
rect 20269 34697 20303 34731
rect 20303 34697 20312 34731
rect 20260 34688 20312 34697
rect 20812 34688 20864 34740
rect 21180 34688 21232 34740
rect 22284 34688 22336 34740
rect 23664 34688 23716 34740
rect 24676 34688 24728 34740
rect 6000 34620 6052 34672
rect 6920 34620 6972 34672
rect 8484 34620 8536 34672
rect 12072 34620 12124 34672
rect 13912 34620 13964 34672
rect 16580 34620 16632 34672
rect 17960 34620 18012 34672
rect 19708 34620 19760 34672
rect 22100 34620 22152 34672
rect 22468 34620 22520 34672
rect 6092 34552 6144 34604
rect 8576 34552 8628 34604
rect 13360 34552 13412 34604
rect 17316 34552 17368 34604
rect 21640 34552 21692 34604
rect 23296 34552 23348 34604
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 9588 34484 9640 34536
rect 10968 34484 11020 34536
rect 13820 34484 13872 34536
rect 14832 34484 14884 34536
rect 10140 34348 10192 34400
rect 11152 34416 11204 34468
rect 13360 34416 13412 34468
rect 10784 34348 10836 34400
rect 11796 34348 11848 34400
rect 13912 34348 13964 34400
rect 15476 34348 15528 34400
rect 15568 34391 15620 34400
rect 15568 34357 15577 34391
rect 15577 34357 15611 34391
rect 15611 34357 15620 34391
rect 15568 34348 15620 34357
rect 15844 34416 15896 34468
rect 19524 34416 19576 34468
rect 22468 34527 22520 34536
rect 22468 34493 22477 34527
rect 22477 34493 22511 34527
rect 22511 34493 22520 34527
rect 22468 34484 22520 34493
rect 22652 34527 22704 34536
rect 22652 34493 22661 34527
rect 22661 34493 22695 34527
rect 22695 34493 22704 34527
rect 22652 34484 22704 34493
rect 23480 34484 23532 34536
rect 23848 34527 23900 34536
rect 23848 34493 23857 34527
rect 23857 34493 23891 34527
rect 23891 34493 23900 34527
rect 23848 34484 23900 34493
rect 20168 34348 20220 34400
rect 22008 34391 22060 34400
rect 22008 34357 22017 34391
rect 22017 34357 22051 34391
rect 22051 34357 22060 34391
rect 22008 34348 22060 34357
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 6920 34144 6972 34196
rect 7748 34187 7800 34196
rect 7748 34153 7757 34187
rect 7757 34153 7791 34187
rect 7791 34153 7800 34187
rect 7748 34144 7800 34153
rect 7840 34144 7892 34196
rect 11152 34144 11204 34196
rect 8484 34119 8536 34128
rect 8484 34085 8493 34119
rect 8493 34085 8527 34119
rect 8527 34085 8536 34119
rect 8484 34076 8536 34085
rect 5540 34051 5592 34060
rect 5540 34017 5549 34051
rect 5549 34017 5583 34051
rect 5583 34017 5592 34051
rect 5540 34008 5592 34017
rect 5816 34008 5868 34060
rect 9220 34008 9272 34060
rect 11704 34008 11756 34060
rect 12624 34008 12676 34060
rect 13912 34144 13964 34196
rect 6920 33940 6972 33992
rect 9588 33940 9640 33992
rect 11796 33940 11848 33992
rect 1216 33804 1268 33856
rect 7656 33872 7708 33924
rect 7748 33804 7800 33856
rect 8392 33804 8444 33856
rect 10968 33804 11020 33856
rect 12348 33804 12400 33856
rect 12532 33804 12584 33856
rect 12808 33804 12860 33856
rect 13176 33804 13228 33856
rect 16948 34144 17000 34196
rect 17960 34144 18012 34196
rect 18052 34187 18104 34196
rect 18052 34153 18061 34187
rect 18061 34153 18095 34187
rect 18095 34153 18104 34187
rect 18052 34144 18104 34153
rect 18420 34144 18472 34196
rect 18788 34144 18840 34196
rect 20720 34144 20772 34196
rect 22468 34144 22520 34196
rect 25320 34187 25372 34196
rect 25320 34153 25329 34187
rect 25329 34153 25363 34187
rect 25363 34153 25372 34187
rect 25320 34144 25372 34153
rect 17868 34076 17920 34128
rect 23848 34076 23900 34128
rect 15936 34051 15988 34060
rect 15936 34017 15945 34051
rect 15945 34017 15979 34051
rect 15979 34017 15988 34051
rect 15936 34008 15988 34017
rect 18420 34008 18472 34060
rect 21364 34008 21416 34060
rect 21916 34008 21968 34060
rect 23388 34008 23440 34060
rect 20076 33940 20128 33992
rect 21456 33940 21508 33992
rect 16212 33915 16264 33924
rect 16212 33881 16221 33915
rect 16221 33881 16255 33915
rect 16255 33881 16264 33915
rect 16212 33872 16264 33881
rect 17592 33872 17644 33924
rect 18052 33872 18104 33924
rect 20260 33872 20312 33924
rect 24768 33983 24820 33992
rect 24768 33949 24777 33983
rect 24777 33949 24811 33983
rect 24811 33949 24820 33983
rect 24768 33940 24820 33949
rect 23388 33872 23440 33924
rect 24032 33872 24084 33924
rect 24308 33872 24360 33924
rect 16304 33804 16356 33856
rect 19156 33804 19208 33856
rect 20628 33847 20680 33856
rect 20628 33813 20637 33847
rect 20637 33813 20671 33847
rect 20671 33813 20680 33847
rect 20628 33804 20680 33813
rect 20720 33804 20772 33856
rect 21456 33847 21508 33856
rect 21456 33813 21465 33847
rect 21465 33813 21499 33847
rect 21499 33813 21508 33847
rect 21456 33804 21508 33813
rect 22468 33804 22520 33856
rect 24584 33847 24636 33856
rect 24584 33813 24593 33847
rect 24593 33813 24627 33847
rect 24627 33813 24636 33847
rect 24584 33804 24636 33813
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 6920 33600 6972 33652
rect 10416 33643 10468 33652
rect 10416 33609 10425 33643
rect 10425 33609 10459 33643
rect 10459 33609 10468 33643
rect 10416 33600 10468 33609
rect 10876 33643 10928 33652
rect 10876 33609 10885 33643
rect 10885 33609 10919 33643
rect 10919 33609 10928 33643
rect 10876 33600 10928 33609
rect 11336 33600 11388 33652
rect 13360 33643 13412 33652
rect 13360 33609 13369 33643
rect 13369 33609 13403 33643
rect 13403 33609 13412 33643
rect 13360 33600 13412 33609
rect 10968 33532 11020 33584
rect 12624 33532 12676 33584
rect 1216 33464 1268 33516
rect 11888 33464 11940 33516
rect 12532 33464 12584 33516
rect 14556 33600 14608 33652
rect 15936 33600 15988 33652
rect 15476 33464 15528 33516
rect 15936 33464 15988 33516
rect 17592 33600 17644 33652
rect 19892 33600 19944 33652
rect 18328 33532 18380 33584
rect 18788 33532 18840 33584
rect 5356 33439 5408 33448
rect 5356 33405 5365 33439
rect 5365 33405 5399 33439
rect 5399 33405 5408 33439
rect 5356 33396 5408 33405
rect 9772 33439 9824 33448
rect 9772 33405 9781 33439
rect 9781 33405 9815 33439
rect 9815 33405 9824 33439
rect 9772 33396 9824 33405
rect 8300 33328 8352 33380
rect 13452 33439 13504 33448
rect 13452 33405 13461 33439
rect 13461 33405 13495 33439
rect 13495 33405 13504 33439
rect 13452 33396 13504 33405
rect 16304 33396 16356 33448
rect 21364 33600 21416 33652
rect 21456 33600 21508 33652
rect 25044 33600 25096 33652
rect 20260 33532 20312 33584
rect 20628 33507 20680 33516
rect 20628 33473 20637 33507
rect 20637 33473 20671 33507
rect 20671 33473 20680 33507
rect 20628 33464 20680 33473
rect 24032 33532 24084 33584
rect 21456 33464 21508 33516
rect 22100 33464 22152 33516
rect 22192 33464 22244 33516
rect 20444 33396 20496 33448
rect 21180 33396 21232 33448
rect 23756 33439 23808 33448
rect 23756 33405 23765 33439
rect 23765 33405 23799 33439
rect 23799 33405 23808 33439
rect 23756 33396 23808 33405
rect 15476 33328 15528 33380
rect 15936 33328 15988 33380
rect 1768 33260 1820 33312
rect 7104 33260 7156 33312
rect 10600 33260 10652 33312
rect 12532 33303 12584 33312
rect 12532 33269 12541 33303
rect 12541 33269 12575 33303
rect 12575 33269 12584 33303
rect 12532 33260 12584 33269
rect 13176 33260 13228 33312
rect 13452 33260 13504 33312
rect 13544 33260 13596 33312
rect 15844 33303 15896 33312
rect 15844 33269 15853 33303
rect 15853 33269 15887 33303
rect 15887 33269 15896 33303
rect 15844 33260 15896 33269
rect 23480 33328 23532 33380
rect 21364 33303 21416 33312
rect 21364 33269 21373 33303
rect 21373 33269 21407 33303
rect 21407 33269 21416 33303
rect 21364 33260 21416 33269
rect 22284 33260 22336 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 7472 33099 7524 33108
rect 7472 33065 7481 33099
rect 7481 33065 7515 33099
rect 7515 33065 7524 33099
rect 7472 33056 7524 33065
rect 9312 33056 9364 33108
rect 10600 33099 10652 33108
rect 10600 33065 10609 33099
rect 10609 33065 10643 33099
rect 10643 33065 10652 33099
rect 10600 33056 10652 33065
rect 11060 33056 11112 33108
rect 12256 33099 12308 33108
rect 12256 33065 12265 33099
rect 12265 33065 12299 33099
rect 12299 33065 12308 33099
rect 12256 33056 12308 33065
rect 12440 33056 12492 33108
rect 13912 33056 13964 33108
rect 14004 33056 14056 33108
rect 7564 32988 7616 33040
rect 5540 32920 5592 32972
rect 1768 32895 1820 32904
rect 1768 32861 1777 32895
rect 1777 32861 1811 32895
rect 1811 32861 1820 32895
rect 1768 32852 1820 32861
rect 6920 32852 6972 32904
rect 8300 32920 8352 32972
rect 10140 32920 10192 32972
rect 11612 32963 11664 32972
rect 11612 32929 11621 32963
rect 11621 32929 11655 32963
rect 11655 32929 11664 32963
rect 11612 32920 11664 32929
rect 14924 32988 14976 33040
rect 14280 32920 14332 32972
rect 14832 32963 14884 32972
rect 14832 32929 14841 32963
rect 14841 32929 14875 32963
rect 14875 32929 14884 32963
rect 14832 32920 14884 32929
rect 16488 32920 16540 32972
rect 18512 32920 18564 32972
rect 1584 32759 1636 32768
rect 1584 32725 1593 32759
rect 1593 32725 1627 32759
rect 1627 32725 1636 32759
rect 1584 32716 1636 32725
rect 9772 32895 9824 32904
rect 9772 32861 9781 32895
rect 9781 32861 9815 32895
rect 9815 32861 9824 32895
rect 9772 32852 9824 32861
rect 10600 32852 10652 32904
rect 11980 32852 12032 32904
rect 12532 32852 12584 32904
rect 13636 32852 13688 32904
rect 7748 32784 7800 32836
rect 7840 32759 7892 32768
rect 7840 32725 7849 32759
rect 7849 32725 7883 32759
rect 7883 32725 7892 32759
rect 7840 32716 7892 32725
rect 9496 32716 9548 32768
rect 11612 32716 11664 32768
rect 14004 32716 14056 32768
rect 15844 32784 15896 32836
rect 16764 32852 16816 32904
rect 14648 32759 14700 32768
rect 14648 32725 14657 32759
rect 14657 32725 14691 32759
rect 14691 32725 14700 32759
rect 14648 32716 14700 32725
rect 16120 32759 16172 32768
rect 16120 32725 16129 32759
rect 16129 32725 16163 32759
rect 16163 32725 16172 32759
rect 16120 32716 16172 32725
rect 17592 32784 17644 32836
rect 22468 33056 22520 33108
rect 23572 33056 23624 33108
rect 22100 32988 22152 33040
rect 21272 32920 21324 32972
rect 21548 32963 21600 32972
rect 21548 32929 21557 32963
rect 21557 32929 21591 32963
rect 21591 32929 21600 32963
rect 21548 32920 21600 32929
rect 22284 32988 22336 33040
rect 23664 32988 23716 33040
rect 21180 32852 21232 32904
rect 24032 32920 24084 32972
rect 20628 32784 20680 32836
rect 18604 32716 18656 32768
rect 21916 32716 21968 32768
rect 22376 32891 22428 32904
rect 22376 32857 22385 32891
rect 22385 32857 22419 32891
rect 22419 32857 22428 32891
rect 22376 32852 22428 32857
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 22744 32759 22796 32768
rect 22744 32725 22753 32759
rect 22753 32725 22787 32759
rect 22787 32725 22796 32759
rect 22744 32716 22796 32725
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 4620 32555 4672 32564
rect 4620 32521 4629 32555
rect 4629 32521 4663 32555
rect 4663 32521 4672 32555
rect 4620 32512 4672 32521
rect 4988 32555 5040 32564
rect 4988 32521 4997 32555
rect 4997 32521 5031 32555
rect 5031 32521 5040 32555
rect 4988 32512 5040 32521
rect 5356 32555 5408 32564
rect 5356 32521 5365 32555
rect 5365 32521 5399 32555
rect 5399 32521 5408 32555
rect 5356 32512 5408 32521
rect 7840 32512 7892 32564
rect 14648 32512 14700 32564
rect 14740 32512 14792 32564
rect 5448 32487 5500 32496
rect 5448 32453 5457 32487
rect 5457 32453 5491 32487
rect 5491 32453 5500 32487
rect 5448 32444 5500 32453
rect 5540 32444 5592 32496
rect 9128 32444 9180 32496
rect 6184 32376 6236 32428
rect 5264 32308 5316 32360
rect 8392 32308 8444 32360
rect 9404 32308 9456 32360
rect 7564 32240 7616 32292
rect 9312 32215 9364 32224
rect 9312 32181 9321 32215
rect 9321 32181 9355 32215
rect 9355 32181 9364 32215
rect 9312 32172 9364 32181
rect 13728 32444 13780 32496
rect 15108 32444 15160 32496
rect 17224 32487 17276 32496
rect 17224 32453 17233 32487
rect 17233 32453 17267 32487
rect 17267 32453 17276 32487
rect 17224 32444 17276 32453
rect 14556 32419 14608 32428
rect 14556 32385 14565 32419
rect 14565 32385 14599 32419
rect 14599 32385 14608 32419
rect 14556 32376 14608 32385
rect 15936 32376 15988 32428
rect 18512 32555 18564 32564
rect 18512 32521 18521 32555
rect 18521 32521 18555 32555
rect 18555 32521 18564 32555
rect 18512 32512 18564 32521
rect 21088 32512 21140 32564
rect 21180 32555 21232 32564
rect 21180 32521 21189 32555
rect 21189 32521 21223 32555
rect 21223 32521 21232 32555
rect 21916 32555 21968 32564
rect 21180 32512 21232 32521
rect 21916 32521 21925 32555
rect 21925 32521 21959 32555
rect 21959 32521 21968 32555
rect 21916 32512 21968 32521
rect 22376 32512 22428 32564
rect 22744 32512 22796 32564
rect 9864 32351 9916 32360
rect 9864 32317 9873 32351
rect 9873 32317 9907 32351
rect 9907 32317 9916 32351
rect 9864 32308 9916 32317
rect 12256 32308 12308 32360
rect 12072 32240 12124 32292
rect 14832 32351 14884 32360
rect 14832 32317 14841 32351
rect 14841 32317 14875 32351
rect 14875 32317 14884 32351
rect 14832 32308 14884 32317
rect 16304 32351 16356 32360
rect 16304 32317 16313 32351
rect 16313 32317 16347 32351
rect 16347 32317 16356 32351
rect 16304 32308 16356 32317
rect 16120 32240 16172 32292
rect 17500 32351 17552 32360
rect 17500 32317 17509 32351
rect 17509 32317 17543 32351
rect 17543 32317 17552 32351
rect 17500 32308 17552 32317
rect 18604 32351 18656 32360
rect 18604 32317 18613 32351
rect 18613 32317 18647 32351
rect 18647 32317 18656 32351
rect 18604 32308 18656 32317
rect 20168 32376 20220 32428
rect 21088 32419 21140 32428
rect 21088 32385 21097 32419
rect 21097 32385 21131 32419
rect 21131 32385 21140 32419
rect 21088 32376 21140 32385
rect 21456 32376 21508 32428
rect 22100 32444 22152 32496
rect 22284 32444 22336 32496
rect 17592 32240 17644 32292
rect 21364 32351 21416 32360
rect 21364 32317 21373 32351
rect 21373 32317 21407 32351
rect 21407 32317 21416 32351
rect 21364 32308 21416 32317
rect 22560 32376 22612 32428
rect 25412 32376 25464 32428
rect 25136 32283 25188 32292
rect 25136 32249 25145 32283
rect 25145 32249 25179 32283
rect 25179 32249 25188 32283
rect 25136 32240 25188 32249
rect 10968 32172 11020 32224
rect 12348 32172 12400 32224
rect 13452 32172 13504 32224
rect 14556 32172 14608 32224
rect 15200 32172 15252 32224
rect 16672 32172 16724 32224
rect 18328 32172 18380 32224
rect 20628 32172 20680 32224
rect 20996 32172 21048 32224
rect 21364 32172 21416 32224
rect 21548 32172 21600 32224
rect 22560 32172 22612 32224
rect 22744 32172 22796 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 8300 31968 8352 32020
rect 8392 32011 8444 32020
rect 8392 31977 8401 32011
rect 8401 31977 8435 32011
rect 8435 31977 8444 32011
rect 8392 31968 8444 31977
rect 9128 31968 9180 32020
rect 9404 31968 9456 32020
rect 9680 31968 9732 32020
rect 10140 31968 10192 32020
rect 11888 31968 11940 32020
rect 17592 31968 17644 32020
rect 18236 31968 18288 32020
rect 18604 31968 18656 32020
rect 6184 31875 6236 31884
rect 6184 31841 6193 31875
rect 6193 31841 6227 31875
rect 6227 31841 6236 31875
rect 6184 31832 6236 31841
rect 7196 31832 7248 31884
rect 9312 31900 9364 31952
rect 12164 31900 12216 31952
rect 13820 31900 13872 31952
rect 13912 31943 13964 31952
rect 13912 31909 13921 31943
rect 13921 31909 13955 31943
rect 13955 31909 13964 31943
rect 13912 31900 13964 31909
rect 9772 31832 9824 31884
rect 14188 31900 14240 31952
rect 18788 31900 18840 31952
rect 19432 31943 19484 31952
rect 19432 31909 19441 31943
rect 19441 31909 19475 31943
rect 19475 31909 19484 31943
rect 19432 31900 19484 31909
rect 19892 31900 19944 31952
rect 15108 31832 15160 31884
rect 15660 31764 15712 31816
rect 16764 31764 16816 31816
rect 9588 31696 9640 31748
rect 10968 31696 11020 31748
rect 9128 31671 9180 31680
rect 9128 31637 9137 31671
rect 9137 31637 9171 31671
rect 9171 31637 9180 31671
rect 9128 31628 9180 31637
rect 17408 31696 17460 31748
rect 18880 31696 18932 31748
rect 11704 31628 11756 31680
rect 12440 31628 12492 31680
rect 12716 31628 12768 31680
rect 13820 31628 13872 31680
rect 14924 31628 14976 31680
rect 17224 31628 17276 31680
rect 18236 31671 18288 31680
rect 18236 31637 18245 31671
rect 18245 31637 18279 31671
rect 18279 31637 18288 31671
rect 18236 31628 18288 31637
rect 19156 31628 19208 31680
rect 22560 31968 22612 32020
rect 24308 31968 24360 32020
rect 20260 31900 20312 31952
rect 20996 31900 21048 31952
rect 23388 31900 23440 31952
rect 23572 31900 23624 31952
rect 23480 31832 23532 31884
rect 20904 31764 20956 31816
rect 21640 31764 21692 31816
rect 23940 31764 23992 31816
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 20720 31696 20772 31748
rect 21824 31696 21876 31748
rect 22284 31739 22336 31748
rect 22284 31705 22293 31739
rect 22293 31705 22327 31739
rect 22327 31705 22336 31739
rect 22284 31696 22336 31705
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 7656 31424 7708 31476
rect 8668 31467 8720 31476
rect 8668 31433 8677 31467
rect 8677 31433 8711 31467
rect 8711 31433 8720 31467
rect 8668 31424 8720 31433
rect 9864 31424 9916 31476
rect 12716 31424 12768 31476
rect 13360 31424 13412 31476
rect 14648 31467 14700 31476
rect 14648 31433 14657 31467
rect 14657 31433 14691 31467
rect 14691 31433 14700 31467
rect 14648 31424 14700 31433
rect 16212 31424 16264 31476
rect 17316 31424 17368 31476
rect 21456 31424 21508 31476
rect 21640 31424 21692 31476
rect 23296 31424 23348 31476
rect 1952 31288 2004 31340
rect 7840 31331 7892 31340
rect 7840 31297 7849 31331
rect 7849 31297 7883 31331
rect 7883 31297 7892 31331
rect 7840 31288 7892 31297
rect 1308 31220 1360 31272
rect 9680 31356 9732 31408
rect 11336 31356 11388 31408
rect 15384 31356 15436 31408
rect 20628 31356 20680 31408
rect 21364 31356 21416 31408
rect 23940 31356 23992 31408
rect 8760 31288 8812 31340
rect 9588 31288 9640 31340
rect 14280 31288 14332 31340
rect 15936 31288 15988 31340
rect 4804 31152 4856 31204
rect 8668 31152 8720 31204
rect 8760 31152 8812 31204
rect 5724 31084 5776 31136
rect 13268 31220 13320 31272
rect 13544 31220 13596 31272
rect 14464 31084 14516 31136
rect 15292 31084 15344 31136
rect 17040 31220 17092 31272
rect 17592 31152 17644 31204
rect 17132 31127 17184 31136
rect 17132 31093 17141 31127
rect 17141 31093 17175 31127
rect 17175 31093 17184 31127
rect 17132 31084 17184 31093
rect 19248 31288 19300 31340
rect 21548 31288 21600 31340
rect 24400 31288 24452 31340
rect 25320 31331 25372 31340
rect 25320 31297 25329 31331
rect 25329 31297 25363 31331
rect 25363 31297 25372 31331
rect 25320 31288 25372 31297
rect 18880 31263 18932 31272
rect 18880 31229 18889 31263
rect 18889 31229 18923 31263
rect 18923 31229 18932 31263
rect 18880 31220 18932 31229
rect 19984 31263 20036 31272
rect 19984 31229 19993 31263
rect 19993 31229 20027 31263
rect 20027 31229 20036 31263
rect 19984 31220 20036 31229
rect 20444 31152 20496 31204
rect 22192 31263 22244 31272
rect 22192 31229 22201 31263
rect 22201 31229 22235 31263
rect 22235 31229 22244 31263
rect 22192 31220 22244 31229
rect 19156 31084 19208 31136
rect 20168 31084 20220 31136
rect 20352 31084 20404 31136
rect 20628 31084 20680 31136
rect 22652 31084 22704 31136
rect 23572 31084 23624 31136
rect 24400 31127 24452 31136
rect 24400 31093 24409 31127
rect 24409 31093 24443 31127
rect 24443 31093 24452 31127
rect 24400 31084 24452 31093
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 12624 30880 12676 30932
rect 11704 30855 11756 30864
rect 1860 30744 1912 30796
rect 4620 30787 4672 30796
rect 4620 30753 4629 30787
rect 4629 30753 4663 30787
rect 4663 30753 4672 30787
rect 4620 30744 4672 30753
rect 7840 30744 7892 30796
rect 9588 30787 9640 30796
rect 9588 30753 9597 30787
rect 9597 30753 9631 30787
rect 9631 30753 9640 30787
rect 9588 30744 9640 30753
rect 10876 30744 10928 30796
rect 11704 30821 11713 30855
rect 11713 30821 11747 30855
rect 11747 30821 11756 30855
rect 11704 30812 11756 30821
rect 14280 30812 14332 30864
rect 11336 30744 11388 30796
rect 11428 30676 11480 30728
rect 18696 30880 18748 30932
rect 19616 30880 19668 30932
rect 20352 30880 20404 30932
rect 15936 30855 15988 30864
rect 15936 30821 15945 30855
rect 15945 30821 15979 30855
rect 15979 30821 15988 30855
rect 15936 30812 15988 30821
rect 17684 30812 17736 30864
rect 25320 30880 25372 30932
rect 15200 30744 15252 30796
rect 16488 30787 16540 30796
rect 16488 30753 16497 30787
rect 16497 30753 16531 30787
rect 16531 30753 16540 30787
rect 16488 30744 16540 30753
rect 19064 30744 19116 30796
rect 19892 30787 19944 30796
rect 19892 30753 19901 30787
rect 19901 30753 19935 30787
rect 19935 30753 19944 30787
rect 19892 30744 19944 30753
rect 19984 30787 20036 30796
rect 19984 30753 19993 30787
rect 19993 30753 20027 30787
rect 20027 30753 20036 30787
rect 19984 30744 20036 30753
rect 20536 30744 20588 30796
rect 15476 30676 15528 30728
rect 15936 30676 15988 30728
rect 3792 30608 3844 30660
rect 16120 30608 16172 30660
rect 20076 30676 20128 30728
rect 20444 30676 20496 30728
rect 22468 30719 22520 30728
rect 22468 30685 22477 30719
rect 22477 30685 22511 30719
rect 22511 30685 22520 30719
rect 22468 30676 22520 30685
rect 23848 30719 23900 30728
rect 23848 30685 23857 30719
rect 23857 30685 23891 30719
rect 23891 30685 23900 30719
rect 23848 30676 23900 30685
rect 25504 30676 25556 30728
rect 24492 30608 24544 30660
rect 8760 30540 8812 30592
rect 11336 30583 11388 30592
rect 11336 30549 11345 30583
rect 11345 30549 11379 30583
rect 11379 30549 11388 30583
rect 11336 30540 11388 30549
rect 14096 30540 14148 30592
rect 15384 30540 15436 30592
rect 17500 30540 17552 30592
rect 19432 30583 19484 30592
rect 19432 30549 19441 30583
rect 19441 30549 19475 30583
rect 19475 30549 19484 30583
rect 19432 30540 19484 30549
rect 21824 30540 21876 30592
rect 25136 30540 25188 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 10048 30379 10100 30388
rect 10048 30345 10057 30379
rect 10057 30345 10091 30379
rect 10091 30345 10100 30379
rect 10048 30336 10100 30345
rect 10324 30336 10376 30388
rect 6276 30268 6328 30320
rect 9588 30268 9640 30320
rect 11152 30132 11204 30184
rect 10416 30039 10468 30048
rect 10416 30005 10425 30039
rect 10425 30005 10459 30039
rect 10459 30005 10468 30039
rect 10416 29996 10468 30005
rect 11888 29996 11940 30048
rect 14372 30268 14424 30320
rect 15476 30268 15528 30320
rect 14464 30243 14516 30252
rect 14464 30209 14473 30243
rect 14473 30209 14507 30243
rect 14507 30209 14516 30243
rect 14464 30200 14516 30209
rect 16120 30336 16172 30388
rect 17960 30336 18012 30388
rect 18880 30336 18932 30388
rect 21088 30336 21140 30388
rect 23940 30336 23992 30388
rect 16304 30268 16356 30320
rect 18696 30200 18748 30252
rect 23572 30268 23624 30320
rect 22192 30200 22244 30252
rect 12440 30132 12492 30184
rect 12624 30132 12676 30184
rect 14832 30132 14884 30184
rect 16212 30175 16264 30184
rect 16212 30141 16221 30175
rect 16221 30141 16255 30175
rect 16255 30141 16264 30175
rect 16212 30132 16264 30141
rect 17224 30132 17276 30184
rect 18052 30175 18104 30184
rect 18052 30141 18061 30175
rect 18061 30141 18095 30175
rect 18095 30141 18104 30175
rect 18052 30132 18104 30141
rect 19524 30132 19576 30184
rect 23756 30132 23808 30184
rect 15844 30064 15896 30116
rect 17684 30064 17736 30116
rect 17960 30064 18012 30116
rect 18696 30064 18748 30116
rect 21640 30064 21692 30116
rect 12348 29996 12400 30048
rect 14464 29996 14516 30048
rect 17500 29996 17552 30048
rect 17592 30039 17644 30048
rect 17592 30005 17601 30039
rect 17601 30005 17635 30039
rect 17635 30005 17644 30039
rect 17592 29996 17644 30005
rect 21732 29996 21784 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 4252 29792 4304 29844
rect 7656 29792 7708 29844
rect 7748 29792 7800 29844
rect 9496 29835 9548 29844
rect 9496 29801 9505 29835
rect 9505 29801 9539 29835
rect 9539 29801 9548 29835
rect 9496 29792 9548 29801
rect 14464 29792 14516 29844
rect 11336 29724 11388 29776
rect 2688 29656 2740 29708
rect 7196 29656 7248 29708
rect 9128 29656 9180 29708
rect 7288 29588 7340 29640
rect 7840 29588 7892 29640
rect 14556 29724 14608 29776
rect 16028 29835 16080 29844
rect 16028 29801 16037 29835
rect 16037 29801 16071 29835
rect 16071 29801 16080 29835
rect 16028 29792 16080 29801
rect 16488 29792 16540 29844
rect 16580 29792 16632 29844
rect 18972 29792 19024 29844
rect 19800 29792 19852 29844
rect 16764 29724 16816 29776
rect 17592 29724 17644 29776
rect 14464 29656 14516 29708
rect 19064 29656 19116 29708
rect 21180 29656 21232 29708
rect 25688 29792 25740 29844
rect 21640 29724 21692 29776
rect 22836 29724 22888 29776
rect 24768 29724 24820 29776
rect 10416 29588 10468 29640
rect 14004 29588 14056 29640
rect 15292 29588 15344 29640
rect 16304 29588 16356 29640
rect 18052 29588 18104 29640
rect 18972 29588 19024 29640
rect 20812 29588 20864 29640
rect 22008 29588 22060 29640
rect 22560 29656 22612 29708
rect 23388 29699 23440 29708
rect 23388 29665 23397 29699
rect 23397 29665 23431 29699
rect 23431 29665 23440 29699
rect 23388 29656 23440 29665
rect 23756 29656 23808 29708
rect 22284 29588 22336 29640
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 3424 29520 3476 29572
rect 5264 29520 5316 29572
rect 7012 29520 7064 29572
rect 9312 29520 9364 29572
rect 9588 29520 9640 29572
rect 12348 29520 12400 29572
rect 12808 29520 12860 29572
rect 14740 29563 14792 29572
rect 14740 29529 14749 29563
rect 14749 29529 14783 29563
rect 14783 29529 14792 29563
rect 14740 29520 14792 29529
rect 7656 29452 7708 29504
rect 10048 29452 10100 29504
rect 10784 29452 10836 29504
rect 11888 29495 11940 29504
rect 11888 29461 11897 29495
rect 11897 29461 11931 29495
rect 11931 29461 11940 29495
rect 11888 29452 11940 29461
rect 12900 29452 12952 29504
rect 16580 29520 16632 29572
rect 17592 29520 17644 29572
rect 19340 29520 19392 29572
rect 15108 29452 15160 29504
rect 17500 29452 17552 29504
rect 18236 29452 18288 29504
rect 18420 29452 18472 29504
rect 18512 29495 18564 29504
rect 18512 29461 18521 29495
rect 18521 29461 18555 29495
rect 18555 29461 18564 29495
rect 18512 29452 18564 29461
rect 20352 29452 20404 29504
rect 20904 29495 20956 29504
rect 20904 29461 20913 29495
rect 20913 29461 20947 29495
rect 20947 29461 20956 29495
rect 20904 29452 20956 29461
rect 21456 29452 21508 29504
rect 23296 29495 23348 29504
rect 23296 29461 23305 29495
rect 23305 29461 23339 29495
rect 23339 29461 23348 29495
rect 23296 29452 23348 29461
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 7748 29248 7800 29300
rect 9496 29180 9548 29232
rect 12900 29291 12952 29300
rect 12900 29257 12909 29291
rect 12909 29257 12943 29291
rect 12943 29257 12952 29291
rect 12900 29248 12952 29257
rect 15568 29248 15620 29300
rect 6552 29044 6604 29096
rect 9404 29044 9456 29096
rect 10876 28976 10928 29028
rect 14004 29112 14056 29164
rect 14096 29155 14148 29164
rect 14096 29121 14105 29155
rect 14105 29121 14139 29155
rect 14139 29121 14148 29155
rect 14096 29112 14148 29121
rect 13544 29044 13596 29096
rect 13636 28976 13688 29028
rect 14648 29044 14700 29096
rect 15384 29087 15436 29096
rect 15384 29053 15393 29087
rect 15393 29053 15427 29087
rect 15427 29053 15436 29087
rect 15384 29044 15436 29053
rect 16396 29248 16448 29300
rect 17224 29291 17276 29300
rect 17224 29257 17233 29291
rect 17233 29257 17267 29291
rect 17267 29257 17276 29291
rect 17224 29248 17276 29257
rect 17500 29248 17552 29300
rect 17592 29248 17644 29300
rect 19800 29248 19852 29300
rect 20168 29248 20220 29300
rect 9680 28908 9732 28960
rect 15200 28908 15252 28960
rect 16028 28908 16080 28960
rect 18880 29180 18932 29232
rect 16764 29112 16816 29164
rect 20076 29180 20128 29232
rect 20536 29180 20588 29232
rect 20904 29248 20956 29300
rect 22836 29248 22888 29300
rect 25320 29291 25372 29300
rect 25320 29257 25329 29291
rect 25329 29257 25363 29291
rect 25363 29257 25372 29291
rect 25320 29248 25372 29257
rect 25504 29291 25556 29300
rect 25504 29257 25513 29291
rect 25513 29257 25547 29291
rect 25547 29257 25556 29291
rect 25504 29248 25556 29257
rect 17408 29087 17460 29096
rect 17408 29053 17417 29087
rect 17417 29053 17451 29087
rect 17451 29053 17460 29087
rect 17408 29044 17460 29053
rect 21548 29223 21600 29232
rect 21548 29189 21557 29223
rect 21557 29189 21591 29223
rect 21591 29189 21600 29223
rect 21548 29180 21600 29189
rect 24584 29180 24636 29232
rect 16396 29019 16448 29028
rect 16396 28985 16405 29019
rect 16405 28985 16439 29019
rect 16439 28985 16448 29019
rect 20168 29044 20220 29096
rect 22744 29112 22796 29164
rect 24124 29155 24176 29164
rect 24124 29121 24133 29155
rect 24133 29121 24167 29155
rect 24167 29121 24176 29155
rect 24124 29112 24176 29121
rect 16396 28976 16448 28985
rect 18512 28976 18564 29028
rect 22468 29044 22520 29096
rect 23572 29044 23624 29096
rect 23296 28976 23348 29028
rect 23388 28976 23440 29028
rect 16856 28951 16908 28960
rect 16856 28917 16865 28951
rect 16865 28917 16899 28951
rect 16899 28917 16908 28951
rect 16856 28908 16908 28917
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 8116 28704 8168 28756
rect 9496 28704 9548 28756
rect 14096 28704 14148 28756
rect 18788 28704 18840 28756
rect 18972 28704 19024 28756
rect 9864 28636 9916 28688
rect 16396 28636 16448 28688
rect 18328 28636 18380 28688
rect 21180 28747 21232 28756
rect 21180 28713 21189 28747
rect 21189 28713 21223 28747
rect 21223 28713 21232 28747
rect 21180 28704 21232 28713
rect 1308 28568 1360 28620
rect 4068 28568 4120 28620
rect 5172 28611 5224 28620
rect 5172 28577 5181 28611
rect 5181 28577 5215 28611
rect 5215 28577 5224 28611
rect 5172 28568 5224 28577
rect 6552 28611 6604 28620
rect 6552 28577 6561 28611
rect 6561 28577 6595 28611
rect 6595 28577 6604 28611
rect 6552 28568 6604 28577
rect 9404 28568 9456 28620
rect 11336 28568 11388 28620
rect 13360 28611 13412 28620
rect 13360 28577 13369 28611
rect 13369 28577 13403 28611
rect 13403 28577 13412 28611
rect 13360 28568 13412 28577
rect 14832 28611 14884 28620
rect 14832 28577 14841 28611
rect 14841 28577 14875 28611
rect 14875 28577 14884 28611
rect 14832 28568 14884 28577
rect 16212 28611 16264 28620
rect 16212 28577 16221 28611
rect 16221 28577 16255 28611
rect 16255 28577 16264 28611
rect 16212 28568 16264 28577
rect 17132 28568 17184 28620
rect 17776 28611 17828 28620
rect 17776 28577 17785 28611
rect 17785 28577 17819 28611
rect 17819 28577 17828 28611
rect 17776 28568 17828 28577
rect 22008 28568 22060 28620
rect 1768 28543 1820 28552
rect 1768 28509 1777 28543
rect 1777 28509 1811 28543
rect 1811 28509 1820 28543
rect 1768 28500 1820 28509
rect 9956 28500 10008 28552
rect 15200 28500 15252 28552
rect 16856 28500 16908 28552
rect 17868 28500 17920 28552
rect 3976 28364 4028 28416
rect 8116 28432 8168 28484
rect 12532 28432 12584 28484
rect 13360 28432 13412 28484
rect 15476 28432 15528 28484
rect 16672 28432 16724 28484
rect 19616 28432 19668 28484
rect 22192 28432 22244 28484
rect 24768 28543 24820 28552
rect 24768 28509 24777 28543
rect 24777 28509 24811 28543
rect 24811 28509 24820 28543
rect 24768 28500 24820 28509
rect 24216 28432 24268 28484
rect 24860 28432 24912 28484
rect 12808 28364 12860 28416
rect 13176 28407 13228 28416
rect 13176 28373 13185 28407
rect 13185 28373 13219 28407
rect 13219 28373 13228 28407
rect 13176 28364 13228 28373
rect 13268 28407 13320 28416
rect 13268 28373 13277 28407
rect 13277 28373 13311 28407
rect 13311 28373 13320 28407
rect 13268 28364 13320 28373
rect 14004 28364 14056 28416
rect 14280 28407 14332 28416
rect 14280 28373 14289 28407
rect 14289 28373 14323 28407
rect 14323 28373 14332 28407
rect 14280 28364 14332 28373
rect 14924 28364 14976 28416
rect 15292 28407 15344 28416
rect 15292 28373 15301 28407
rect 15301 28373 15335 28407
rect 15335 28373 15344 28407
rect 15292 28364 15344 28373
rect 15752 28364 15804 28416
rect 16764 28407 16816 28416
rect 16764 28373 16773 28407
rect 16773 28373 16807 28407
rect 16807 28373 16816 28407
rect 16764 28364 16816 28373
rect 16948 28364 17000 28416
rect 24584 28407 24636 28416
rect 24584 28373 24593 28407
rect 24593 28373 24627 28407
rect 24627 28373 24636 28407
rect 24584 28364 24636 28373
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 1952 28160 2004 28212
rect 3792 28160 3844 28212
rect 13176 28160 13228 28212
rect 13360 28203 13412 28212
rect 13360 28169 13369 28203
rect 13369 28169 13403 28203
rect 13403 28169 13412 28203
rect 13360 28160 13412 28169
rect 15476 28160 15528 28212
rect 15936 28203 15988 28212
rect 15936 28169 15945 28203
rect 15945 28169 15979 28203
rect 15979 28169 15988 28203
rect 15936 28160 15988 28169
rect 18328 28203 18380 28212
rect 18328 28169 18337 28203
rect 18337 28169 18371 28203
rect 18371 28169 18380 28203
rect 18328 28160 18380 28169
rect 19064 28160 19116 28212
rect 16396 28092 16448 28144
rect 3332 28024 3384 28076
rect 3608 28067 3660 28076
rect 3608 28033 3652 28067
rect 3652 28033 3660 28067
rect 3608 28024 3660 28033
rect 8576 27999 8628 28008
rect 8576 27965 8585 27999
rect 8585 27965 8619 27999
rect 8619 27965 8628 27999
rect 8576 27956 8628 27965
rect 9680 27888 9732 27940
rect 10600 27888 10652 27940
rect 13268 28024 13320 28076
rect 15936 28024 15988 28076
rect 16028 27999 16080 28008
rect 16028 27965 16037 27999
rect 16037 27965 16071 27999
rect 16071 27965 16080 27999
rect 16028 27956 16080 27965
rect 21088 28092 21140 28144
rect 22192 28092 22244 28144
rect 24676 28135 24728 28144
rect 24676 28101 24685 28135
rect 24685 28101 24719 28135
rect 24719 28101 24728 28135
rect 24676 28092 24728 28101
rect 9956 27820 10008 27872
rect 10692 27820 10744 27872
rect 14924 27820 14976 27872
rect 15568 27863 15620 27872
rect 15568 27829 15577 27863
rect 15577 27829 15611 27863
rect 15611 27829 15620 27863
rect 15568 27820 15620 27829
rect 15844 27820 15896 27872
rect 19340 28024 19392 28076
rect 22008 28067 22060 28076
rect 22008 28033 22017 28067
rect 22017 28033 22051 28067
rect 22051 28033 22060 28067
rect 22008 28024 22060 28033
rect 18604 27956 18656 28008
rect 18788 27956 18840 28008
rect 17868 27863 17920 27872
rect 17868 27829 17877 27863
rect 17877 27829 17911 27863
rect 17911 27829 17920 27863
rect 17868 27820 17920 27829
rect 19064 27863 19116 27872
rect 19064 27829 19073 27863
rect 19073 27829 19107 27863
rect 19107 27829 19116 27863
rect 19064 27820 19116 27829
rect 19984 27956 20036 28008
rect 24676 27956 24728 28008
rect 20076 27863 20128 27872
rect 20076 27829 20085 27863
rect 20085 27829 20119 27863
rect 20119 27829 20128 27863
rect 20076 27820 20128 27829
rect 22744 27820 22796 27872
rect 23388 27820 23440 27872
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 9864 27616 9916 27668
rect 12532 27616 12584 27668
rect 13268 27616 13320 27668
rect 18328 27616 18380 27668
rect 18604 27616 18656 27668
rect 21640 27616 21692 27668
rect 22192 27616 22244 27668
rect 22836 27616 22888 27668
rect 23388 27616 23440 27668
rect 24216 27659 24268 27668
rect 24216 27625 24225 27659
rect 24225 27625 24259 27659
rect 24259 27625 24268 27659
rect 24216 27616 24268 27625
rect 7840 27548 7892 27600
rect 8300 27591 8352 27600
rect 8300 27557 8309 27591
rect 8309 27557 8343 27591
rect 8343 27557 8352 27591
rect 8300 27548 8352 27557
rect 21548 27548 21600 27600
rect 6552 27480 6604 27532
rect 9956 27412 10008 27464
rect 12072 27480 12124 27532
rect 12808 27480 12860 27532
rect 12532 27412 12584 27464
rect 15844 27412 15896 27464
rect 17684 27412 17736 27464
rect 20444 27480 20496 27532
rect 20628 27523 20680 27532
rect 20628 27489 20637 27523
rect 20637 27489 20671 27523
rect 20671 27489 20680 27523
rect 20628 27480 20680 27489
rect 21916 27523 21968 27532
rect 21916 27489 21925 27523
rect 21925 27489 21959 27523
rect 21959 27489 21968 27523
rect 21916 27480 21968 27489
rect 22652 27480 22704 27532
rect 21272 27412 21324 27464
rect 8300 27344 8352 27396
rect 11428 27387 11480 27396
rect 11428 27353 11437 27387
rect 11437 27353 11471 27387
rect 11471 27353 11480 27387
rect 11428 27344 11480 27353
rect 15384 27344 15436 27396
rect 10232 27276 10284 27328
rect 12900 27319 12952 27328
rect 12900 27285 12909 27319
rect 12909 27285 12943 27319
rect 12943 27285 12952 27319
rect 12900 27276 12952 27285
rect 15016 27276 15068 27328
rect 17224 27344 17276 27396
rect 17132 27276 17184 27328
rect 19340 27276 19392 27328
rect 22100 27344 22152 27396
rect 22192 27387 22244 27396
rect 22192 27353 22201 27387
rect 22201 27353 22235 27387
rect 22235 27353 22244 27387
rect 22192 27344 22244 27353
rect 22836 27344 22888 27396
rect 25596 27344 25648 27396
rect 23112 27276 23164 27328
rect 25228 27319 25280 27328
rect 25228 27285 25237 27319
rect 25237 27285 25271 27319
rect 25271 27285 25280 27319
rect 25228 27276 25280 27285
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 3424 27072 3476 27124
rect 10692 27072 10744 27124
rect 1584 27004 1636 27056
rect 4344 27004 4396 27056
rect 8116 27004 8168 27056
rect 8300 27004 8352 27056
rect 11244 27004 11296 27056
rect 3424 26936 3476 26988
rect 6552 26979 6604 26988
rect 6552 26945 6561 26979
rect 6561 26945 6595 26979
rect 6595 26945 6604 26979
rect 6552 26936 6604 26945
rect 9128 26979 9180 26988
rect 9128 26945 9137 26979
rect 9137 26945 9171 26979
rect 9171 26945 9180 26979
rect 9128 26936 9180 26945
rect 7840 26868 7892 26920
rect 8668 26868 8720 26920
rect 9404 26911 9456 26920
rect 9404 26877 9413 26911
rect 9413 26877 9447 26911
rect 9447 26877 9456 26911
rect 9404 26868 9456 26877
rect 4528 26800 4580 26852
rect 8300 26843 8352 26852
rect 8300 26809 8309 26843
rect 8309 26809 8343 26843
rect 8343 26809 8352 26843
rect 8300 26800 8352 26809
rect 9680 26800 9732 26852
rect 10140 26800 10192 26852
rect 12900 27072 12952 27124
rect 12072 27004 12124 27056
rect 12808 27047 12860 27056
rect 12808 27013 12817 27047
rect 12817 27013 12851 27047
rect 12851 27013 12860 27047
rect 12808 27004 12860 27013
rect 13268 27004 13320 27056
rect 15108 27072 15160 27124
rect 20168 27072 20220 27124
rect 20444 27072 20496 27124
rect 14188 26936 14240 26988
rect 18972 27004 19024 27056
rect 24584 27072 24636 27124
rect 23112 27047 23164 27056
rect 23112 27013 23121 27047
rect 23121 27013 23155 27047
rect 23155 27013 23164 27047
rect 23112 27004 23164 27013
rect 23388 27004 23440 27056
rect 25136 27047 25188 27056
rect 25136 27013 25145 27047
rect 25145 27013 25179 27047
rect 25179 27013 25188 27047
rect 25136 27004 25188 27013
rect 12532 26800 12584 26852
rect 10508 26732 10560 26784
rect 10600 26732 10652 26784
rect 12348 26732 12400 26784
rect 14372 26732 14424 26784
rect 14740 26775 14792 26784
rect 14740 26741 14749 26775
rect 14749 26741 14783 26775
rect 14783 26741 14792 26775
rect 14740 26732 14792 26741
rect 19340 26868 19392 26920
rect 19524 26868 19576 26920
rect 21180 26868 21232 26920
rect 22008 26868 22060 26920
rect 20628 26800 20680 26852
rect 23112 26868 23164 26920
rect 23480 26868 23532 26920
rect 25412 26800 25464 26852
rect 18328 26732 18380 26784
rect 19524 26775 19576 26784
rect 19524 26741 19533 26775
rect 19533 26741 19567 26775
rect 19567 26741 19576 26775
rect 19524 26732 19576 26741
rect 23848 26732 23900 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 4068 26571 4120 26580
rect 4068 26537 4077 26571
rect 4077 26537 4111 26571
rect 4111 26537 4120 26571
rect 4068 26528 4120 26537
rect 7104 26528 7156 26580
rect 7748 26528 7800 26580
rect 9220 26528 9272 26580
rect 6460 26435 6512 26444
rect 6460 26401 6469 26435
rect 6469 26401 6503 26435
rect 6503 26401 6512 26435
rect 6460 26392 6512 26401
rect 8300 26392 8352 26444
rect 9128 26435 9180 26444
rect 9128 26401 9137 26435
rect 9137 26401 9171 26435
rect 9171 26401 9180 26435
rect 9128 26392 9180 26401
rect 10232 26435 10284 26444
rect 10232 26401 10241 26435
rect 10241 26401 10275 26435
rect 10275 26401 10284 26435
rect 10232 26392 10284 26401
rect 2044 26324 2096 26376
rect 9956 26367 10008 26376
rect 9956 26333 9965 26367
rect 9965 26333 9999 26367
rect 9999 26333 10008 26367
rect 9956 26324 10008 26333
rect 12532 26528 12584 26580
rect 14648 26528 14700 26580
rect 16672 26528 16724 26580
rect 17776 26528 17828 26580
rect 21916 26528 21968 26580
rect 12256 26460 12308 26512
rect 12348 26460 12400 26512
rect 19708 26460 19760 26512
rect 22008 26460 22060 26512
rect 22192 26460 22244 26512
rect 22560 26460 22612 26512
rect 17040 26392 17092 26444
rect 14280 26324 14332 26376
rect 15384 26367 15436 26376
rect 15384 26333 15393 26367
rect 15393 26333 15427 26367
rect 15427 26333 15436 26367
rect 15384 26324 15436 26333
rect 2780 26299 2832 26308
rect 2780 26265 2789 26299
rect 2789 26265 2823 26299
rect 2823 26265 2832 26299
rect 2780 26256 2832 26265
rect 8116 26256 8168 26308
rect 8484 26256 8536 26308
rect 8668 26299 8720 26308
rect 8668 26265 8677 26299
rect 8677 26265 8711 26299
rect 8711 26265 8720 26299
rect 8668 26256 8720 26265
rect 9588 26256 9640 26308
rect 10692 26256 10744 26308
rect 14832 26256 14884 26308
rect 17868 26392 17920 26444
rect 20168 26392 20220 26444
rect 20260 26324 20312 26376
rect 23572 26528 23624 26580
rect 25044 26528 25096 26580
rect 25228 26528 25280 26580
rect 24492 26392 24544 26444
rect 24400 26324 24452 26376
rect 14648 26188 14700 26240
rect 17684 26256 17736 26308
rect 21180 26256 21232 26308
rect 21640 26256 21692 26308
rect 22468 26256 22520 26308
rect 25228 26256 25280 26308
rect 17592 26231 17644 26240
rect 17592 26197 17601 26231
rect 17601 26197 17635 26231
rect 17635 26197 17644 26231
rect 17592 26188 17644 26197
rect 22652 26188 22704 26240
rect 23388 26188 23440 26240
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 1768 25984 1820 26036
rect 6736 25984 6788 26036
rect 8852 25984 8904 26036
rect 9220 26027 9272 26036
rect 9220 25993 9229 26027
rect 9229 25993 9263 26027
rect 9263 25993 9272 26027
rect 9220 25984 9272 25993
rect 10508 25984 10560 26036
rect 10876 26027 10928 26036
rect 10876 25993 10885 26027
rect 10885 25993 10919 26027
rect 10919 25993 10928 26027
rect 10876 25984 10928 25993
rect 3516 25916 3568 25968
rect 4068 25916 4120 25968
rect 2872 25848 2924 25900
rect 8484 25959 8536 25968
rect 8484 25925 8493 25959
rect 8493 25925 8527 25959
rect 8527 25925 8536 25959
rect 8484 25916 8536 25925
rect 9772 25916 9824 25968
rect 10692 25916 10744 25968
rect 2780 25780 2832 25832
rect 3608 25780 3660 25832
rect 9404 25848 9456 25900
rect 15384 25984 15436 26036
rect 15568 25984 15620 26036
rect 17592 25984 17644 26036
rect 14648 25916 14700 25968
rect 19340 26027 19392 26036
rect 19340 25993 19349 26027
rect 19349 25993 19383 26027
rect 19383 25993 19392 26027
rect 19340 25984 19392 25993
rect 19524 25984 19576 26036
rect 20352 26027 20404 26036
rect 20352 25993 20361 26027
rect 20361 25993 20395 26027
rect 20395 25993 20404 26027
rect 20352 25984 20404 25993
rect 22376 25984 22428 26036
rect 21364 25916 21416 25968
rect 6184 25780 6236 25832
rect 7840 25780 7892 25832
rect 3332 25712 3384 25764
rect 4252 25687 4304 25696
rect 4252 25653 4261 25687
rect 4261 25653 4295 25687
rect 4295 25653 4304 25687
rect 4252 25644 4304 25653
rect 5448 25644 5500 25696
rect 8760 25780 8812 25832
rect 8576 25712 8628 25764
rect 9588 25712 9640 25764
rect 9864 25780 9916 25832
rect 11796 25780 11848 25832
rect 14372 25780 14424 25832
rect 14464 25823 14516 25832
rect 14464 25789 14473 25823
rect 14473 25789 14507 25823
rect 14507 25789 14516 25823
rect 14464 25780 14516 25789
rect 12348 25644 12400 25696
rect 15108 25644 15160 25696
rect 16028 25823 16080 25832
rect 16028 25789 16037 25823
rect 16037 25789 16071 25823
rect 16071 25789 16080 25823
rect 16028 25780 16080 25789
rect 17868 25823 17920 25832
rect 17868 25789 17877 25823
rect 17877 25789 17911 25823
rect 17911 25789 17920 25823
rect 17868 25780 17920 25789
rect 22192 25848 22244 25900
rect 22284 25848 22336 25900
rect 23388 25848 23440 25900
rect 23848 25848 23900 25900
rect 21272 25823 21324 25832
rect 21272 25789 21281 25823
rect 21281 25789 21315 25823
rect 21315 25789 21324 25823
rect 21272 25780 21324 25789
rect 22284 25712 22336 25764
rect 25136 25823 25188 25832
rect 25136 25789 25145 25823
rect 25145 25789 25179 25823
rect 25179 25789 25188 25823
rect 25136 25780 25188 25789
rect 24400 25712 24452 25764
rect 18420 25644 18472 25696
rect 18880 25644 18932 25696
rect 21364 25644 21416 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 14188 25440 14240 25492
rect 16764 25440 16816 25492
rect 17592 25440 17644 25492
rect 17776 25440 17828 25492
rect 22376 25440 22428 25492
rect 23388 25483 23440 25492
rect 23388 25449 23397 25483
rect 23397 25449 23431 25483
rect 23431 25449 23440 25483
rect 23388 25440 23440 25449
rect 24860 25440 24912 25492
rect 25044 25440 25096 25492
rect 25504 25483 25556 25492
rect 25504 25449 25513 25483
rect 25513 25449 25547 25483
rect 25547 25449 25556 25483
rect 25504 25440 25556 25449
rect 7656 25304 7708 25356
rect 9404 25347 9456 25356
rect 9404 25313 9413 25347
rect 9413 25313 9447 25347
rect 9447 25313 9456 25347
rect 9404 25304 9456 25313
rect 9680 25304 9732 25356
rect 11428 25304 11480 25356
rect 14464 25372 14516 25424
rect 12808 25304 12860 25356
rect 13820 25304 13872 25356
rect 14188 25304 14240 25356
rect 15384 25304 15436 25356
rect 24952 25372 25004 25424
rect 16672 25304 16724 25356
rect 19064 25304 19116 25356
rect 20076 25347 20128 25356
rect 20076 25313 20085 25347
rect 20085 25313 20119 25347
rect 20119 25313 20128 25347
rect 20076 25304 20128 25313
rect 22652 25347 22704 25356
rect 22652 25313 22661 25347
rect 22661 25313 22695 25347
rect 22695 25313 22704 25347
rect 22652 25304 22704 25313
rect 4068 25279 4120 25288
rect 4068 25245 4086 25279
rect 4086 25245 4120 25279
rect 4068 25236 4120 25245
rect 8392 25236 8444 25288
rect 10784 25236 10836 25288
rect 11796 25279 11848 25288
rect 11796 25245 11805 25279
rect 11805 25245 11839 25279
rect 11839 25245 11848 25279
rect 11796 25236 11848 25245
rect 12624 25236 12676 25288
rect 19432 25236 19484 25288
rect 21272 25236 21324 25288
rect 24032 25236 24084 25288
rect 24308 25236 24360 25288
rect 7104 25211 7156 25220
rect 7104 25177 7113 25211
rect 7113 25177 7147 25211
rect 7147 25177 7156 25211
rect 7104 25168 7156 25177
rect 9772 25168 9824 25220
rect 3976 25100 4028 25152
rect 8576 25143 8628 25152
rect 8576 25109 8585 25143
rect 8585 25109 8619 25143
rect 8619 25109 8628 25143
rect 8576 25100 8628 25109
rect 13452 25168 13504 25220
rect 14648 25168 14700 25220
rect 22100 25168 22152 25220
rect 25044 25168 25096 25220
rect 11152 25143 11204 25152
rect 11152 25109 11161 25143
rect 11161 25109 11195 25143
rect 11195 25109 11204 25143
rect 11152 25100 11204 25109
rect 11980 25100 12032 25152
rect 12624 25143 12676 25152
rect 12624 25109 12633 25143
rect 12633 25109 12667 25143
rect 12667 25109 12676 25143
rect 12624 25100 12676 25109
rect 12808 25100 12860 25152
rect 14924 25100 14976 25152
rect 16856 25100 16908 25152
rect 17040 25100 17092 25152
rect 17868 25100 17920 25152
rect 18328 25100 18380 25152
rect 19524 25100 19576 25152
rect 23940 25143 23992 25152
rect 23940 25109 23949 25143
rect 23949 25109 23983 25143
rect 23983 25109 23992 25143
rect 23940 25100 23992 25109
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 4252 24896 4304 24948
rect 7840 24896 7892 24948
rect 9496 24896 9548 24948
rect 11152 24896 11204 24948
rect 12624 24896 12676 24948
rect 16856 24939 16908 24948
rect 16856 24905 16865 24939
rect 16865 24905 16899 24939
rect 16899 24905 16908 24939
rect 16856 24896 16908 24905
rect 7104 24828 7156 24880
rect 6000 24692 6052 24744
rect 3976 24556 4028 24608
rect 7564 24760 7616 24812
rect 7748 24760 7800 24812
rect 12992 24828 13044 24880
rect 17224 24871 17276 24880
rect 17224 24837 17233 24871
rect 17233 24837 17267 24871
rect 17267 24837 17276 24871
rect 17224 24828 17276 24837
rect 8116 24735 8168 24744
rect 8116 24701 8125 24735
rect 8125 24701 8159 24735
rect 8159 24701 8168 24735
rect 8116 24692 8168 24701
rect 9312 24735 9364 24744
rect 9312 24701 9321 24735
rect 9321 24701 9355 24735
rect 9355 24701 9364 24735
rect 9312 24692 9364 24701
rect 12440 24760 12492 24812
rect 12624 24760 12676 24812
rect 13268 24760 13320 24812
rect 13820 24803 13872 24812
rect 13820 24769 13829 24803
rect 13829 24769 13863 24803
rect 13863 24769 13872 24803
rect 13820 24760 13872 24769
rect 9680 24692 9732 24744
rect 8392 24624 8444 24676
rect 6920 24556 6972 24608
rect 7472 24556 7524 24608
rect 11152 24556 11204 24608
rect 12072 24556 12124 24608
rect 12532 24692 12584 24744
rect 14648 24760 14700 24812
rect 15016 24760 15068 24812
rect 16856 24760 16908 24812
rect 18328 24828 18380 24880
rect 18512 24828 18564 24880
rect 22652 24828 22704 24880
rect 14372 24692 14424 24744
rect 14924 24624 14976 24676
rect 17684 24760 17736 24812
rect 17868 24760 17920 24812
rect 19892 24760 19944 24812
rect 17592 24692 17644 24744
rect 18788 24692 18840 24744
rect 19248 24692 19300 24744
rect 22008 24760 22060 24812
rect 22100 24760 22152 24812
rect 24308 24760 24360 24812
rect 24860 24760 24912 24812
rect 25504 24760 25556 24812
rect 12992 24599 13044 24608
rect 12992 24565 13001 24599
rect 13001 24565 13035 24599
rect 13035 24565 13044 24599
rect 12992 24556 13044 24565
rect 13728 24556 13780 24608
rect 14648 24556 14700 24608
rect 18696 24624 18748 24676
rect 20536 24624 20588 24676
rect 22836 24692 22888 24744
rect 22100 24624 22152 24676
rect 24676 24735 24728 24744
rect 24676 24701 24685 24735
rect 24685 24701 24719 24735
rect 24719 24701 24728 24735
rect 24676 24692 24728 24701
rect 16856 24556 16908 24608
rect 17316 24556 17368 24608
rect 18512 24556 18564 24608
rect 19892 24599 19944 24608
rect 19892 24565 19901 24599
rect 19901 24565 19935 24599
rect 19935 24565 19944 24599
rect 19892 24556 19944 24565
rect 24584 24556 24636 24608
rect 24768 24556 24820 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 3424 24395 3476 24404
rect 3424 24361 3433 24395
rect 3433 24361 3467 24395
rect 3467 24361 3476 24395
rect 3424 24352 3476 24361
rect 4436 24352 4488 24404
rect 6184 24395 6236 24404
rect 6184 24361 6193 24395
rect 6193 24361 6227 24395
rect 6227 24361 6236 24395
rect 6184 24352 6236 24361
rect 8760 24395 8812 24404
rect 8760 24361 8769 24395
rect 8769 24361 8803 24395
rect 8803 24361 8812 24395
rect 8760 24352 8812 24361
rect 9312 24352 9364 24404
rect 10324 24352 10376 24404
rect 6368 24284 6420 24336
rect 8576 24284 8628 24336
rect 4252 24259 4304 24268
rect 4252 24225 4261 24259
rect 4261 24225 4295 24259
rect 4295 24225 4304 24259
rect 4252 24216 4304 24225
rect 9864 24216 9916 24268
rect 10416 24216 10468 24268
rect 2780 24148 2832 24200
rect 3516 24148 3568 24200
rect 3976 24191 4028 24200
rect 3976 24157 3985 24191
rect 3985 24157 4019 24191
rect 4019 24157 4028 24191
rect 3976 24148 4028 24157
rect 7104 24148 7156 24200
rect 4252 24080 4304 24132
rect 1860 24012 1912 24064
rect 11060 24216 11112 24268
rect 12532 24352 12584 24404
rect 13360 24352 13412 24404
rect 12808 24216 12860 24268
rect 11152 24191 11204 24200
rect 11152 24157 11161 24191
rect 11161 24157 11195 24191
rect 11195 24157 11204 24191
rect 11152 24148 11204 24157
rect 13544 24148 13596 24200
rect 11520 24080 11572 24132
rect 11796 24080 11848 24132
rect 6920 24012 6972 24064
rect 7840 24012 7892 24064
rect 8484 24012 8536 24064
rect 9312 24012 9364 24064
rect 9404 24055 9456 24064
rect 9404 24021 9413 24055
rect 9413 24021 9447 24055
rect 9447 24021 9456 24055
rect 9404 24012 9456 24021
rect 9772 24055 9824 24064
rect 9772 24021 9781 24055
rect 9781 24021 9815 24055
rect 9815 24021 9824 24055
rect 9772 24012 9824 24021
rect 10784 24055 10836 24064
rect 10784 24021 10793 24055
rect 10793 24021 10827 24055
rect 10827 24021 10836 24055
rect 10784 24012 10836 24021
rect 11980 24055 12032 24064
rect 11980 24021 11989 24055
rect 11989 24021 12023 24055
rect 12023 24021 12032 24055
rect 11980 24012 12032 24021
rect 15200 24352 15252 24404
rect 15660 24352 15712 24404
rect 17592 24352 17644 24404
rect 21824 24352 21876 24404
rect 24676 24352 24728 24404
rect 14648 24284 14700 24336
rect 17684 24284 17736 24336
rect 18696 24284 18748 24336
rect 13820 24216 13872 24268
rect 16948 24216 17000 24268
rect 17040 24259 17092 24268
rect 17040 24225 17049 24259
rect 17049 24225 17083 24259
rect 17083 24225 17092 24259
rect 17040 24216 17092 24225
rect 22100 24216 22152 24268
rect 16764 24191 16816 24200
rect 16764 24157 16773 24191
rect 16773 24157 16807 24191
rect 16807 24157 16816 24191
rect 16764 24148 16816 24157
rect 14556 24080 14608 24132
rect 21732 24148 21784 24200
rect 24768 24284 24820 24336
rect 24860 24216 24912 24268
rect 18788 24080 18840 24132
rect 19248 24080 19300 24132
rect 21640 24080 21692 24132
rect 21824 24080 21876 24132
rect 23296 24148 23348 24200
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 25688 24148 25740 24200
rect 22192 24123 22244 24132
rect 22192 24089 22201 24123
rect 22201 24089 22235 24123
rect 22235 24089 22244 24123
rect 22192 24080 22244 24089
rect 17132 24012 17184 24064
rect 17408 24012 17460 24064
rect 17684 24012 17736 24064
rect 19432 24012 19484 24064
rect 20260 24012 20312 24064
rect 23572 24012 23624 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 6000 23851 6052 23860
rect 6000 23817 6009 23851
rect 6009 23817 6043 23851
rect 6043 23817 6052 23851
rect 6000 23808 6052 23817
rect 6828 23808 6880 23860
rect 9680 23808 9732 23860
rect 9772 23808 9824 23860
rect 10784 23808 10836 23860
rect 14832 23808 14884 23860
rect 19248 23808 19300 23860
rect 4160 23740 4212 23792
rect 4436 23740 4488 23792
rect 6920 23740 6972 23792
rect 8484 23740 8536 23792
rect 9312 23740 9364 23792
rect 11796 23783 11848 23792
rect 11796 23749 11805 23783
rect 11805 23749 11839 23783
rect 11839 23749 11848 23783
rect 11796 23740 11848 23749
rect 11888 23740 11940 23792
rect 17868 23740 17920 23792
rect 1768 23715 1820 23724
rect 1768 23681 1777 23715
rect 1777 23681 1811 23715
rect 1811 23681 1820 23715
rect 1768 23672 1820 23681
rect 9864 23672 9916 23724
rect 12164 23672 12216 23724
rect 1308 23604 1360 23656
rect 3976 23604 4028 23656
rect 7564 23604 7616 23656
rect 7656 23647 7708 23656
rect 7656 23613 7665 23647
rect 7665 23613 7699 23647
rect 7699 23613 7708 23647
rect 7656 23604 7708 23613
rect 8576 23604 8628 23656
rect 11704 23604 11756 23656
rect 12624 23604 12676 23656
rect 13728 23672 13780 23724
rect 17224 23672 17276 23724
rect 14372 23604 14424 23656
rect 14924 23604 14976 23656
rect 17040 23647 17092 23656
rect 17040 23613 17049 23647
rect 17049 23613 17083 23647
rect 17083 23613 17092 23647
rect 17040 23604 17092 23613
rect 5724 23468 5776 23520
rect 9956 23468 10008 23520
rect 10968 23468 11020 23520
rect 16488 23536 16540 23588
rect 12164 23511 12216 23520
rect 12164 23477 12173 23511
rect 12173 23477 12207 23511
rect 12207 23477 12216 23511
rect 12164 23468 12216 23477
rect 12440 23468 12492 23520
rect 13728 23468 13780 23520
rect 13912 23511 13964 23520
rect 13912 23477 13921 23511
rect 13921 23477 13955 23511
rect 13955 23477 13964 23511
rect 18972 23740 19024 23792
rect 19340 23740 19392 23792
rect 21640 23851 21692 23860
rect 21640 23817 21649 23851
rect 21649 23817 21683 23851
rect 21683 23817 21692 23851
rect 21640 23808 21692 23817
rect 22836 23808 22888 23860
rect 20536 23740 20588 23792
rect 23204 23740 23256 23792
rect 18604 23604 18656 23656
rect 19064 23647 19116 23656
rect 19064 23613 19073 23647
rect 19073 23613 19107 23647
rect 19107 23613 19116 23647
rect 19064 23604 19116 23613
rect 19432 23604 19484 23656
rect 22008 23672 22060 23724
rect 22100 23672 22152 23724
rect 13912 23468 13964 23477
rect 21088 23511 21140 23520
rect 21088 23477 21097 23511
rect 21097 23477 21131 23511
rect 21131 23477 21140 23511
rect 21088 23468 21140 23477
rect 24308 23672 24360 23724
rect 25320 23715 25372 23724
rect 25320 23681 25329 23715
rect 25329 23681 25363 23715
rect 25363 23681 25372 23715
rect 25320 23672 25372 23681
rect 23204 23647 23256 23656
rect 23204 23613 23213 23647
rect 23213 23613 23247 23647
rect 23247 23613 23256 23647
rect 23204 23604 23256 23613
rect 23664 23604 23716 23656
rect 24492 23604 24544 23656
rect 24216 23468 24268 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 2044 23307 2096 23316
rect 2044 23273 2053 23307
rect 2053 23273 2087 23307
rect 2087 23273 2096 23307
rect 2044 23264 2096 23273
rect 2872 23264 2924 23316
rect 3884 23264 3936 23316
rect 7564 23307 7616 23316
rect 7564 23273 7573 23307
rect 7573 23273 7607 23307
rect 7607 23273 7616 23307
rect 7564 23264 7616 23273
rect 12624 23264 12676 23316
rect 12808 23264 12860 23316
rect 14556 23264 14608 23316
rect 16028 23307 16080 23316
rect 16028 23273 16037 23307
rect 16037 23273 16071 23307
rect 16071 23273 16080 23307
rect 16028 23264 16080 23273
rect 16396 23264 16448 23316
rect 17776 23264 17828 23316
rect 19340 23264 19392 23316
rect 20076 23264 20128 23316
rect 20444 23264 20496 23316
rect 7840 23239 7892 23248
rect 7840 23205 7849 23239
rect 7849 23205 7883 23239
rect 7883 23205 7892 23239
rect 7840 23196 7892 23205
rect 9772 23196 9824 23248
rect 12440 23196 12492 23248
rect 24492 23196 24544 23248
rect 2872 23128 2924 23180
rect 3424 23128 3476 23180
rect 5080 23128 5132 23180
rect 5724 23128 5776 23180
rect 6460 23128 6512 23180
rect 3700 23060 3752 23112
rect 4344 23060 4396 23112
rect 7380 23128 7432 23180
rect 10048 23128 10100 23180
rect 10784 23128 10836 23180
rect 11612 23128 11664 23180
rect 12624 23128 12676 23180
rect 14280 23171 14332 23180
rect 14280 23137 14289 23171
rect 14289 23137 14323 23171
rect 14323 23137 14332 23171
rect 14280 23128 14332 23137
rect 15292 23128 15344 23180
rect 18604 23128 18656 23180
rect 10968 23060 11020 23112
rect 11704 23103 11756 23112
rect 11704 23069 11713 23103
rect 11713 23069 11747 23103
rect 11747 23069 11756 23103
rect 11704 23060 11756 23069
rect 12164 23060 12216 23112
rect 13912 23060 13964 23112
rect 16120 23060 16172 23112
rect 16396 23060 16448 23112
rect 23848 23171 23900 23180
rect 23848 23137 23857 23171
rect 23857 23137 23891 23171
rect 23891 23137 23900 23171
rect 23848 23128 23900 23137
rect 24584 23128 24636 23180
rect 3792 22992 3844 23044
rect 7748 22992 7800 23044
rect 9956 22924 10008 22976
rect 10784 22992 10836 23044
rect 12624 22967 12676 22976
rect 12624 22933 12633 22967
rect 12633 22933 12667 22967
rect 12667 22933 12676 22967
rect 12624 22924 12676 22933
rect 13084 22924 13136 22976
rect 15936 22992 15988 23044
rect 17776 22992 17828 23044
rect 15384 22924 15436 22976
rect 15476 22924 15528 22976
rect 15844 22924 15896 22976
rect 16212 22924 16264 22976
rect 16488 22924 16540 22976
rect 19984 22992 20036 23044
rect 19340 22924 19392 22976
rect 25412 22992 25464 23044
rect 21088 22924 21140 22976
rect 22836 22924 22888 22976
rect 23480 22924 23532 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 1768 22720 1820 22772
rect 9404 22720 9456 22772
rect 10048 22720 10100 22772
rect 12072 22720 12124 22772
rect 12808 22720 12860 22772
rect 13084 22763 13136 22772
rect 13084 22729 13093 22763
rect 13093 22729 13127 22763
rect 13127 22729 13136 22763
rect 13084 22720 13136 22729
rect 15108 22720 15160 22772
rect 15384 22720 15436 22772
rect 16028 22720 16080 22772
rect 11520 22652 11572 22704
rect 11888 22652 11940 22704
rect 2872 22584 2924 22636
rect 7840 22584 7892 22636
rect 9680 22584 9732 22636
rect 15292 22652 15344 22704
rect 16120 22652 16172 22704
rect 6000 22516 6052 22568
rect 7288 22559 7340 22568
rect 7288 22525 7297 22559
rect 7297 22525 7331 22559
rect 7331 22525 7340 22559
rect 7288 22516 7340 22525
rect 7564 22516 7616 22568
rect 8852 22559 8904 22568
rect 8852 22525 8861 22559
rect 8861 22525 8895 22559
rect 8895 22525 8904 22559
rect 8852 22516 8904 22525
rect 11152 22516 11204 22568
rect 13820 22584 13872 22636
rect 16580 22720 16632 22772
rect 17500 22763 17552 22772
rect 17500 22729 17509 22763
rect 17509 22729 17543 22763
rect 17543 22729 17552 22763
rect 17500 22720 17552 22729
rect 20352 22720 20404 22772
rect 23296 22720 23348 22772
rect 18604 22695 18656 22704
rect 18604 22661 18613 22695
rect 18613 22661 18647 22695
rect 18647 22661 18656 22695
rect 18604 22652 18656 22661
rect 19708 22695 19760 22704
rect 19708 22661 19717 22695
rect 19717 22661 19751 22695
rect 19751 22661 19760 22695
rect 19708 22652 19760 22661
rect 23664 22720 23716 22772
rect 24308 22763 24360 22772
rect 24308 22729 24317 22763
rect 24317 22729 24351 22763
rect 24351 22729 24360 22763
rect 24308 22720 24360 22729
rect 25320 22720 25372 22772
rect 18328 22584 18380 22636
rect 19340 22584 19392 22636
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 23664 22584 23716 22636
rect 24492 22584 24544 22636
rect 13084 22516 13136 22568
rect 13912 22559 13964 22568
rect 13912 22525 13921 22559
rect 13921 22525 13955 22559
rect 13955 22525 13964 22559
rect 13912 22516 13964 22525
rect 15936 22516 15988 22568
rect 19064 22516 19116 22568
rect 21180 22516 21232 22568
rect 21640 22516 21692 22568
rect 9404 22448 9456 22500
rect 14004 22448 14056 22500
rect 4252 22380 4304 22432
rect 6920 22380 6972 22432
rect 10784 22380 10836 22432
rect 11520 22380 11572 22432
rect 15568 22380 15620 22432
rect 18788 22380 18840 22432
rect 18972 22380 19024 22432
rect 19248 22423 19300 22432
rect 19248 22389 19257 22423
rect 19257 22389 19291 22423
rect 19291 22389 19300 22423
rect 19248 22380 19300 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 16120 22176 16172 22228
rect 16396 22176 16448 22228
rect 7472 22108 7524 22160
rect 11520 22108 11572 22160
rect 12164 22040 12216 22092
rect 11152 22015 11204 22024
rect 11152 21981 11161 22015
rect 11161 21981 11195 22015
rect 11195 21981 11204 22015
rect 11152 21972 11204 21981
rect 11888 21972 11940 22024
rect 13636 21972 13688 22024
rect 4436 21879 4488 21888
rect 4436 21845 4445 21879
rect 4445 21845 4479 21879
rect 4479 21845 4488 21879
rect 4436 21836 4488 21845
rect 4712 21836 4764 21888
rect 8576 21836 8628 21888
rect 8760 21836 8812 21888
rect 10232 21836 10284 21888
rect 11428 21879 11480 21888
rect 11428 21845 11437 21879
rect 11437 21845 11471 21879
rect 11471 21845 11480 21879
rect 11428 21836 11480 21845
rect 13544 21904 13596 21956
rect 14280 22083 14332 22092
rect 14280 22049 14289 22083
rect 14289 22049 14323 22083
rect 14323 22049 14332 22083
rect 14280 22040 14332 22049
rect 16120 22040 16172 22092
rect 13360 21836 13412 21888
rect 14556 21947 14608 21956
rect 14556 21913 14565 21947
rect 14565 21913 14599 21947
rect 14599 21913 14608 21947
rect 14556 21904 14608 21913
rect 16396 21904 16448 21956
rect 18604 22176 18656 22228
rect 17040 21972 17092 22024
rect 18512 22083 18564 22092
rect 18512 22049 18521 22083
rect 18521 22049 18555 22083
rect 18555 22049 18564 22083
rect 18512 22040 18564 22049
rect 20260 22176 20312 22228
rect 21180 22219 21232 22228
rect 21180 22185 21189 22219
rect 21189 22185 21223 22219
rect 21223 22185 21232 22219
rect 21180 22176 21232 22185
rect 22008 22083 22060 22092
rect 22008 22049 22017 22083
rect 22017 22049 22051 22083
rect 22051 22049 22060 22083
rect 22008 22040 22060 22049
rect 22284 22083 22336 22092
rect 22284 22049 22293 22083
rect 22293 22049 22327 22083
rect 22327 22049 22336 22083
rect 22284 22040 22336 22049
rect 22376 22040 22428 22092
rect 23296 22040 23348 22092
rect 24216 22040 24268 22092
rect 19340 21972 19392 22024
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 24124 21972 24176 22024
rect 22376 21904 22428 21956
rect 15384 21836 15436 21888
rect 15936 21836 15988 21888
rect 19984 21836 20036 21888
rect 21548 21836 21600 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 7104 21675 7156 21684
rect 7104 21641 7113 21675
rect 7113 21641 7147 21675
rect 7147 21641 7156 21675
rect 7104 21632 7156 21641
rect 9772 21632 9824 21684
rect 11980 21632 12032 21684
rect 13820 21632 13872 21684
rect 13912 21675 13964 21684
rect 13912 21641 13921 21675
rect 13921 21641 13955 21675
rect 13955 21641 13964 21675
rect 13912 21632 13964 21641
rect 14004 21675 14056 21684
rect 14004 21641 14013 21675
rect 14013 21641 14047 21675
rect 14047 21641 14056 21675
rect 14004 21632 14056 21641
rect 14740 21632 14792 21684
rect 7656 21564 7708 21616
rect 1860 21496 1912 21548
rect 4436 21496 4488 21548
rect 4712 21496 4764 21548
rect 8944 21496 8996 21548
rect 1308 21428 1360 21480
rect 3608 21471 3660 21480
rect 3608 21437 3617 21471
rect 3617 21437 3651 21471
rect 3651 21437 3660 21471
rect 3608 21428 3660 21437
rect 4068 21428 4120 21480
rect 7656 21471 7708 21480
rect 7656 21437 7665 21471
rect 7665 21437 7699 21471
rect 7699 21437 7708 21471
rect 7656 21428 7708 21437
rect 8760 21471 8812 21480
rect 8760 21437 8769 21471
rect 8769 21437 8803 21471
rect 8803 21437 8812 21471
rect 8760 21428 8812 21437
rect 9036 21428 9088 21480
rect 12256 21564 12308 21616
rect 13636 21496 13688 21548
rect 16120 21496 16172 21548
rect 16212 21539 16264 21548
rect 16212 21505 16221 21539
rect 16221 21505 16255 21539
rect 16255 21505 16264 21539
rect 16212 21496 16264 21505
rect 17224 21564 17276 21616
rect 17684 21564 17736 21616
rect 22560 21675 22612 21684
rect 22560 21641 22569 21675
rect 22569 21641 22603 21675
rect 22603 21641 22612 21675
rect 22560 21632 22612 21641
rect 22008 21564 22060 21616
rect 20168 21496 20220 21548
rect 20444 21496 20496 21548
rect 23296 21496 23348 21548
rect 23664 21607 23716 21616
rect 23664 21573 23673 21607
rect 23673 21573 23707 21607
rect 23707 21573 23716 21607
rect 23664 21564 23716 21573
rect 24216 21564 24268 21616
rect 3792 21403 3844 21412
rect 3792 21369 3801 21403
rect 3801 21369 3835 21403
rect 3835 21369 3844 21403
rect 3792 21360 3844 21369
rect 3976 21360 4028 21412
rect 7472 21360 7524 21412
rect 7840 21360 7892 21412
rect 12256 21471 12308 21480
rect 12256 21437 12265 21471
rect 12265 21437 12299 21471
rect 12299 21437 12308 21471
rect 12256 21428 12308 21437
rect 14556 21428 14608 21480
rect 14648 21428 14700 21480
rect 15384 21471 15436 21480
rect 15384 21437 15393 21471
rect 15393 21437 15427 21471
rect 15427 21437 15436 21471
rect 15384 21428 15436 21437
rect 17592 21428 17644 21480
rect 22284 21428 22336 21480
rect 11060 21360 11112 21412
rect 5816 21292 5868 21344
rect 5908 21292 5960 21344
rect 15936 21360 15988 21412
rect 17224 21360 17276 21412
rect 13820 21292 13872 21344
rect 16856 21335 16908 21344
rect 16856 21301 16865 21335
rect 16865 21301 16899 21335
rect 16899 21301 16908 21335
rect 16856 21292 16908 21301
rect 17040 21292 17092 21344
rect 20260 21360 20312 21412
rect 18420 21292 18472 21344
rect 20444 21335 20496 21344
rect 20444 21301 20453 21335
rect 20453 21301 20487 21335
rect 20487 21301 20496 21335
rect 20444 21292 20496 21301
rect 21272 21292 21324 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 2872 21088 2924 21140
rect 7288 21088 7340 21140
rect 10508 21088 10560 21140
rect 14188 21088 14240 21140
rect 16856 21088 16908 21140
rect 7748 20952 7800 21004
rect 10416 20952 10468 21004
rect 12256 21020 12308 21072
rect 12348 21020 12400 21072
rect 16212 21020 16264 21072
rect 1860 20816 1912 20868
rect 3700 20884 3752 20936
rect 4068 20884 4120 20936
rect 4252 20927 4304 20936
rect 4252 20893 4261 20927
rect 4261 20893 4295 20927
rect 4295 20893 4304 20927
rect 4252 20884 4304 20893
rect 1768 20748 1820 20800
rect 2872 20816 2924 20868
rect 7748 20816 7800 20868
rect 11888 20884 11940 20936
rect 17040 21020 17092 21072
rect 19340 21020 19392 21072
rect 22376 21088 22428 21140
rect 24216 21088 24268 21140
rect 23480 21020 23532 21072
rect 12348 20884 12400 20936
rect 12624 20884 12676 20936
rect 14188 20884 14240 20936
rect 17316 20952 17368 21004
rect 9956 20816 10008 20868
rect 10324 20816 10376 20868
rect 8576 20748 8628 20800
rect 9588 20748 9640 20800
rect 10508 20816 10560 20868
rect 10692 20748 10744 20800
rect 15752 20927 15804 20936
rect 15752 20893 15761 20927
rect 15761 20893 15795 20927
rect 15795 20893 15804 20927
rect 15752 20884 15804 20893
rect 16120 20927 16172 20936
rect 16120 20893 16129 20927
rect 16129 20893 16163 20927
rect 16163 20893 16172 20927
rect 16120 20884 16172 20893
rect 15200 20816 15252 20868
rect 16948 20816 17000 20868
rect 17592 20927 17644 20936
rect 17592 20893 17601 20927
rect 17601 20893 17635 20927
rect 17635 20893 17644 20927
rect 17592 20884 17644 20893
rect 19156 20816 19208 20868
rect 19432 20952 19484 21004
rect 24860 20952 24912 21004
rect 22376 20884 22428 20936
rect 22652 20927 22704 20936
rect 22652 20893 22661 20927
rect 22661 20893 22695 20927
rect 22695 20893 22704 20927
rect 22652 20884 22704 20893
rect 20168 20859 20220 20868
rect 20168 20825 20177 20859
rect 20177 20825 20211 20859
rect 20211 20825 20220 20859
rect 20168 20816 20220 20825
rect 14280 20748 14332 20800
rect 15660 20748 15712 20800
rect 16856 20791 16908 20800
rect 16856 20757 16865 20791
rect 16865 20757 16899 20791
rect 16899 20757 16908 20791
rect 16856 20748 16908 20757
rect 25044 20816 25096 20868
rect 21640 20791 21692 20800
rect 21640 20757 21649 20791
rect 21649 20757 21683 20791
rect 21683 20757 21692 20791
rect 21640 20748 21692 20757
rect 22376 20791 22428 20800
rect 22376 20757 22385 20791
rect 22385 20757 22419 20791
rect 22419 20757 22428 20791
rect 22376 20748 22428 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 5724 20544 5776 20596
rect 4344 20476 4396 20528
rect 6460 20476 6512 20528
rect 8852 20544 8904 20596
rect 8944 20544 8996 20596
rect 17316 20587 17368 20596
rect 17316 20553 17325 20587
rect 17325 20553 17359 20587
rect 17359 20553 17368 20587
rect 17316 20544 17368 20553
rect 5724 20408 5776 20460
rect 7288 20476 7340 20528
rect 9036 20476 9088 20528
rect 8668 20408 8720 20460
rect 8760 20315 8812 20324
rect 8760 20281 8769 20315
rect 8769 20281 8803 20315
rect 8803 20281 8812 20315
rect 8760 20272 8812 20281
rect 9312 20340 9364 20392
rect 11520 20476 11572 20528
rect 11704 20408 11756 20460
rect 10600 20340 10652 20392
rect 16856 20476 16908 20528
rect 19340 20587 19392 20596
rect 19340 20553 19349 20587
rect 19349 20553 19383 20587
rect 19383 20553 19392 20587
rect 19340 20544 19392 20553
rect 19524 20544 19576 20596
rect 17960 20476 18012 20528
rect 18604 20476 18656 20528
rect 19616 20476 19668 20528
rect 23388 20476 23440 20528
rect 13452 20408 13504 20460
rect 18512 20451 18564 20460
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 25136 20476 25188 20528
rect 25228 20408 25280 20460
rect 11612 20272 11664 20324
rect 5816 20204 5868 20256
rect 6460 20204 6512 20256
rect 7288 20204 7340 20256
rect 8300 20247 8352 20256
rect 8300 20213 8309 20247
rect 8309 20213 8343 20247
rect 8343 20213 8352 20247
rect 8300 20204 8352 20213
rect 9036 20204 9088 20256
rect 12072 20247 12124 20256
rect 12072 20213 12081 20247
rect 12081 20213 12115 20247
rect 12115 20213 12124 20247
rect 12072 20204 12124 20213
rect 12716 20383 12768 20392
rect 12716 20349 12725 20383
rect 12725 20349 12759 20383
rect 12759 20349 12768 20383
rect 12716 20340 12768 20349
rect 21640 20340 21692 20392
rect 24676 20383 24728 20392
rect 24676 20349 24685 20383
rect 24685 20349 24719 20383
rect 24719 20349 24728 20383
rect 24676 20340 24728 20349
rect 17868 20315 17920 20324
rect 17868 20281 17877 20315
rect 17877 20281 17911 20315
rect 17911 20281 17920 20315
rect 17868 20272 17920 20281
rect 13360 20204 13412 20256
rect 14004 20204 14056 20256
rect 14096 20204 14148 20256
rect 14648 20247 14700 20256
rect 14648 20213 14657 20247
rect 14657 20213 14691 20247
rect 14691 20213 14700 20247
rect 14648 20204 14700 20213
rect 17316 20204 17368 20256
rect 18788 20204 18840 20256
rect 19800 20204 19852 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 5080 20043 5132 20052
rect 5080 20009 5089 20043
rect 5089 20009 5123 20043
rect 5123 20009 5132 20043
rect 5080 20000 5132 20009
rect 11704 20043 11756 20052
rect 11704 20009 11713 20043
rect 11713 20009 11747 20043
rect 11747 20009 11756 20043
rect 11704 20000 11756 20009
rect 13636 20000 13688 20052
rect 20536 20000 20588 20052
rect 5724 19907 5776 19916
rect 5724 19873 5733 19907
rect 5733 19873 5767 19907
rect 5767 19873 5776 19907
rect 5724 19864 5776 19873
rect 8300 19864 8352 19916
rect 8852 19864 8904 19916
rect 12164 19932 12216 19984
rect 14648 19932 14700 19984
rect 17960 19932 18012 19984
rect 7288 19796 7340 19848
rect 8944 19796 8996 19848
rect 11612 19796 11664 19848
rect 14464 19864 14516 19916
rect 17408 19864 17460 19916
rect 12440 19796 12492 19848
rect 6460 19728 6512 19780
rect 7380 19660 7432 19712
rect 7656 19728 7708 19780
rect 8668 19703 8720 19712
rect 8668 19669 8677 19703
rect 8677 19669 8711 19703
rect 8711 19669 8720 19703
rect 8668 19660 8720 19669
rect 8944 19660 8996 19712
rect 14188 19728 14240 19780
rect 14648 19771 14700 19780
rect 14648 19737 14657 19771
rect 14657 19737 14691 19771
rect 14691 19737 14700 19771
rect 14648 19728 14700 19737
rect 17776 19839 17828 19848
rect 17776 19805 17785 19839
rect 17785 19805 17819 19839
rect 17819 19805 17828 19839
rect 17776 19796 17828 19805
rect 18880 19796 18932 19848
rect 24952 19864 25004 19916
rect 25596 19796 25648 19848
rect 17592 19728 17644 19780
rect 18420 19728 18472 19780
rect 23848 19728 23900 19780
rect 9588 19660 9640 19712
rect 14740 19703 14792 19712
rect 14740 19669 14749 19703
rect 14749 19669 14783 19703
rect 14783 19669 14792 19703
rect 14740 19660 14792 19669
rect 19064 19660 19116 19712
rect 19340 19703 19392 19712
rect 19340 19669 19349 19703
rect 19349 19669 19383 19703
rect 19383 19669 19392 19703
rect 19340 19660 19392 19669
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 1492 19456 1544 19508
rect 3608 19456 3660 19508
rect 4436 19456 4488 19508
rect 9404 19456 9456 19508
rect 4528 19388 4580 19440
rect 7288 19388 7340 19440
rect 9312 19388 9364 19440
rect 13452 19456 13504 19508
rect 14004 19388 14056 19440
rect 16304 19388 16356 19440
rect 18696 19456 18748 19508
rect 3884 19363 3936 19372
rect 3884 19329 3893 19363
rect 3893 19329 3927 19363
rect 3927 19329 3936 19363
rect 3884 19320 3936 19329
rect 6276 19320 6328 19372
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 8392 19320 8444 19372
rect 8668 19320 8720 19372
rect 12164 19363 12216 19372
rect 12164 19329 12173 19363
rect 12173 19329 12207 19363
rect 12207 19329 12216 19363
rect 12164 19320 12216 19329
rect 14648 19320 14700 19372
rect 14832 19320 14884 19372
rect 17592 19320 17644 19372
rect 19248 19388 19300 19440
rect 19524 19456 19576 19508
rect 20536 19456 20588 19508
rect 21364 19456 21416 19508
rect 21916 19456 21968 19508
rect 22560 19388 22612 19440
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 9036 19252 9088 19304
rect 9588 19252 9640 19304
rect 12348 19252 12400 19304
rect 14004 19295 14056 19304
rect 14004 19261 14013 19295
rect 14013 19261 14047 19295
rect 14047 19261 14056 19295
rect 14004 19252 14056 19261
rect 14464 19252 14516 19304
rect 16580 19252 16632 19304
rect 17776 19252 17828 19304
rect 19156 19252 19208 19304
rect 10324 19184 10376 19236
rect 10968 19184 11020 19236
rect 19248 19184 19300 19236
rect 20812 19320 20864 19372
rect 21088 19363 21140 19372
rect 21088 19329 21097 19363
rect 21097 19329 21131 19363
rect 21131 19329 21140 19363
rect 21088 19320 21140 19329
rect 20628 19252 20680 19304
rect 21916 19252 21968 19304
rect 22008 19295 22060 19304
rect 22008 19261 22017 19295
rect 22017 19261 22051 19295
rect 22051 19261 22060 19295
rect 22008 19252 22060 19261
rect 22284 19295 22336 19304
rect 22284 19261 22293 19295
rect 22293 19261 22327 19295
rect 22327 19261 22336 19295
rect 22284 19252 22336 19261
rect 22836 19252 22888 19304
rect 20996 19184 21048 19236
rect 7840 19116 7892 19168
rect 8760 19159 8812 19168
rect 8760 19125 8769 19159
rect 8769 19125 8803 19159
rect 8803 19125 8812 19159
rect 8760 19116 8812 19125
rect 10784 19116 10836 19168
rect 11152 19116 11204 19168
rect 12440 19116 12492 19168
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 14832 19159 14884 19168
rect 14832 19125 14841 19159
rect 14841 19125 14875 19159
rect 14875 19125 14884 19159
rect 14832 19116 14884 19125
rect 24032 19159 24084 19168
rect 24032 19125 24041 19159
rect 24041 19125 24075 19159
rect 24075 19125 24084 19159
rect 24032 19116 24084 19125
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 8944 18955 8996 18964
rect 8944 18921 8953 18955
rect 8953 18921 8987 18955
rect 8987 18921 8996 18955
rect 8944 18912 8996 18921
rect 3792 18844 3844 18896
rect 10600 18912 10652 18964
rect 10784 18912 10836 18964
rect 12164 18912 12216 18964
rect 14188 18912 14240 18964
rect 18328 18912 18380 18964
rect 18972 18955 19024 18964
rect 18972 18921 18981 18955
rect 18981 18921 19015 18955
rect 19015 18921 19024 18955
rect 18972 18912 19024 18921
rect 22284 18912 22336 18964
rect 13360 18844 13412 18896
rect 13912 18844 13964 18896
rect 1308 18776 1360 18828
rect 4896 18776 4948 18828
rect 5908 18776 5960 18828
rect 12716 18776 12768 18828
rect 14188 18776 14240 18828
rect 14832 18819 14884 18828
rect 14832 18785 14841 18819
rect 14841 18785 14875 18819
rect 14875 18785 14884 18819
rect 14832 18776 14884 18785
rect 19064 18844 19116 18896
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 5172 18708 5224 18760
rect 11152 18708 11204 18760
rect 12808 18708 12860 18760
rect 13820 18708 13872 18760
rect 17776 18776 17828 18828
rect 16212 18751 16264 18760
rect 16212 18717 16221 18751
rect 16221 18717 16255 18751
rect 16255 18717 16264 18751
rect 16212 18708 16264 18717
rect 18972 18708 19024 18760
rect 20444 18708 20496 18760
rect 22008 18708 22060 18760
rect 8484 18615 8536 18624
rect 8484 18581 8493 18615
rect 8493 18581 8527 18615
rect 8527 18581 8536 18615
rect 8484 18572 8536 18581
rect 8668 18615 8720 18624
rect 8668 18581 8677 18615
rect 8677 18581 8711 18615
rect 8711 18581 8720 18615
rect 8668 18572 8720 18581
rect 9312 18572 9364 18624
rect 9588 18572 9640 18624
rect 10876 18572 10928 18624
rect 11612 18572 11664 18624
rect 11980 18572 12032 18624
rect 13636 18640 13688 18692
rect 13360 18615 13412 18624
rect 13360 18581 13369 18615
rect 13369 18581 13403 18615
rect 13403 18581 13412 18615
rect 13360 18572 13412 18581
rect 19432 18640 19484 18692
rect 20904 18640 20956 18692
rect 22560 18683 22612 18692
rect 22560 18649 22569 18683
rect 22569 18649 22603 18683
rect 22603 18649 22612 18683
rect 22560 18640 22612 18649
rect 18420 18572 18472 18624
rect 19524 18572 19576 18624
rect 20720 18572 20772 18624
rect 22376 18572 22428 18624
rect 22928 18572 22980 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 7564 18368 7616 18420
rect 9680 18411 9732 18420
rect 9680 18377 9689 18411
rect 9689 18377 9723 18411
rect 9723 18377 9732 18411
rect 9680 18368 9732 18377
rect 11060 18368 11112 18420
rect 12440 18300 12492 18352
rect 5264 18232 5316 18284
rect 3792 18207 3844 18216
rect 3792 18173 3801 18207
rect 3801 18173 3835 18207
rect 3835 18173 3844 18207
rect 3792 18164 3844 18173
rect 4988 18028 5040 18080
rect 7748 18232 7800 18284
rect 7104 18164 7156 18216
rect 7840 18207 7892 18216
rect 7840 18173 7849 18207
rect 7849 18173 7883 18207
rect 7883 18173 7892 18207
rect 7840 18164 7892 18173
rect 8484 18096 8536 18148
rect 11980 18232 12032 18284
rect 12900 18368 12952 18420
rect 13360 18368 13412 18420
rect 18328 18368 18380 18420
rect 12716 18232 12768 18284
rect 19156 18343 19208 18352
rect 19156 18309 19165 18343
rect 19165 18309 19199 18343
rect 19199 18309 19208 18343
rect 19156 18300 19208 18309
rect 19432 18300 19484 18352
rect 10692 18164 10744 18216
rect 10968 18207 11020 18216
rect 10968 18173 10977 18207
rect 10977 18173 11011 18207
rect 11011 18173 11020 18207
rect 10968 18164 11020 18173
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 12256 18207 12308 18216
rect 12256 18173 12265 18207
rect 12265 18173 12299 18207
rect 12299 18173 12308 18207
rect 12256 18164 12308 18173
rect 12440 18164 12492 18216
rect 14464 18164 14516 18216
rect 15016 18232 15068 18284
rect 17500 18275 17552 18284
rect 17500 18241 17509 18275
rect 17509 18241 17543 18275
rect 17543 18241 17552 18275
rect 17500 18232 17552 18241
rect 15384 18164 15436 18216
rect 16028 18164 16080 18216
rect 16212 18164 16264 18216
rect 16488 18164 16540 18216
rect 24032 18232 24084 18284
rect 12348 18096 12400 18148
rect 12532 18096 12584 18148
rect 13636 18096 13688 18148
rect 18512 18096 18564 18148
rect 22928 18164 22980 18216
rect 23664 18164 23716 18216
rect 21456 18139 21508 18148
rect 21456 18105 21465 18139
rect 21465 18105 21499 18139
rect 21499 18105 21508 18139
rect 21456 18096 21508 18105
rect 7748 18028 7800 18080
rect 10692 18028 10744 18080
rect 11612 18028 11664 18080
rect 12256 18028 12308 18080
rect 13544 18071 13596 18080
rect 13544 18037 13553 18071
rect 13553 18037 13587 18071
rect 13587 18037 13596 18071
rect 13544 18028 13596 18037
rect 14004 18028 14056 18080
rect 14740 18028 14792 18080
rect 16580 18028 16632 18080
rect 17500 18028 17552 18080
rect 20168 18028 20220 18080
rect 24032 18028 24084 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 6276 17867 6328 17876
rect 6276 17833 6285 17867
rect 6285 17833 6319 17867
rect 6319 17833 6328 17867
rect 6276 17824 6328 17833
rect 7380 17824 7432 17876
rect 11888 17824 11940 17876
rect 12532 17867 12584 17876
rect 12532 17833 12541 17867
rect 12541 17833 12575 17867
rect 12575 17833 12584 17867
rect 12532 17824 12584 17833
rect 12716 17824 12768 17876
rect 12900 17824 12952 17876
rect 15108 17824 15160 17876
rect 19248 17824 19300 17876
rect 20628 17824 20680 17876
rect 6920 17688 6972 17740
rect 8392 17688 8444 17740
rect 9404 17688 9456 17740
rect 11980 17688 12032 17740
rect 14464 17688 14516 17740
rect 14832 17731 14884 17740
rect 14832 17697 14841 17731
rect 14841 17697 14875 17731
rect 14875 17697 14884 17731
rect 14832 17688 14884 17697
rect 16396 17688 16448 17740
rect 17040 17688 17092 17740
rect 20904 17688 20956 17740
rect 22560 17824 22612 17876
rect 4712 17620 4764 17672
rect 8760 17620 8812 17672
rect 9588 17620 9640 17672
rect 12532 17620 12584 17672
rect 14648 17663 14700 17672
rect 14648 17629 14657 17663
rect 14657 17629 14691 17663
rect 14691 17629 14700 17663
rect 14648 17620 14700 17629
rect 15108 17620 15160 17672
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 15660 17620 15712 17672
rect 16212 17620 16264 17672
rect 25044 17620 25096 17672
rect 7288 17484 7340 17536
rect 9680 17552 9732 17604
rect 10508 17595 10560 17604
rect 10508 17561 10517 17595
rect 10517 17561 10551 17595
rect 10551 17561 10560 17595
rect 10508 17552 10560 17561
rect 11336 17595 11388 17604
rect 11336 17561 11345 17595
rect 11345 17561 11379 17595
rect 11379 17561 11388 17595
rect 11336 17552 11388 17561
rect 8576 17484 8628 17536
rect 8760 17527 8812 17536
rect 8760 17493 8769 17527
rect 8769 17493 8803 17527
rect 8803 17493 8812 17527
rect 8760 17484 8812 17493
rect 9496 17527 9548 17536
rect 9496 17493 9505 17527
rect 9505 17493 9539 17527
rect 9539 17493 9548 17527
rect 9496 17484 9548 17493
rect 10140 17484 10192 17536
rect 12716 17484 12768 17536
rect 13544 17484 13596 17536
rect 14740 17527 14792 17536
rect 14740 17493 14749 17527
rect 14749 17493 14783 17527
rect 14783 17493 14792 17527
rect 14740 17484 14792 17493
rect 15384 17484 15436 17536
rect 18880 17552 18932 17604
rect 20168 17595 20220 17604
rect 20168 17561 20177 17595
rect 20177 17561 20211 17595
rect 20211 17561 20220 17595
rect 20168 17552 20220 17561
rect 20720 17552 20772 17604
rect 23664 17552 23716 17604
rect 16396 17484 16448 17536
rect 24216 17484 24268 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 8852 17280 8904 17332
rect 3700 17212 3752 17264
rect 3976 17255 4028 17264
rect 3976 17221 3985 17255
rect 3985 17221 4019 17255
rect 4019 17221 4028 17255
rect 3976 17212 4028 17221
rect 8116 17212 8168 17264
rect 8944 17212 8996 17264
rect 9496 17280 9548 17332
rect 10508 17280 10560 17332
rect 16580 17280 16632 17332
rect 4620 17144 4672 17196
rect 8760 17144 8812 17196
rect 6552 17119 6604 17128
rect 6552 17085 6561 17119
rect 6561 17085 6595 17119
rect 6595 17085 6604 17119
rect 6552 17076 6604 17085
rect 6920 17076 6972 17128
rect 8852 17076 8904 17128
rect 12072 17212 12124 17264
rect 12808 17212 12860 17264
rect 13360 17212 13412 17264
rect 15108 17255 15160 17264
rect 15108 17221 15117 17255
rect 15117 17221 15151 17255
rect 15151 17221 15160 17255
rect 15108 17212 15160 17221
rect 17132 17144 17184 17196
rect 20904 17280 20956 17332
rect 17960 17212 18012 17264
rect 20720 17212 20772 17264
rect 24860 17212 24912 17264
rect 9956 17008 10008 17060
rect 10508 17119 10560 17128
rect 10508 17085 10517 17119
rect 10517 17085 10551 17119
rect 10551 17085 10560 17119
rect 10508 17076 10560 17085
rect 10968 17076 11020 17128
rect 11336 17076 11388 17128
rect 12900 17119 12952 17128
rect 12900 17085 12909 17119
rect 12909 17085 12943 17119
rect 12943 17085 12952 17119
rect 12900 17076 12952 17085
rect 13360 17076 13412 17128
rect 18604 17076 18656 17128
rect 19156 17076 19208 17128
rect 20444 17119 20496 17128
rect 20444 17085 20453 17119
rect 20453 17085 20487 17119
rect 20487 17085 20496 17119
rect 20444 17076 20496 17085
rect 11060 17008 11112 17060
rect 12440 17008 12492 17060
rect 14188 17008 14240 17060
rect 15016 17008 15068 17060
rect 16396 17008 16448 17060
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 11612 16940 11664 16992
rect 14464 16940 14516 16992
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 17224 16940 17276 16992
rect 22100 17187 22152 17196
rect 22100 17153 22109 17187
rect 22109 17153 22143 17187
rect 22143 17153 22152 17187
rect 22100 17144 22152 17153
rect 23940 17187 23992 17196
rect 23940 17153 23949 17187
rect 23949 17153 23983 17187
rect 23983 17153 23992 17187
rect 23940 17144 23992 17153
rect 23296 17076 23348 17128
rect 21732 17008 21784 17060
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 6920 16736 6972 16788
rect 7196 16736 7248 16788
rect 8116 16736 8168 16788
rect 8392 16668 8444 16720
rect 8576 16736 8628 16788
rect 10140 16736 10192 16788
rect 8760 16668 8812 16720
rect 9956 16668 10008 16720
rect 6644 16600 6696 16652
rect 8484 16600 8536 16652
rect 1492 16532 1544 16584
rect 8300 16532 8352 16584
rect 9036 16532 9088 16584
rect 12808 16736 12860 16788
rect 10968 16600 11020 16652
rect 14280 16668 14332 16720
rect 12808 16600 12860 16652
rect 14924 16643 14976 16652
rect 14924 16609 14933 16643
rect 14933 16609 14967 16643
rect 14967 16609 14976 16643
rect 19708 16736 19760 16788
rect 20168 16736 20220 16788
rect 18696 16668 18748 16720
rect 14924 16600 14976 16609
rect 16028 16600 16080 16652
rect 9588 16532 9640 16584
rect 1308 16464 1360 16516
rect 7196 16464 7248 16516
rect 10324 16532 10376 16584
rect 10876 16575 10928 16584
rect 10876 16541 10885 16575
rect 10885 16541 10919 16575
rect 10919 16541 10928 16575
rect 10876 16532 10928 16541
rect 12716 16532 12768 16584
rect 20444 16575 20496 16584
rect 20444 16541 20453 16575
rect 20453 16541 20487 16575
rect 20487 16541 20496 16575
rect 20444 16532 20496 16541
rect 20904 16600 20956 16652
rect 22008 16643 22060 16652
rect 22008 16609 22017 16643
rect 22017 16609 22051 16643
rect 22051 16609 22060 16643
rect 22008 16600 22060 16609
rect 22652 16600 22704 16652
rect 23664 16600 23716 16652
rect 5172 16396 5224 16448
rect 10232 16464 10284 16516
rect 22652 16464 22704 16516
rect 8484 16439 8536 16448
rect 8484 16405 8493 16439
rect 8493 16405 8527 16439
rect 8527 16405 8536 16439
rect 8484 16396 8536 16405
rect 9956 16396 10008 16448
rect 11704 16396 11756 16448
rect 11796 16439 11848 16448
rect 11796 16405 11805 16439
rect 11805 16405 11839 16439
rect 11839 16405 11848 16439
rect 11796 16396 11848 16405
rect 15292 16439 15344 16448
rect 15292 16405 15301 16439
rect 15301 16405 15335 16439
rect 15335 16405 15344 16439
rect 15292 16396 15344 16405
rect 16304 16396 16356 16448
rect 17132 16396 17184 16448
rect 17224 16396 17276 16448
rect 17960 16396 18012 16448
rect 18696 16396 18748 16448
rect 20168 16396 20220 16448
rect 21180 16396 21232 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 7288 16192 7340 16244
rect 10508 16192 10560 16244
rect 11428 16192 11480 16244
rect 11520 16192 11572 16244
rect 13544 16192 13596 16244
rect 13728 16235 13780 16244
rect 13728 16201 13737 16235
rect 13737 16201 13771 16235
rect 13771 16201 13780 16235
rect 13728 16192 13780 16201
rect 14740 16235 14792 16244
rect 14740 16201 14749 16235
rect 14749 16201 14783 16235
rect 14783 16201 14792 16235
rect 14740 16192 14792 16201
rect 17316 16192 17368 16244
rect 2504 16167 2556 16176
rect 2504 16133 2513 16167
rect 2513 16133 2547 16167
rect 2547 16133 2556 16167
rect 2504 16124 2556 16133
rect 7196 16124 7248 16176
rect 11796 16124 11848 16176
rect 13360 16124 13412 16176
rect 15936 16167 15988 16176
rect 15936 16133 15945 16167
rect 15945 16133 15979 16167
rect 15979 16133 15988 16167
rect 15936 16124 15988 16133
rect 17040 16124 17092 16176
rect 17224 16124 17276 16176
rect 18604 16235 18656 16244
rect 18604 16201 18613 16235
rect 18613 16201 18647 16235
rect 18647 16201 18656 16235
rect 18604 16192 18656 16201
rect 18696 16192 18748 16244
rect 21088 16192 21140 16244
rect 6644 16099 6696 16108
rect 6644 16065 6653 16099
rect 6653 16065 6687 16099
rect 6687 16065 6696 16099
rect 6644 16056 6696 16065
rect 3792 15988 3844 16040
rect 4068 15988 4120 16040
rect 8300 15988 8352 16040
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 10324 16056 10376 16108
rect 12716 16056 12768 16108
rect 16580 16056 16632 16108
rect 20812 16124 20864 16176
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 23480 16099 23532 16108
rect 23480 16065 23489 16099
rect 23489 16065 23523 16099
rect 23523 16065 23532 16099
rect 23480 16056 23532 16065
rect 24400 16124 24452 16176
rect 10232 15988 10284 16040
rect 11428 15988 11480 16040
rect 12256 16031 12308 16040
rect 12256 15997 12265 16031
rect 12265 15997 12299 16031
rect 12299 15997 12308 16031
rect 12256 15988 12308 15997
rect 19708 16031 19760 16040
rect 19708 15997 19717 16031
rect 19717 15997 19751 16031
rect 19751 15997 19760 16031
rect 19708 15988 19760 15997
rect 12072 15920 12124 15972
rect 22284 15988 22336 16040
rect 22560 16031 22612 16040
rect 22560 15997 22569 16031
rect 22569 15997 22603 16031
rect 22603 15997 22612 16031
rect 22560 15988 22612 15997
rect 23388 15988 23440 16040
rect 23664 15920 23716 15972
rect 1768 15852 1820 15904
rect 14280 15895 14332 15904
rect 14280 15861 14289 15895
rect 14289 15861 14323 15895
rect 14323 15861 14332 15895
rect 14280 15852 14332 15861
rect 15568 15852 15620 15904
rect 22192 15852 22244 15904
rect 22468 15852 22520 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 8760 15691 8812 15700
rect 8760 15657 8769 15691
rect 8769 15657 8803 15691
rect 8803 15657 8812 15691
rect 8760 15648 8812 15657
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 10140 15648 10192 15700
rect 11704 15648 11756 15700
rect 19892 15580 19944 15632
rect 11336 15512 11388 15564
rect 11428 15512 11480 15564
rect 14188 15512 14240 15564
rect 17408 15512 17460 15564
rect 20996 15580 21048 15632
rect 8484 15351 8536 15360
rect 8484 15317 8493 15351
rect 8493 15317 8527 15351
rect 8527 15317 8536 15351
rect 8484 15308 8536 15317
rect 10324 15308 10376 15360
rect 10876 15308 10928 15360
rect 11980 15308 12032 15360
rect 12256 15308 12308 15360
rect 13360 15444 13412 15496
rect 13728 15444 13780 15496
rect 15292 15444 15344 15496
rect 17684 15444 17736 15496
rect 21180 15512 21232 15564
rect 21272 15444 21324 15496
rect 24216 15444 24268 15496
rect 12624 15376 12676 15428
rect 15476 15376 15528 15428
rect 12808 15351 12860 15360
rect 12808 15317 12817 15351
rect 12817 15317 12851 15351
rect 12851 15317 12860 15351
rect 12808 15308 12860 15317
rect 15660 15308 15712 15360
rect 16764 15308 16816 15360
rect 18696 15351 18748 15360
rect 18696 15317 18705 15351
rect 18705 15317 18739 15351
rect 18739 15317 18748 15351
rect 18696 15308 18748 15317
rect 21548 15376 21600 15428
rect 24952 15376 25004 15428
rect 19708 15308 19760 15360
rect 20628 15351 20680 15360
rect 20628 15317 20637 15351
rect 20637 15317 20671 15351
rect 20671 15317 20680 15351
rect 20628 15308 20680 15317
rect 21916 15351 21968 15360
rect 21916 15317 21925 15351
rect 21925 15317 21959 15351
rect 21959 15317 21968 15351
rect 21916 15308 21968 15317
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 8760 15104 8812 15156
rect 9588 15104 9640 15156
rect 9404 15079 9456 15088
rect 9404 15045 9413 15079
rect 9413 15045 9447 15079
rect 9447 15045 9456 15079
rect 9404 15036 9456 15045
rect 12164 15104 12216 15156
rect 17316 15104 17368 15156
rect 18696 15104 18748 15156
rect 18880 15147 18932 15156
rect 18880 15113 18889 15147
rect 18889 15113 18923 15147
rect 18923 15113 18932 15147
rect 18880 15104 18932 15113
rect 22376 15104 22428 15156
rect 12256 15036 12308 15088
rect 15384 15036 15436 15088
rect 16120 15079 16172 15088
rect 16120 15045 16129 15079
rect 16129 15045 16163 15079
rect 16163 15045 16172 15079
rect 16120 15036 16172 15045
rect 16304 15036 16356 15088
rect 19708 15036 19760 15088
rect 12440 14968 12492 15020
rect 10876 14900 10928 14952
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 15476 14968 15528 15020
rect 16764 14968 16816 15020
rect 16948 14968 17000 15020
rect 18604 14968 18656 15020
rect 14832 14943 14884 14952
rect 14832 14909 14841 14943
rect 14841 14909 14875 14943
rect 14875 14909 14884 14943
rect 14832 14900 14884 14909
rect 13636 14832 13688 14884
rect 17868 14900 17920 14952
rect 18788 14900 18840 14952
rect 19800 15011 19852 15020
rect 19800 14977 19809 15011
rect 19809 14977 19843 15011
rect 19843 14977 19852 15011
rect 19800 14968 19852 14977
rect 23572 14968 23624 15020
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 24768 14943 24820 14952
rect 24768 14909 24777 14943
rect 24777 14909 24811 14943
rect 24811 14909 24820 14943
rect 24768 14900 24820 14909
rect 17592 14832 17644 14884
rect 9956 14764 10008 14816
rect 16672 14764 16724 14816
rect 18880 14764 18932 14816
rect 19800 14764 19852 14816
rect 21272 14764 21324 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 10416 14560 10468 14612
rect 10692 14560 10744 14612
rect 11336 14492 11388 14544
rect 9956 14467 10008 14476
rect 9956 14433 9965 14467
rect 9965 14433 9999 14467
rect 9999 14433 10008 14467
rect 9956 14424 10008 14433
rect 11980 14356 12032 14408
rect 12256 14492 12308 14544
rect 12716 14560 12768 14612
rect 14556 14492 14608 14544
rect 14464 14424 14516 14476
rect 15384 14560 15436 14612
rect 15844 14560 15896 14612
rect 17040 14560 17092 14612
rect 21640 14560 21692 14612
rect 15384 14467 15436 14476
rect 15384 14433 15393 14467
rect 15393 14433 15427 14467
rect 15427 14433 15436 14467
rect 15384 14424 15436 14433
rect 16396 14424 16448 14476
rect 17132 14424 17184 14476
rect 20812 14424 20864 14476
rect 21180 14467 21232 14476
rect 21180 14433 21189 14467
rect 21189 14433 21223 14467
rect 21223 14433 21232 14467
rect 21180 14424 21232 14433
rect 18512 14356 18564 14408
rect 20904 14399 20956 14408
rect 20904 14365 20913 14399
rect 20913 14365 20947 14399
rect 20947 14365 20956 14399
rect 20904 14356 20956 14365
rect 22284 14356 22336 14408
rect 22652 14356 22704 14408
rect 10232 14331 10284 14340
rect 10232 14297 10241 14331
rect 10241 14297 10275 14331
rect 10275 14297 10284 14331
rect 10232 14288 10284 14297
rect 12532 14331 12584 14340
rect 12532 14297 12541 14331
rect 12541 14297 12575 14331
rect 12575 14297 12584 14331
rect 12532 14288 12584 14297
rect 13636 14288 13688 14340
rect 15936 14288 15988 14340
rect 9864 14220 9916 14272
rect 10968 14220 11020 14272
rect 15752 14220 15804 14272
rect 17224 14220 17276 14272
rect 19432 14263 19484 14272
rect 19432 14229 19441 14263
rect 19441 14229 19475 14263
rect 19475 14229 19484 14263
rect 19432 14220 19484 14229
rect 19708 14220 19760 14272
rect 21824 14220 21876 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 9956 14016 10008 14068
rect 10140 14016 10192 14068
rect 10324 14016 10376 14068
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 9588 13948 9640 14000
rect 10324 13880 10376 13932
rect 10600 13880 10652 13932
rect 12440 14016 12492 14068
rect 17224 14016 17276 14068
rect 13544 13991 13596 14000
rect 13544 13957 13553 13991
rect 13553 13957 13587 13991
rect 13587 13957 13596 13991
rect 13544 13948 13596 13957
rect 17408 13991 17460 14000
rect 17408 13957 17417 13991
rect 17417 13957 17451 13991
rect 17451 13957 17460 13991
rect 17408 13948 17460 13957
rect 18420 14016 18472 14068
rect 19248 14016 19300 14068
rect 22376 14016 22428 14068
rect 22652 14016 22704 14068
rect 17868 13948 17920 14000
rect 19708 13991 19760 14000
rect 19708 13957 19717 13991
rect 19717 13957 19751 13991
rect 19751 13957 19760 13991
rect 19708 13948 19760 13957
rect 19984 13948 20036 14000
rect 16580 13880 16632 13932
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 20260 13880 20312 13932
rect 20720 13880 20772 13932
rect 22744 13880 22796 13932
rect 23848 13880 23900 13932
rect 1308 13812 1360 13864
rect 9496 13812 9548 13864
rect 11796 13744 11848 13796
rect 13636 13812 13688 13864
rect 17408 13812 17460 13864
rect 19340 13812 19392 13864
rect 20352 13812 20404 13864
rect 22100 13812 22152 13864
rect 24676 13855 24728 13864
rect 24676 13821 24685 13855
rect 24685 13821 24719 13855
rect 24719 13821 24728 13855
rect 24676 13812 24728 13821
rect 13544 13744 13596 13796
rect 14280 13744 14332 13796
rect 9864 13676 9916 13728
rect 15108 13676 15160 13728
rect 17868 13676 17920 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 5816 13472 5868 13524
rect 8484 13336 8536 13388
rect 6828 13311 6880 13320
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 8392 13268 8444 13320
rect 9588 13404 9640 13456
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 11612 13515 11664 13524
rect 11612 13481 11621 13515
rect 11621 13481 11655 13515
rect 11655 13481 11664 13515
rect 11612 13472 11664 13481
rect 11980 13515 12032 13524
rect 11980 13481 11989 13515
rect 11989 13481 12023 13515
rect 12023 13481 12032 13515
rect 11980 13472 12032 13481
rect 12072 13472 12124 13524
rect 12440 13472 12492 13524
rect 12808 13336 12860 13388
rect 15384 13336 15436 13388
rect 15936 13472 15988 13524
rect 19248 13472 19300 13524
rect 19340 13404 19392 13456
rect 14464 13268 14516 13320
rect 18512 13336 18564 13388
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 19432 13268 19484 13320
rect 20996 13268 21048 13320
rect 7104 13243 7156 13252
rect 7104 13209 7113 13243
rect 7113 13209 7147 13243
rect 7147 13209 7156 13243
rect 7104 13200 7156 13209
rect 11520 13200 11572 13252
rect 11980 13200 12032 13252
rect 14004 13200 14056 13252
rect 14556 13200 14608 13252
rect 14832 13243 14884 13252
rect 14832 13209 14841 13243
rect 14841 13209 14875 13243
rect 14875 13209 14884 13243
rect 14832 13200 14884 13209
rect 15292 13200 15344 13252
rect 16120 13200 16172 13252
rect 8760 13132 8812 13184
rect 17224 13132 17276 13184
rect 19892 13243 19944 13252
rect 19892 13209 19901 13243
rect 19901 13209 19935 13243
rect 19935 13209 19944 13243
rect 19892 13200 19944 13209
rect 21364 13200 21416 13252
rect 21180 13132 21232 13184
rect 22284 13472 22336 13524
rect 21732 13268 21784 13320
rect 25504 13200 25556 13252
rect 22008 13175 22060 13184
rect 22008 13141 22017 13175
rect 22017 13141 22051 13175
rect 22051 13141 22060 13175
rect 22008 13132 22060 13141
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 7748 12928 7800 12980
rect 11796 12928 11848 12980
rect 6644 12860 6696 12912
rect 8392 12860 8444 12912
rect 6552 12792 6604 12844
rect 9680 12860 9732 12912
rect 9956 12860 10008 12912
rect 11520 12903 11572 12912
rect 11520 12869 11529 12903
rect 11529 12869 11563 12903
rect 11563 12869 11572 12903
rect 11520 12860 11572 12869
rect 12808 12860 12860 12912
rect 15292 12928 15344 12980
rect 15752 12928 15804 12980
rect 13912 12860 13964 12912
rect 14372 12860 14424 12912
rect 15200 12860 15252 12912
rect 16120 12971 16172 12980
rect 16120 12937 16129 12971
rect 16129 12937 16163 12971
rect 16163 12937 16172 12971
rect 16120 12928 16172 12937
rect 17224 12971 17276 12980
rect 17224 12937 17233 12971
rect 17233 12937 17267 12971
rect 17267 12937 17276 12971
rect 17224 12928 17276 12937
rect 17316 12971 17368 12980
rect 17316 12937 17325 12971
rect 17325 12937 17359 12971
rect 17359 12937 17368 12971
rect 17316 12928 17368 12937
rect 18328 12928 18380 12980
rect 15936 12792 15988 12844
rect 8760 12767 8812 12776
rect 8760 12733 8769 12767
rect 8769 12733 8803 12767
rect 8803 12733 8812 12767
rect 8760 12724 8812 12733
rect 14832 12724 14884 12776
rect 18328 12724 18380 12776
rect 20904 12928 20956 12980
rect 20996 12928 21048 12980
rect 21456 12860 21508 12912
rect 13360 12656 13412 12708
rect 13728 12656 13780 12708
rect 14280 12656 14332 12708
rect 14648 12699 14700 12708
rect 14648 12665 14657 12699
rect 14657 12665 14691 12699
rect 14691 12665 14700 12699
rect 14648 12656 14700 12665
rect 15936 12656 15988 12708
rect 16120 12656 16172 12708
rect 21180 12724 21232 12776
rect 22468 12792 22520 12844
rect 23296 12835 23348 12844
rect 23296 12801 23305 12835
rect 23305 12801 23339 12835
rect 23339 12801 23348 12835
rect 23296 12792 23348 12801
rect 24768 12767 24820 12776
rect 24768 12733 24777 12767
rect 24777 12733 24811 12767
rect 24811 12733 24820 12767
rect 24768 12724 24820 12733
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 15476 12588 15528 12597
rect 18604 12631 18656 12640
rect 18604 12597 18613 12631
rect 18613 12597 18647 12631
rect 18647 12597 18656 12631
rect 18604 12588 18656 12597
rect 21824 12656 21876 12708
rect 20536 12588 20588 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 10876 12384 10928 12436
rect 9680 12248 9732 12300
rect 10968 12248 11020 12300
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 13912 12384 13964 12436
rect 14464 12427 14516 12436
rect 14464 12393 14473 12427
rect 14473 12393 14507 12427
rect 14507 12393 14516 12427
rect 14464 12384 14516 12393
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 15660 12384 15712 12393
rect 16028 12384 16080 12436
rect 15936 12316 15988 12368
rect 15292 12248 15344 12300
rect 17500 12384 17552 12436
rect 24860 12316 24912 12368
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 19984 12248 20036 12300
rect 21548 12291 21600 12300
rect 21548 12257 21557 12291
rect 21557 12257 21591 12291
rect 21591 12257 21600 12291
rect 21548 12248 21600 12257
rect 21824 12248 21876 12300
rect 22192 12248 22244 12300
rect 16948 12180 17000 12232
rect 18880 12180 18932 12232
rect 22008 12180 22060 12232
rect 12808 12112 12860 12164
rect 16488 12112 16540 12164
rect 13268 12087 13320 12096
rect 13268 12053 13277 12087
rect 13277 12053 13311 12087
rect 13311 12053 13320 12087
rect 13268 12044 13320 12053
rect 13728 12087 13780 12096
rect 13728 12053 13737 12087
rect 13737 12053 13771 12087
rect 13771 12053 13780 12087
rect 13728 12044 13780 12053
rect 17408 12044 17460 12096
rect 17868 12112 17920 12164
rect 20168 12112 20220 12164
rect 19800 12044 19852 12096
rect 20996 12044 21048 12096
rect 21088 12087 21140 12096
rect 21088 12053 21097 12087
rect 21097 12053 21131 12087
rect 21131 12053 21140 12087
rect 21088 12044 21140 12053
rect 25044 12044 25096 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 13268 11840 13320 11892
rect 13176 11772 13228 11824
rect 15108 11840 15160 11892
rect 15752 11840 15804 11892
rect 17868 11840 17920 11892
rect 10968 11704 11020 11756
rect 15108 11704 15160 11756
rect 16764 11772 16816 11824
rect 18328 11840 18380 11892
rect 19984 11883 20036 11892
rect 19984 11849 19993 11883
rect 19993 11849 20027 11883
rect 20027 11849 20036 11883
rect 19984 11840 20036 11849
rect 18512 11815 18564 11824
rect 18512 11781 18521 11815
rect 18521 11781 18555 11815
rect 18555 11781 18564 11815
rect 18512 11772 18564 11781
rect 19800 11772 19852 11824
rect 21180 11840 21232 11892
rect 20812 11772 20864 11824
rect 22836 11704 22888 11756
rect 16488 11636 16540 11688
rect 19892 11636 19944 11688
rect 24032 11679 24084 11688
rect 24032 11645 24041 11679
rect 24041 11645 24075 11679
rect 24075 11645 24084 11679
rect 24032 11636 24084 11645
rect 14556 11611 14608 11620
rect 14556 11577 14565 11611
rect 14565 11577 14599 11611
rect 14599 11577 14608 11611
rect 14556 11568 14608 11577
rect 22008 11568 22060 11620
rect 17040 11543 17092 11552
rect 17040 11509 17049 11543
rect 17049 11509 17083 11543
rect 17083 11509 17092 11543
rect 17040 11500 17092 11509
rect 18328 11500 18380 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 14004 11296 14056 11348
rect 15108 11160 15160 11212
rect 15292 11160 15344 11212
rect 20628 11092 20680 11144
rect 15200 11024 15252 11076
rect 16304 11024 16356 11076
rect 20812 11067 20864 11076
rect 20812 11033 20821 11067
rect 20821 11033 20855 11067
rect 20855 11033 20864 11067
rect 20812 11024 20864 11033
rect 23940 11024 23992 11076
rect 19616 10999 19668 11008
rect 19616 10965 19625 10999
rect 19625 10965 19659 10999
rect 19659 10965 19668 10999
rect 19616 10956 19668 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 15292 10795 15344 10804
rect 15292 10761 15301 10795
rect 15301 10761 15335 10795
rect 15335 10761 15344 10795
rect 15292 10752 15344 10761
rect 19616 10752 19668 10804
rect 10232 10684 10284 10736
rect 14832 10659 14884 10668
rect 14832 10625 14841 10659
rect 14841 10625 14875 10659
rect 14875 10625 14884 10659
rect 14832 10616 14884 10625
rect 18328 10616 18380 10668
rect 19340 10616 19392 10668
rect 20536 10659 20588 10668
rect 20536 10625 20545 10659
rect 20545 10625 20579 10659
rect 20579 10625 20588 10659
rect 20536 10616 20588 10625
rect 23664 10616 23716 10668
rect 19984 10548 20036 10600
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 12440 10480 12492 10532
rect 20812 10480 20864 10532
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 18236 10455 18288 10464
rect 18236 10421 18245 10455
rect 18245 10421 18279 10455
rect 18279 10421 18288 10455
rect 18236 10412 18288 10421
rect 20628 10412 20680 10464
rect 23296 10412 23348 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 20996 10140 21048 10192
rect 18236 10072 18288 10124
rect 13452 10004 13504 10056
rect 18696 10004 18748 10056
rect 21364 10004 21416 10056
rect 19432 9936 19484 9988
rect 24952 10004 25004 10056
rect 16856 9911 16908 9920
rect 16856 9877 16865 9911
rect 16865 9877 16899 9911
rect 16899 9877 16908 9911
rect 16856 9868 16908 9877
rect 21732 9868 21784 9920
rect 24032 9868 24084 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 16212 9596 16264 9648
rect 21916 9596 21968 9648
rect 19064 9528 19116 9580
rect 21088 9528 21140 9580
rect 4436 9460 4488 9512
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 23388 9460 23440 9512
rect 6552 9435 6604 9444
rect 6552 9401 6561 9435
rect 6561 9401 6595 9435
rect 6595 9401 6604 9435
rect 6552 9392 6604 9401
rect 17592 9392 17644 9444
rect 17684 9324 17736 9376
rect 22744 9367 22796 9376
rect 22744 9333 22753 9367
rect 22753 9333 22787 9367
rect 22787 9333 22796 9367
rect 22744 9324 22796 9333
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 3608 9052 3660 9104
rect 4896 9052 4948 9104
rect 22468 9052 22520 9104
rect 20628 8916 20680 8968
rect 22652 8916 22704 8968
rect 24860 8959 24912 8968
rect 24860 8925 24869 8959
rect 24869 8925 24903 8959
rect 24903 8925 24912 8959
rect 24860 8916 24912 8925
rect 22560 8780 22612 8832
rect 23480 8780 23532 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 19156 8551 19208 8560
rect 19156 8517 19165 8551
rect 19165 8517 19199 8551
rect 19199 8517 19208 8551
rect 19156 8508 19208 8517
rect 21272 8508 21324 8560
rect 22652 8440 22704 8492
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 23296 8415 23348 8424
rect 23296 8381 23305 8415
rect 23305 8381 23339 8415
rect 23339 8381 23348 8415
rect 23296 8372 23348 8381
rect 24676 8415 24728 8424
rect 24676 8381 24685 8415
rect 24685 8381 24719 8415
rect 24719 8381 24728 8415
rect 24676 8372 24728 8381
rect 20720 8304 20772 8356
rect 21272 8304 21324 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 6552 8032 6604 8084
rect 6828 8032 6880 8084
rect 22836 8032 22888 8084
rect 6552 7828 6604 7880
rect 19892 7828 19944 7880
rect 20536 7828 20588 7880
rect 23480 7828 23532 7880
rect 24860 7828 24912 7880
rect 4344 7803 4396 7812
rect 4344 7769 4353 7803
rect 4353 7769 4387 7803
rect 4387 7769 4396 7803
rect 4344 7760 4396 7769
rect 9220 7760 9272 7812
rect 24492 7760 24544 7812
rect 20812 7692 20864 7744
rect 21088 7735 21140 7744
rect 21088 7701 21097 7735
rect 21097 7701 21131 7735
rect 21131 7701 21140 7735
rect 21088 7692 21140 7701
rect 22468 7692 22520 7744
rect 22836 7692 22888 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 16948 7420 17000 7472
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 20720 7352 20772 7404
rect 23388 7352 23440 7404
rect 20904 7284 20956 7336
rect 21364 7284 21416 7336
rect 22284 7284 22336 7336
rect 20628 7216 20680 7268
rect 22560 7148 22612 7200
rect 23388 7148 23440 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 15844 6740 15896 6792
rect 20812 6783 20864 6792
rect 20812 6749 20821 6783
rect 20821 6749 20855 6783
rect 20855 6749 20864 6783
rect 20812 6740 20864 6749
rect 22836 6783 22888 6792
rect 22836 6749 22845 6783
rect 22845 6749 22879 6783
rect 22879 6749 22888 6783
rect 22836 6740 22888 6749
rect 24952 6740 25004 6792
rect 21824 6715 21876 6724
rect 21824 6681 21833 6715
rect 21833 6681 21867 6715
rect 21867 6681 21876 6715
rect 21824 6672 21876 6681
rect 25044 6672 25096 6724
rect 18328 6604 18380 6656
rect 24676 6647 24728 6656
rect 24676 6613 24685 6647
rect 24685 6613 24719 6647
rect 24719 6613 24728 6647
rect 24676 6604 24728 6613
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 1860 6443 1912 6452
rect 1860 6409 1869 6443
rect 1869 6409 1903 6443
rect 1903 6409 1912 6443
rect 1860 6400 1912 6409
rect 4344 6400 4396 6452
rect 11612 6400 11664 6452
rect 2412 6264 2464 6316
rect 3332 6264 3384 6316
rect 21088 6264 21140 6316
rect 22008 6307 22060 6316
rect 22008 6273 22017 6307
rect 22017 6273 22051 6307
rect 22051 6273 22060 6307
rect 22008 6264 22060 6273
rect 22560 6264 22612 6316
rect 2780 6196 2832 6248
rect 20720 6196 20772 6248
rect 21456 6196 21508 6248
rect 21916 6196 21968 6248
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 2504 6060 2556 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 3332 5856 3384 5908
rect 4160 5856 4212 5908
rect 9312 5856 9364 5908
rect 20904 5856 20956 5908
rect 4988 5788 5040 5840
rect 5908 5720 5960 5772
rect 10784 5720 10836 5772
rect 20444 5720 20496 5772
rect 21548 5720 21600 5772
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 3056 5652 3108 5704
rect 8668 5652 8720 5704
rect 17684 5695 17736 5704
rect 17684 5661 17693 5695
rect 17693 5661 17727 5695
rect 17727 5661 17736 5695
rect 17684 5652 17736 5661
rect 20352 5652 20404 5704
rect 20628 5652 20680 5704
rect 1860 5627 1912 5636
rect 1860 5593 1869 5627
rect 1869 5593 1903 5627
rect 1903 5593 1912 5627
rect 1860 5584 1912 5593
rect 2136 5584 2188 5636
rect 9312 5584 9364 5636
rect 3608 5559 3660 5568
rect 3608 5525 3617 5559
rect 3617 5525 3651 5559
rect 3651 5525 3660 5559
rect 3608 5516 3660 5525
rect 3884 5516 3936 5568
rect 4804 5516 4856 5568
rect 6368 5516 6420 5568
rect 8852 5516 8904 5568
rect 10324 5516 10376 5568
rect 21180 5584 21232 5636
rect 14096 5516 14148 5568
rect 21732 5516 21784 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 3792 5355 3844 5364
rect 3792 5321 3801 5355
rect 3801 5321 3835 5355
rect 3835 5321 3844 5355
rect 3792 5312 3844 5321
rect 4436 5312 4488 5364
rect 5172 5355 5224 5364
rect 5172 5321 5181 5355
rect 5181 5321 5215 5355
rect 5215 5321 5224 5355
rect 5172 5312 5224 5321
rect 1676 5176 1728 5228
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 19340 5244 19392 5296
rect 2320 5108 2372 5160
rect 6000 5176 6052 5228
rect 17776 5219 17828 5228
rect 17776 5185 17785 5219
rect 17785 5185 17819 5219
rect 17819 5185 17828 5219
rect 17776 5176 17828 5185
rect 19524 5219 19576 5228
rect 19524 5185 19533 5219
rect 19533 5185 19567 5219
rect 19567 5185 19576 5219
rect 19524 5176 19576 5185
rect 22192 5219 22244 5228
rect 22192 5185 22201 5219
rect 22201 5185 22235 5219
rect 22235 5185 22244 5219
rect 22192 5176 22244 5185
rect 24032 5219 24084 5228
rect 24032 5185 24041 5219
rect 24041 5185 24075 5219
rect 24075 5185 24084 5219
rect 24032 5176 24084 5185
rect 20260 5108 20312 5160
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 22468 5108 22520 5117
rect 24584 5151 24636 5160
rect 24584 5117 24593 5151
rect 24593 5117 24627 5151
rect 24627 5117 24636 5151
rect 24584 5108 24636 5117
rect 1676 4972 1728 5024
rect 5356 4972 5408 5024
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 4160 4811 4212 4820
rect 4160 4777 4169 4811
rect 4169 4777 4203 4811
rect 4203 4777 4212 4811
rect 4160 4768 4212 4777
rect 5908 4811 5960 4820
rect 5908 4777 5917 4811
rect 5917 4777 5951 4811
rect 5951 4777 5960 4811
rect 5908 4768 5960 4777
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 7012 4768 7064 4820
rect 8484 4811 8536 4820
rect 8484 4777 8493 4811
rect 8493 4777 8527 4811
rect 8527 4777 8536 4811
rect 8484 4768 8536 4777
rect 12348 4768 12400 4820
rect 17776 4768 17828 4820
rect 10048 4700 10100 4752
rect 15200 4700 15252 4752
rect 22652 4700 22704 4752
rect 19892 4675 19944 4684
rect 19892 4641 19901 4675
rect 19901 4641 19935 4675
rect 19935 4641 19944 4675
rect 19892 4632 19944 4641
rect 21732 4675 21784 4684
rect 21732 4641 21741 4675
rect 21741 4641 21775 4675
rect 21775 4641 21784 4675
rect 21732 4632 21784 4641
rect 3424 4564 3476 4616
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 7196 4564 7248 4616
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 9864 4564 9916 4616
rect 11612 4564 11664 4616
rect 18328 4564 18380 4616
rect 18604 4564 18656 4616
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 22744 4564 22796 4616
rect 7656 4539 7708 4548
rect 7656 4505 7665 4539
rect 7665 4505 7699 4539
rect 7699 4505 7708 4539
rect 7656 4496 7708 4505
rect 7840 4496 7892 4548
rect 9036 4496 9088 4548
rect 20168 4496 20220 4548
rect 23388 4496 23440 4548
rect 1768 4428 1820 4480
rect 6552 4428 6604 4480
rect 8484 4428 8536 4480
rect 10232 4428 10284 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 3884 3952 3936 4004
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 6000 4131 6052 4140
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 7196 4131 7248 4140
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 8576 4088 8628 4140
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 11244 4088 11296 4140
rect 13636 4131 13688 4140
rect 13636 4097 13645 4131
rect 13645 4097 13679 4131
rect 13679 4097 13688 4131
rect 13636 4088 13688 4097
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 16672 4088 16724 4140
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 20260 4088 20312 4140
rect 22100 4088 22152 4140
rect 22376 4088 22428 4140
rect 24676 4088 24728 4140
rect 13452 4020 13504 4072
rect 16396 4020 16448 4072
rect 17500 4020 17552 4072
rect 20076 4020 20128 4072
rect 24768 4063 24820 4072
rect 24768 4029 24777 4063
rect 24777 4029 24811 4063
rect 24811 4029 24820 4063
rect 24768 4020 24820 4029
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 5448 3952 5500 4004
rect 6920 3952 6972 4004
rect 8852 3995 8904 4004
rect 8852 3961 8861 3995
rect 8861 3961 8895 3995
rect 8895 3961 8904 3995
rect 8852 3952 8904 3961
rect 10324 3952 10376 4004
rect 20720 3952 20772 4004
rect 24952 3952 25004 4004
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 5540 3884 5592 3936
rect 6828 3884 6880 3936
rect 10048 3884 10100 3936
rect 10876 3927 10928 3936
rect 10876 3893 10885 3927
rect 10885 3893 10919 3927
rect 10919 3893 10928 3927
rect 10876 3884 10928 3893
rect 11244 3927 11296 3936
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 11704 3884 11756 3936
rect 22560 3884 22612 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 1860 3680 1912 3732
rect 2872 3680 2924 3732
rect 4988 3680 5040 3732
rect 5724 3680 5776 3732
rect 8576 3723 8628 3732
rect 8576 3689 8585 3723
rect 8585 3689 8619 3723
rect 8619 3689 8628 3723
rect 8576 3680 8628 3689
rect 9312 3723 9364 3732
rect 9312 3689 9321 3723
rect 9321 3689 9355 3723
rect 9355 3689 9364 3723
rect 9312 3680 9364 3689
rect 12532 3680 12584 3732
rect 12716 3680 12768 3732
rect 18696 3680 18748 3732
rect 16120 3612 16172 3664
rect 18972 3612 19024 3664
rect 10876 3544 10928 3596
rect 1492 3476 1544 3528
rect 2044 3476 2096 3528
rect 2780 3519 2832 3528
rect 2780 3485 2789 3519
rect 2789 3485 2823 3519
rect 2823 3485 2832 3519
rect 2780 3476 2832 3485
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4988 3476 5040 3528
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 7840 3476 7892 3528
rect 9772 3476 9824 3528
rect 10048 3476 10100 3528
rect 12532 3519 12584 3528
rect 12532 3485 12541 3519
rect 12541 3485 12575 3519
rect 12575 3485 12584 3519
rect 12532 3476 12584 3485
rect 12716 3544 12768 3596
rect 14924 3544 14976 3596
rect 16028 3544 16080 3596
rect 17868 3544 17920 3596
rect 14832 3476 14884 3528
rect 15568 3476 15620 3528
rect 15476 3408 15528 3460
rect 17408 3476 17460 3528
rect 21640 3476 21692 3528
rect 23112 3476 23164 3528
rect 19708 3408 19760 3460
rect 21732 3408 21784 3460
rect 4620 3340 4672 3392
rect 18604 3340 18656 3392
rect 19892 3340 19944 3392
rect 21824 3340 21876 3392
rect 22836 3340 22888 3392
rect 24584 3340 24636 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 2872 3136 2924 3188
rect 4160 3136 4212 3188
rect 8300 3136 8352 3188
rect 13360 3136 13412 3188
rect 21456 3136 21508 3188
rect 22652 3136 22704 3188
rect 23112 3179 23164 3188
rect 23112 3145 23121 3179
rect 23121 3145 23155 3179
rect 23155 3145 23164 3179
rect 23112 3136 23164 3145
rect 24860 3136 24912 3188
rect 2136 3043 2188 3052
rect 2136 3009 2145 3043
rect 2145 3009 2179 3043
rect 2179 3009 2188 3043
rect 2136 3000 2188 3009
rect 2412 3000 2464 3052
rect 4620 3043 4672 3052
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4620 3000 4672 3009
rect 5540 3000 5592 3052
rect 6092 3000 6144 3052
rect 7196 3000 7248 3052
rect 8484 3000 8536 3052
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9588 3000 9640 3052
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 10508 3000 10560 3052
rect 13728 3068 13780 3120
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 13544 3000 13596 3052
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 2780 2932 2832 2984
rect 3332 2932 3384 2984
rect 10140 2932 10192 2984
rect 13360 2975 13412 2984
rect 13360 2941 13369 2975
rect 13369 2941 13403 2975
rect 13403 2941 13412 2975
rect 13360 2932 13412 2941
rect 14188 2932 14240 2984
rect 15660 2932 15712 2984
rect 4804 2907 4856 2916
rect 4804 2873 4813 2907
rect 4813 2873 4847 2907
rect 4847 2873 4856 2907
rect 4804 2864 4856 2873
rect 17132 2864 17184 2916
rect 20168 2932 20220 2984
rect 23388 2932 23440 2984
rect 4712 2796 4764 2848
rect 7472 2839 7524 2848
rect 7472 2805 7481 2839
rect 7481 2805 7515 2839
rect 7515 2805 7524 2839
rect 7472 2796 7524 2805
rect 16764 2796 16816 2848
rect 17960 2796 18012 2848
rect 20812 2796 20864 2848
rect 22468 2796 22520 2848
rect 25320 3043 25372 3052
rect 25320 3009 25329 3043
rect 25329 3009 25363 3043
rect 25363 3009 25372 3043
rect 25320 3000 25372 3009
rect 24124 2796 24176 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 2320 2635 2372 2644
rect 2320 2601 2329 2635
rect 2329 2601 2363 2635
rect 2363 2601 2372 2635
rect 2320 2592 2372 2601
rect 3976 2592 4028 2644
rect 3516 2456 3568 2508
rect 3792 2456 3844 2508
rect 7472 2592 7524 2644
rect 9864 2635 9916 2644
rect 9864 2601 9873 2635
rect 9873 2601 9907 2635
rect 9907 2601 9916 2635
rect 9864 2592 9916 2601
rect 15936 2592 15988 2644
rect 18788 2592 18840 2644
rect 25320 2592 25372 2644
rect 7104 2524 7156 2576
rect 7656 2524 7708 2576
rect 12348 2524 12400 2576
rect 17684 2524 17736 2576
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 7380 2388 7432 2440
rect 3608 2320 3660 2372
rect 4068 2320 4120 2372
rect 7288 2320 7340 2372
rect 7564 2388 7616 2440
rect 8208 2320 8260 2372
rect 10232 2388 10284 2440
rect 11980 2456 12032 2508
rect 14556 2456 14608 2508
rect 15292 2456 15344 2508
rect 17960 2456 18012 2508
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 14648 2431 14700 2440
rect 14648 2397 14657 2431
rect 14657 2397 14691 2431
rect 14691 2397 14700 2431
rect 14648 2388 14700 2397
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 19524 2431 19576 2440
rect 19524 2397 19533 2431
rect 19533 2397 19567 2431
rect 19567 2397 19576 2431
rect 19524 2388 19576 2397
rect 5724 2252 5776 2304
rect 7104 2252 7156 2304
rect 10416 2252 10468 2304
rect 12624 2320 12676 2372
rect 13820 2320 13872 2372
rect 18328 2320 18380 2372
rect 24860 2456 24912 2508
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 15016 2252 15068 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 7288 2048 7340 2100
rect 11796 2048 11848 2100
<< metal2 >>
rect 1490 56200 1546 57000
rect 1858 56200 1914 57000
rect 2226 56200 2282 57000
rect 2594 56200 2650 57000
rect 2962 56200 3018 57000
rect 3330 56200 3386 57000
rect 3698 56200 3754 57000
rect 4066 56200 4122 57000
rect 4434 56200 4490 57000
rect 4802 56200 4858 57000
rect 5170 56200 5226 57000
rect 5276 56222 5488 56250
rect 1306 53000 1362 53009
rect 1306 52935 1362 52944
rect 1320 52630 1348 52935
rect 1308 52624 1360 52630
rect 1308 52566 1360 52572
rect 1306 50552 1362 50561
rect 1306 50487 1362 50496
rect 1320 50386 1348 50487
rect 1308 50380 1360 50386
rect 1308 50322 1360 50328
rect 1504 49298 1532 56200
rect 1768 52896 1820 52902
rect 1768 52838 1820 52844
rect 1676 52012 1728 52018
rect 1676 51954 1728 51960
rect 1688 51066 1716 51954
rect 1676 51060 1728 51066
rect 1676 51002 1728 51008
rect 1780 50930 1808 52838
rect 1872 52698 1900 56200
rect 2240 53718 2268 56200
rect 2320 54188 2372 54194
rect 2320 54130 2372 54136
rect 2228 53712 2280 53718
rect 2228 53654 2280 53660
rect 2228 53576 2280 53582
rect 2226 53544 2228 53553
rect 2280 53544 2282 53553
rect 2226 53479 2282 53488
rect 1860 52692 1912 52698
rect 1860 52634 1912 52640
rect 2332 50998 2360 54130
rect 2608 52986 2636 56200
rect 2976 55214 3004 56200
rect 2884 55186 3004 55214
rect 2608 52958 2820 52986
rect 2320 50992 2372 50998
rect 2320 50934 2372 50940
rect 1768 50924 1820 50930
rect 1768 50866 1820 50872
rect 2792 50862 2820 52958
rect 2884 51474 2912 55186
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 3344 51950 3372 56200
rect 3424 53712 3476 53718
rect 3424 53654 3476 53660
rect 3332 51944 3384 51950
rect 3332 51886 3384 51892
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 2872 51468 2924 51474
rect 2872 51410 2924 51416
rect 2780 50856 2832 50862
rect 2780 50798 2832 50804
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 3436 50386 3464 53654
rect 3516 52692 3568 52698
rect 3516 52634 3568 52640
rect 3424 50380 3476 50386
rect 3424 50322 3476 50328
rect 3528 49910 3556 52634
rect 3712 52562 3740 56200
rect 3974 55448 4030 55457
rect 3974 55383 4030 55392
rect 3988 54330 4016 55383
rect 3976 54324 4028 54330
rect 3976 54266 4028 54272
rect 3792 53984 3844 53990
rect 3792 53926 3844 53932
rect 3804 52630 3832 53926
rect 3988 53582 4016 54266
rect 3976 53576 4028 53582
rect 3976 53518 4028 53524
rect 4080 52986 4108 56200
rect 4448 53174 4476 56200
rect 4816 55214 4844 56200
rect 5184 56114 5212 56200
rect 5276 56114 5304 56222
rect 5184 56086 5304 56114
rect 4816 55186 4936 55214
rect 4620 54188 4672 54194
rect 4620 54130 4672 54136
rect 4436 53168 4488 53174
rect 4436 53110 4488 53116
rect 4528 53100 4580 53106
rect 4528 53042 4580 53048
rect 4080 52958 4384 52986
rect 3792 52624 3844 52630
rect 3792 52566 3844 52572
rect 3700 52556 3752 52562
rect 3700 52498 3752 52504
rect 3976 51808 4028 51814
rect 3976 51750 4028 51756
rect 3988 51406 4016 51750
rect 3976 51400 4028 51406
rect 3976 51342 4028 51348
rect 4252 51264 4304 51270
rect 4252 51206 4304 51212
rect 4160 50788 4212 50794
rect 4160 50730 4212 50736
rect 3516 49904 3568 49910
rect 3516 49846 3568 49852
rect 1952 49836 2004 49842
rect 1952 49778 2004 49784
rect 1492 49292 1544 49298
rect 1492 49234 1544 49240
rect 1306 48104 1362 48113
rect 1306 48039 1308 48048
rect 1360 48039 1362 48048
rect 1308 48010 1360 48016
rect 1308 45960 1360 45966
rect 1308 45902 1360 45908
rect 1320 45665 1348 45902
rect 1306 45656 1362 45665
rect 1306 45591 1308 45600
rect 1360 45591 1362 45600
rect 1308 45562 1360 45568
rect 1216 43648 1268 43654
rect 1216 43590 1268 43596
rect 1228 43314 1256 43590
rect 1216 43308 1268 43314
rect 1216 43250 1268 43256
rect 1228 43217 1256 43250
rect 1214 43208 1270 43217
rect 1214 43143 1270 43152
rect 1400 41472 1452 41478
rect 1400 41414 1452 41420
rect 1412 41154 1440 41414
rect 1964 41274 1992 49778
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 4068 48000 4120 48006
rect 4068 47942 4120 47948
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 2228 43104 2280 43110
rect 2228 43046 2280 43052
rect 2240 42702 2268 43046
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2228 42696 2280 42702
rect 2228 42638 2280 42644
rect 3976 42628 4028 42634
rect 3976 42570 4028 42576
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 1952 41268 2004 41274
rect 1952 41210 2004 41216
rect 1320 41138 1440 41154
rect 1308 41132 1440 41138
rect 1360 41126 1440 41132
rect 1308 41074 1360 41080
rect 1320 40769 1348 41074
rect 1768 40928 1820 40934
rect 1768 40870 1820 40876
rect 1306 40760 1362 40769
rect 1306 40695 1362 40704
rect 1780 40526 1808 40870
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 1768 40520 1820 40526
rect 1768 40462 1820 40468
rect 1860 40384 1912 40390
rect 1860 40326 1912 40332
rect 1400 38752 1452 38758
rect 1400 38694 1452 38700
rect 1412 38434 1440 38694
rect 1320 38406 1440 38434
rect 1320 38350 1348 38406
rect 1308 38344 1360 38350
rect 1306 38312 1308 38321
rect 1360 38312 1362 38321
rect 1306 38247 1362 38256
rect 1768 38208 1820 38214
rect 1768 38150 1820 38156
rect 1780 37874 1808 38150
rect 1768 37868 1820 37874
rect 1768 37810 1820 37816
rect 1584 36576 1636 36582
rect 1584 36518 1636 36524
rect 1596 36174 1624 36518
rect 1584 36168 1636 36174
rect 1584 36110 1636 36116
rect 1596 35873 1624 36110
rect 1768 36032 1820 36038
rect 1768 35974 1820 35980
rect 1582 35864 1638 35873
rect 1582 35799 1638 35808
rect 1780 35698 1808 35974
rect 1768 35692 1820 35698
rect 1768 35634 1820 35640
rect 1216 33856 1268 33862
rect 1216 33798 1268 33804
rect 1228 33522 1256 33798
rect 1216 33516 1268 33522
rect 1216 33458 1268 33464
rect 1228 33425 1256 33458
rect 1214 33416 1270 33425
rect 1214 33351 1270 33360
rect 1768 33312 1820 33318
rect 1768 33254 1820 33260
rect 1780 32910 1808 33254
rect 1768 32904 1820 32910
rect 1768 32846 1820 32852
rect 1584 32768 1636 32774
rect 1584 32710 1636 32716
rect 1308 31272 1360 31278
rect 1308 31214 1360 31220
rect 1320 30977 1348 31214
rect 1306 30968 1362 30977
rect 1306 30903 1362 30912
rect 1308 28620 1360 28626
rect 1308 28562 1360 28568
rect 1320 28529 1348 28562
rect 1306 28520 1362 28529
rect 1306 28455 1362 28464
rect 1596 27062 1624 32710
rect 1872 30802 1900 40326
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 2688 37664 2740 37670
rect 2688 37606 2740 37612
rect 1952 31340 2004 31346
rect 1952 31282 2004 31288
rect 1860 30796 1912 30802
rect 1860 30738 1912 30744
rect 1768 28552 1820 28558
rect 1768 28494 1820 28500
rect 1584 27056 1636 27062
rect 1584 26998 1636 27004
rect 1780 26042 1808 28494
rect 1964 28218 1992 31282
rect 2700 29714 2728 37606
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 3792 30660 3844 30666
rect 3792 30602 3844 30608
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 2688 29708 2740 29714
rect 2688 29650 2740 29656
rect 3424 29572 3476 29578
rect 3424 29514 3476 29520
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 1952 28212 2004 28218
rect 1952 28154 2004 28160
rect 3332 28076 3384 28082
rect 3332 28018 3384 28024
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2044 26376 2096 26382
rect 2044 26318 2096 26324
rect 1768 26036 1820 26042
rect 1768 25978 1820 25984
rect 1860 24064 1912 24070
rect 1860 24006 1912 24012
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1308 23656 1360 23662
rect 1306 23624 1308 23633
rect 1360 23624 1362 23633
rect 1306 23559 1362 23568
rect 1780 22778 1808 23666
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 1872 21554 1900 24006
rect 2056 23322 2084 26318
rect 2780 26308 2832 26314
rect 2780 26250 2832 26256
rect 2792 26081 2820 26250
rect 2778 26072 2834 26081
rect 2778 26007 2834 26016
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 2780 25832 2832 25838
rect 2780 25774 2832 25780
rect 2792 24206 2820 25774
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2884 23322 2912 25842
rect 3344 25770 3372 28018
rect 3436 27130 3464 29514
rect 3804 28218 3832 30602
rect 3988 28506 4016 42570
rect 4080 38962 4108 47942
rect 4172 42362 4200 50730
rect 4264 49910 4292 51206
rect 4356 50862 4384 52958
rect 4540 52154 4568 53042
rect 4528 52148 4580 52154
rect 4528 52090 4580 52096
rect 4344 50856 4396 50862
rect 4344 50798 4396 50804
rect 4436 50312 4488 50318
rect 4436 50254 4488 50260
rect 4252 49904 4304 49910
rect 4252 49846 4304 49852
rect 4160 42356 4212 42362
rect 4160 42298 4212 42304
rect 4252 42220 4304 42226
rect 4252 42162 4304 42168
rect 4068 38956 4120 38962
rect 4068 38898 4120 38904
rect 4068 35488 4120 35494
rect 4068 35430 4120 35436
rect 4080 28626 4108 35430
rect 4264 29850 4292 42162
rect 4448 40769 4476 50254
rect 4632 43382 4660 54130
rect 4712 53100 4764 53106
rect 4712 53042 4764 53048
rect 4724 45014 4752 53042
rect 4908 51950 4936 55186
rect 5460 53258 5488 56222
rect 5538 56200 5594 57000
rect 5906 56200 5962 57000
rect 6274 56200 6330 57000
rect 6642 56200 6698 57000
rect 7010 56200 7066 57000
rect 7378 56200 7434 57000
rect 7746 56200 7802 57000
rect 7852 56222 8064 56250
rect 5552 53718 5580 56200
rect 5920 54126 5948 56200
rect 5908 54120 5960 54126
rect 5908 54062 5960 54068
rect 5540 53712 5592 53718
rect 5540 53654 5592 53660
rect 5460 53230 5580 53258
rect 5172 52488 5224 52494
rect 5172 52430 5224 52436
rect 4896 51944 4948 51950
rect 4896 51886 4948 51892
rect 4896 51808 4948 51814
rect 4896 51750 4948 51756
rect 4712 45008 4764 45014
rect 4712 44950 4764 44956
rect 4620 43376 4672 43382
rect 4620 43318 4672 43324
rect 4908 42770 4936 51750
rect 5080 50244 5132 50250
rect 5080 50186 5132 50192
rect 4896 42764 4948 42770
rect 4896 42706 4948 42712
rect 4804 42628 4856 42634
rect 4804 42570 4856 42576
rect 4620 41132 4672 41138
rect 4620 41074 4672 41080
rect 4434 40760 4490 40769
rect 4434 40695 4490 40704
rect 4632 32570 4660 41074
rect 4620 32564 4672 32570
rect 4620 32506 4672 32512
rect 4816 31210 4844 42570
rect 5092 42362 5120 50186
rect 5080 42356 5132 42362
rect 5080 42298 5132 42304
rect 5184 41818 5212 52430
rect 5552 51406 5580 53230
rect 6288 53174 6316 56200
rect 6552 53440 6604 53446
rect 6552 53382 6604 53388
rect 6276 53168 6328 53174
rect 6276 53110 6328 53116
rect 6564 53106 6592 53382
rect 6552 53100 6604 53106
rect 6552 53042 6604 53048
rect 6656 52494 6684 56200
rect 6828 53576 6880 53582
rect 6828 53518 6880 53524
rect 5908 52488 5960 52494
rect 5908 52430 5960 52436
rect 6644 52488 6696 52494
rect 6644 52430 6696 52436
rect 5540 51400 5592 51406
rect 5540 51342 5592 51348
rect 5448 50924 5500 50930
rect 5448 50866 5500 50872
rect 5264 44396 5316 44402
rect 5264 44338 5316 44344
rect 5172 41812 5224 41818
rect 5172 41754 5224 41760
rect 5276 38010 5304 44338
rect 5460 42362 5488 50866
rect 5816 50312 5868 50318
rect 5816 50254 5868 50260
rect 5828 44538 5856 50254
rect 5920 46170 5948 52430
rect 6736 51332 6788 51338
rect 6736 51274 6788 51280
rect 5908 46164 5960 46170
rect 5908 46106 5960 46112
rect 6644 44736 6696 44742
rect 6644 44678 6696 44684
rect 5816 44532 5868 44538
rect 5816 44474 5868 44480
rect 6656 44418 6684 44678
rect 6748 44538 6776 51274
rect 6840 50522 6868 53518
rect 7024 51474 7052 56200
rect 7392 53650 7420 56200
rect 7380 53644 7432 53650
rect 7380 53586 7432 53592
rect 7378 53544 7434 53553
rect 7378 53479 7434 53488
rect 7288 52488 7340 52494
rect 7288 52430 7340 52436
rect 7196 52012 7248 52018
rect 7196 51954 7248 51960
rect 6920 51468 6972 51474
rect 6920 51410 6972 51416
rect 7012 51468 7064 51474
rect 7012 51410 7064 51416
rect 6932 51066 6960 51410
rect 7104 51400 7156 51406
rect 7104 51342 7156 51348
rect 7012 51332 7064 51338
rect 7012 51274 7064 51280
rect 6920 51060 6972 51066
rect 6920 51002 6972 51008
rect 6828 50516 6880 50522
rect 6828 50458 6880 50464
rect 6920 45892 6972 45898
rect 6920 45834 6972 45840
rect 6736 44532 6788 44538
rect 6736 44474 6788 44480
rect 6656 44402 6776 44418
rect 6656 44396 6788 44402
rect 6656 44390 6736 44396
rect 6736 44338 6788 44344
rect 5448 42356 5500 42362
rect 5448 42298 5500 42304
rect 6092 42016 6144 42022
rect 6092 41958 6144 41964
rect 5724 41472 5776 41478
rect 5724 41414 5776 41420
rect 5264 38004 5316 38010
rect 5264 37946 5316 37952
rect 4988 37868 5040 37874
rect 4988 37810 5040 37816
rect 5000 32570 5028 37810
rect 5540 36916 5592 36922
rect 5540 36858 5592 36864
rect 5264 36712 5316 36718
rect 5264 36654 5316 36660
rect 4988 32564 5040 32570
rect 4988 32506 5040 32512
rect 5276 32366 5304 36654
rect 5552 35834 5580 36858
rect 5632 36848 5684 36854
rect 5632 36790 5684 36796
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 5552 35154 5580 35770
rect 5644 35698 5672 36790
rect 5632 35692 5684 35698
rect 5632 35634 5684 35640
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 5552 34066 5580 35090
rect 5540 34060 5592 34066
rect 5540 34002 5592 34008
rect 5356 33448 5408 33454
rect 5356 33390 5408 33396
rect 5368 32570 5396 33390
rect 5552 32978 5580 34002
rect 5540 32972 5592 32978
rect 5540 32914 5592 32920
rect 5356 32564 5408 32570
rect 5356 32506 5408 32512
rect 5552 32502 5580 32914
rect 5448 32496 5500 32502
rect 5446 32464 5448 32473
rect 5540 32496 5592 32502
rect 5500 32464 5502 32473
rect 5540 32438 5592 32444
rect 5446 32399 5502 32408
rect 5264 32360 5316 32366
rect 5264 32302 5316 32308
rect 4804 31204 4856 31210
rect 4804 31146 4856 31152
rect 5736 31142 5764 41414
rect 5816 39296 5868 39302
rect 5816 39238 5868 39244
rect 5828 37806 5856 39238
rect 5816 37800 5868 37806
rect 5816 37742 5868 37748
rect 5828 36718 5856 37742
rect 5816 36712 5868 36718
rect 5816 36654 5868 36660
rect 6000 36712 6052 36718
rect 6000 36654 6052 36660
rect 6012 35834 6040 36654
rect 6104 36530 6132 41958
rect 6184 41676 6236 41682
rect 6184 41618 6236 41624
rect 6196 41274 6224 41618
rect 6748 41414 6776 44338
rect 6656 41386 6776 41414
rect 6184 41268 6236 41274
rect 6184 41210 6236 41216
rect 6196 40526 6224 41210
rect 6552 40588 6604 40594
rect 6552 40530 6604 40536
rect 6184 40520 6236 40526
rect 6184 40462 6236 40468
rect 6196 39506 6224 40462
rect 6564 39642 6592 40530
rect 6552 39636 6604 39642
rect 6552 39578 6604 39584
rect 6184 39500 6236 39506
rect 6184 39442 6236 39448
rect 6552 38208 6604 38214
rect 6552 38150 6604 38156
rect 6564 37806 6592 38150
rect 6552 37800 6604 37806
rect 6552 37742 6604 37748
rect 6564 37262 6592 37742
rect 6656 37670 6684 41386
rect 6932 38554 6960 45834
rect 7024 43926 7052 51274
rect 7116 44470 7144 51342
rect 7208 51338 7236 51954
rect 7196 51332 7248 51338
rect 7196 51274 7248 51280
rect 7196 45960 7248 45966
rect 7196 45902 7248 45908
rect 7104 44464 7156 44470
rect 7104 44406 7156 44412
rect 7012 43920 7064 43926
rect 7012 43862 7064 43868
rect 7104 43648 7156 43654
rect 7104 43590 7156 43596
rect 7012 42220 7064 42226
rect 7012 42162 7064 42168
rect 7024 42022 7052 42162
rect 7012 42016 7064 42022
rect 7012 41958 7064 41964
rect 6920 38548 6972 38554
rect 6920 38490 6972 38496
rect 6920 38412 6972 38418
rect 6920 38354 6972 38360
rect 6932 37942 6960 38354
rect 6920 37936 6972 37942
rect 6920 37878 6972 37884
rect 6644 37664 6696 37670
rect 6644 37606 6696 37612
rect 6552 37256 6604 37262
rect 6552 37198 6604 37204
rect 6564 36922 6592 37198
rect 6552 36916 6604 36922
rect 6552 36858 6604 36864
rect 6104 36502 6224 36530
rect 6000 35828 6052 35834
rect 6000 35770 6052 35776
rect 5816 35624 5868 35630
rect 5816 35566 5868 35572
rect 5828 34066 5856 35566
rect 6012 34678 6040 35770
rect 6092 35148 6144 35154
rect 6092 35090 6144 35096
rect 6000 34672 6052 34678
rect 6000 34614 6052 34620
rect 6104 34610 6132 35090
rect 6092 34604 6144 34610
rect 6092 34546 6144 34552
rect 5816 34060 5868 34066
rect 5816 34002 5868 34008
rect 6196 33810 6224 36502
rect 6920 35692 6972 35698
rect 6920 35634 6972 35640
rect 6932 35018 6960 35634
rect 7024 35034 7052 41958
rect 7116 36310 7144 43590
rect 7208 40186 7236 45902
rect 7300 45082 7328 52430
rect 7288 45076 7340 45082
rect 7288 45018 7340 45024
rect 7288 44736 7340 44742
rect 7288 44678 7340 44684
rect 7300 44418 7328 44678
rect 7392 44538 7420 53479
rect 7564 53100 7616 53106
rect 7564 53042 7616 53048
rect 7472 50856 7524 50862
rect 7472 50798 7524 50804
rect 7484 46714 7512 50798
rect 7576 48006 7604 53042
rect 7760 52562 7788 56200
rect 7852 54262 7880 56222
rect 8036 56114 8064 56222
rect 8114 56200 8170 57000
rect 8482 56200 8538 57000
rect 8850 56200 8906 57000
rect 9218 56200 9274 57000
rect 9586 56200 9642 57000
rect 9954 56200 10010 57000
rect 10322 56200 10378 57000
rect 10690 56200 10746 57000
rect 11058 56200 11114 57000
rect 11426 56200 11482 57000
rect 11794 56200 11850 57000
rect 12162 56200 12218 57000
rect 12530 56200 12586 57000
rect 12898 56200 12954 57000
rect 13266 56200 13322 57000
rect 13634 56200 13690 57000
rect 14002 56200 14058 57000
rect 14370 56200 14426 57000
rect 14476 56222 14688 56250
rect 8128 56114 8156 56200
rect 8036 56086 8156 56114
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 7840 54256 7892 54262
rect 7840 54198 7892 54204
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7748 52556 7800 52562
rect 7748 52498 7800 52504
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 8496 51950 8524 56200
rect 8864 53650 8892 56200
rect 8852 53644 8904 53650
rect 8852 53586 8904 53592
rect 8668 53576 8720 53582
rect 8668 53518 8720 53524
rect 8576 52488 8628 52494
rect 8576 52430 8628 52436
rect 8484 51944 8536 51950
rect 8484 51886 8536 51892
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7656 50924 7708 50930
rect 7656 50866 7708 50872
rect 7840 50924 7892 50930
rect 7840 50866 7892 50872
rect 7564 48000 7616 48006
rect 7564 47942 7616 47948
rect 7472 46708 7524 46714
rect 7472 46650 7524 46656
rect 7564 46572 7616 46578
rect 7564 46514 7616 46520
rect 7380 44532 7432 44538
rect 7380 44474 7432 44480
rect 7300 44402 7420 44418
rect 7300 44396 7432 44402
rect 7300 44390 7380 44396
rect 7380 44338 7432 44344
rect 7472 44396 7524 44402
rect 7472 44338 7524 44344
rect 7288 40384 7340 40390
rect 7288 40326 7340 40332
rect 7196 40180 7248 40186
rect 7196 40122 7248 40128
rect 7300 39370 7328 40326
rect 7392 39953 7420 44338
rect 7378 39944 7434 39953
rect 7378 39879 7434 39888
rect 7288 39364 7340 39370
rect 7288 39306 7340 39312
rect 7300 39098 7328 39306
rect 7288 39092 7340 39098
rect 7288 39034 7340 39040
rect 7196 38548 7248 38554
rect 7196 38490 7248 38496
rect 7208 38214 7236 38490
rect 7380 38276 7432 38282
rect 7380 38218 7432 38224
rect 7196 38208 7248 38214
rect 7196 38150 7248 38156
rect 7392 37806 7420 38218
rect 7380 37800 7432 37806
rect 7380 37742 7432 37748
rect 7484 36922 7512 44338
rect 7576 42634 7604 46514
rect 7668 46102 7696 50866
rect 7748 49836 7800 49842
rect 7748 49778 7800 49784
rect 7656 46096 7708 46102
rect 7656 46038 7708 46044
rect 7760 43450 7788 49778
rect 7852 44538 7880 50866
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 7840 44532 7892 44538
rect 7840 44474 7892 44480
rect 8484 43784 8536 43790
rect 8484 43726 8536 43732
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 7748 43444 7800 43450
rect 7748 43386 7800 43392
rect 7656 43308 7708 43314
rect 7656 43250 7708 43256
rect 8392 43308 8444 43314
rect 8392 43250 8444 43256
rect 7564 42628 7616 42634
rect 7564 42570 7616 42576
rect 7564 41472 7616 41478
rect 7564 41414 7616 41420
rect 7576 40730 7604 41414
rect 7564 40724 7616 40730
rect 7564 40666 7616 40672
rect 7576 38282 7604 40666
rect 7564 38276 7616 38282
rect 7564 38218 7616 38224
rect 7564 37936 7616 37942
rect 7564 37878 7616 37884
rect 7576 37806 7604 37878
rect 7564 37800 7616 37806
rect 7564 37742 7616 37748
rect 7576 37194 7604 37742
rect 7564 37188 7616 37194
rect 7564 37130 7616 37136
rect 7472 36916 7524 36922
rect 7472 36858 7524 36864
rect 7576 36854 7604 37130
rect 7564 36848 7616 36854
rect 7564 36790 7616 36796
rect 7380 36644 7432 36650
rect 7380 36586 7432 36592
rect 7104 36304 7156 36310
rect 7104 36246 7156 36252
rect 7392 36174 7420 36586
rect 7668 36378 7696 43250
rect 8404 42566 8432 43250
rect 8392 42560 8444 42566
rect 8392 42502 8444 42508
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 8116 42356 8168 42362
rect 8116 42298 8168 42304
rect 7748 42152 7800 42158
rect 7748 42094 7800 42100
rect 7760 41818 7788 42094
rect 8128 41818 8156 42298
rect 7748 41812 7800 41818
rect 7748 41754 7800 41760
rect 7840 41812 7892 41818
rect 7840 41754 7892 41760
rect 8116 41812 8168 41818
rect 8116 41754 8168 41760
rect 7748 41540 7800 41546
rect 7748 41482 7800 41488
rect 7760 38554 7788 41482
rect 7852 41274 7880 41754
rect 8300 41744 8352 41750
rect 8300 41686 8352 41692
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7840 41268 7892 41274
rect 7840 41210 7892 41216
rect 7852 40066 7880 41210
rect 8312 40390 8340 41686
rect 8300 40384 8352 40390
rect 8300 40326 8352 40332
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 7852 40050 7972 40066
rect 7852 40044 7984 40050
rect 7852 40038 7932 40044
rect 7932 39986 7984 39992
rect 7840 39976 7892 39982
rect 7840 39918 7892 39924
rect 7748 38548 7800 38554
rect 7748 38490 7800 38496
rect 7852 38418 7880 39918
rect 8300 39296 8352 39302
rect 8300 39238 8352 39244
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7840 38412 7892 38418
rect 7840 38354 7892 38360
rect 8312 38350 8340 39238
rect 8300 38344 8352 38350
rect 8206 38312 8262 38321
rect 8300 38286 8352 38292
rect 8206 38247 8262 38256
rect 8220 38214 8248 38247
rect 8208 38208 8260 38214
rect 8208 38150 8260 38156
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 7840 37800 7892 37806
rect 7760 37760 7840 37788
rect 7656 36372 7708 36378
rect 7656 36314 7708 36320
rect 7564 36236 7616 36242
rect 7564 36178 7616 36184
rect 7380 36168 7432 36174
rect 7380 36110 7432 36116
rect 7288 35828 7340 35834
rect 7288 35770 7340 35776
rect 6920 35012 6972 35018
rect 7024 35006 7144 35034
rect 6920 34954 6972 34960
rect 6932 34898 6960 34954
rect 7012 34944 7064 34950
rect 6932 34892 7012 34898
rect 6932 34886 7064 34892
rect 6932 34870 7052 34886
rect 6932 34678 6960 34870
rect 6920 34672 6972 34678
rect 6920 34614 6972 34620
rect 6932 34202 6960 34614
rect 6920 34196 6972 34202
rect 6920 34138 6972 34144
rect 6932 33998 6960 34138
rect 6920 33992 6972 33998
rect 6920 33934 6972 33940
rect 6196 33782 6316 33810
rect 6184 32428 6236 32434
rect 6184 32370 6236 32376
rect 6196 31890 6224 32370
rect 6184 31884 6236 31890
rect 6184 31826 6236 31832
rect 5724 31136 5776 31142
rect 5724 31078 5776 31084
rect 4620 30796 4672 30802
rect 4620 30738 4672 30744
rect 4252 29844 4304 29850
rect 4252 29786 4304 29792
rect 4068 28620 4120 28626
rect 4068 28562 4120 28568
rect 3988 28478 4108 28506
rect 3976 28416 4028 28422
rect 3976 28358 4028 28364
rect 3792 28212 3844 28218
rect 3792 28154 3844 28160
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3424 27124 3476 27130
rect 3424 27066 3476 27072
rect 3424 26988 3476 26994
rect 3424 26930 3476 26936
rect 3332 25764 3384 25770
rect 3332 25706 3384 25712
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 3436 24410 3464 26930
rect 3516 25968 3568 25974
rect 3516 25910 3568 25916
rect 3424 24404 3476 24410
rect 3424 24346 3476 24352
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2044 23316 2096 23322
rect 2044 23258 2096 23264
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 3436 23186 3464 24346
rect 3528 24206 3556 25910
rect 3620 25838 3648 28018
rect 3608 25832 3660 25838
rect 3608 25774 3660 25780
rect 3988 25158 4016 28358
rect 4080 26586 4108 28478
rect 4344 27056 4396 27062
rect 4344 26998 4396 27004
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 4080 25974 4108 26522
rect 4068 25968 4120 25974
rect 4068 25910 4120 25916
rect 4252 25696 4304 25702
rect 4252 25638 4304 25644
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3988 24206 4016 24550
rect 3516 24200 3568 24206
rect 3516 24142 3568 24148
rect 3976 24200 4028 24206
rect 3976 24142 4028 24148
rect 3988 23662 4016 24142
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3884 23316 3936 23322
rect 3884 23258 3936 23264
rect 2872 23180 2924 23186
rect 2792 23140 2872 23168
rect 1860 21548 1912 21554
rect 1860 21490 1912 21496
rect 1308 21480 1360 21486
rect 1308 21422 1360 21428
rect 1320 21185 1348 21422
rect 1306 21176 1362 21185
rect 1306 21111 1362 21120
rect 2792 20890 2820 23140
rect 2872 23122 2924 23128
rect 3424 23180 3476 23186
rect 3424 23122 3476 23128
rect 3700 23112 3752 23118
rect 3700 23054 3752 23060
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2884 21146 2912 22578
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 2792 20874 2912 20890
rect 1860 20868 1912 20874
rect 2792 20868 2924 20874
rect 2792 20862 2872 20868
rect 1860 20810 1912 20816
rect 2872 20810 2924 20816
rect 1768 20800 1820 20806
rect 1768 20742 1820 20748
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 1308 18828 1360 18834
rect 1308 18770 1360 18776
rect 1320 18737 1348 18770
rect 1306 18728 1362 18737
rect 1306 18663 1362 18672
rect 1504 16590 1532 19450
rect 1780 18766 1808 20742
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1492 16584 1544 16590
rect 1492 16526 1544 16532
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 13938 1808 15846
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1308 13864 1360 13870
rect 1306 13832 1308 13841
rect 1360 13832 1362 13841
rect 1306 13767 1362 13776
rect 1872 6458 1900 20810
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3620 19514 3648 21422
rect 3712 20942 3740 23054
rect 3792 23044 3844 23050
rect 3792 22986 3844 22992
rect 3804 21418 3832 22986
rect 3792 21412 3844 21418
rect 3792 21354 3844 21360
rect 3700 20936 3752 20942
rect 3700 20878 3752 20884
rect 3608 19508 3660 19514
rect 3608 19450 3660 19456
rect 3896 19378 3924 23258
rect 4080 21486 4108 25230
rect 4264 24954 4292 25638
rect 4252 24948 4304 24954
rect 4252 24890 4304 24896
rect 4264 24274 4292 24890
rect 4252 24268 4304 24274
rect 4252 24210 4304 24216
rect 4252 24132 4304 24138
rect 4252 24074 4304 24080
rect 4160 23792 4212 23798
rect 4160 23734 4212 23740
rect 4172 22522 4200 23734
rect 4264 22964 4292 24074
rect 4356 23118 4384 26998
rect 4528 26852 4580 26858
rect 4528 26794 4580 26800
rect 4436 24404 4488 24410
rect 4436 24346 4488 24352
rect 4448 23798 4476 24346
rect 4436 23792 4488 23798
rect 4436 23734 4488 23740
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4264 22936 4476 22964
rect 4172 22494 4384 22522
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 3976 21412 4028 21418
rect 3976 21354 4028 21360
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3792 18896 3844 18902
rect 3792 18838 3844 18844
rect 3804 18222 3832 18838
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3700 17264 3752 17270
rect 3700 17206 3752 17212
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2502 16552 2558 16561
rect 2502 16487 2558 16496
rect 2516 16182 2544 16487
rect 2504 16176 2556 16182
rect 2504 16118 2556 16124
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3620 8945 3648 9046
rect 3606 8936 3662 8945
rect 3606 8871 3662 8880
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1688 5030 1716 5170
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1504 3534 1532 3878
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1688 800 1716 4966
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1780 4146 1808 4422
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1872 3738 1900 5578
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2056 800 2084 3470
rect 2148 3058 2176 5578
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2332 2650 2360 5102
rect 2424 4146 2452 6258
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2516 5710 2544 6054
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2792 3618 2820 6190
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 3344 5914 3372 6258
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3068 5370 3096 5646
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2884 3738 2912 5170
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2792 3590 2912 3618
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2424 800 2452 2994
rect 2792 2990 2820 3470
rect 2884 3194 2912 3590
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 2792 800 2820 2926
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 3344 2632 3372 2926
rect 3160 2604 3372 2632
rect 3160 800 3188 2604
rect 3436 1601 3464 4558
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3422 1592 3478 1601
rect 3422 1527 3478 1536
rect 3528 800 3556 2450
rect 3620 2378 3648 5510
rect 3712 4049 3740 17206
rect 3804 16046 3832 18158
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3896 11665 3924 19314
rect 3988 17270 4016 21354
rect 4264 20942 4292 22374
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 3976 17264 4028 17270
rect 3976 17206 4028 17212
rect 4080 16561 4108 20878
rect 4356 20534 4384 22494
rect 4448 21894 4476 22936
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 4436 21548 4488 21554
rect 4436 21490 4488 21496
rect 4344 20528 4396 20534
rect 4344 20470 4396 20476
rect 4448 19514 4476 21490
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4540 19446 4568 26794
rect 4528 19440 4580 19446
rect 4528 19382 4580 19388
rect 4632 17202 4660 30738
rect 6288 30326 6316 33782
rect 6932 33658 6960 33934
rect 6920 33652 6972 33658
rect 6920 33594 6972 33600
rect 6932 32910 6960 33594
rect 7116 33318 7144 35006
rect 7196 34740 7248 34746
rect 7196 34682 7248 34688
rect 7104 33312 7156 33318
rect 7104 33254 7156 33260
rect 6920 32904 6972 32910
rect 6920 32846 6972 32852
rect 7208 31890 7236 34682
rect 7196 31884 7248 31890
rect 7196 31826 7248 31832
rect 6276 30320 6328 30326
rect 6276 30262 6328 30268
rect 7208 29714 7236 31826
rect 7196 29708 7248 29714
rect 7196 29650 7248 29656
rect 7300 29646 7328 35770
rect 7392 35290 7420 36110
rect 7472 36032 7524 36038
rect 7472 35974 7524 35980
rect 7380 35284 7432 35290
rect 7380 35226 7432 35232
rect 7484 33114 7512 35974
rect 7472 33108 7524 33114
rect 7472 33050 7524 33056
rect 7576 33046 7604 36178
rect 7760 34202 7788 37760
rect 7840 37742 7892 37748
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 7840 36780 7892 36786
rect 7840 36722 7892 36728
rect 7852 34202 7880 36722
rect 8404 36122 8432 42502
rect 8496 40934 8524 43726
rect 8588 43450 8616 52430
rect 8680 50522 8708 53518
rect 9232 53174 9260 56200
rect 9600 53564 9628 56200
rect 9968 54330 9996 56200
rect 9956 54324 10008 54330
rect 9956 54266 10008 54272
rect 9956 54188 10008 54194
rect 9956 54130 10008 54136
rect 9600 53536 9812 53564
rect 9220 53168 9272 53174
rect 9220 53110 9272 53116
rect 9312 53100 9364 53106
rect 9312 53042 9364 53048
rect 9128 52080 9180 52086
rect 9128 52022 9180 52028
rect 8668 50516 8720 50522
rect 8668 50458 8720 50464
rect 9036 49904 9088 49910
rect 9036 49846 9088 49852
rect 8852 49768 8904 49774
rect 8852 49710 8904 49716
rect 8864 45558 8892 49710
rect 9048 46986 9076 49846
rect 9140 47802 9168 52022
rect 9220 51400 9272 51406
rect 9220 51342 9272 51348
rect 9128 47796 9180 47802
rect 9128 47738 9180 47744
rect 9036 46980 9088 46986
rect 9036 46922 9088 46928
rect 9232 46170 9260 51342
rect 9324 49910 9352 53042
rect 9588 52488 9640 52494
rect 9588 52430 9640 52436
rect 9600 50998 9628 52430
rect 9680 52012 9732 52018
rect 9680 51954 9732 51960
rect 9588 50992 9640 50998
rect 9588 50934 9640 50940
rect 9404 50312 9456 50318
rect 9404 50254 9456 50260
rect 9312 49904 9364 49910
rect 9312 49846 9364 49852
rect 9220 46164 9272 46170
rect 9220 46106 9272 46112
rect 8852 45552 8904 45558
rect 8852 45494 8904 45500
rect 8668 44736 8720 44742
rect 8668 44678 8720 44684
rect 8576 43444 8628 43450
rect 8576 43386 8628 43392
rect 8588 42906 8616 43386
rect 8576 42900 8628 42906
rect 8576 42842 8628 42848
rect 8576 42764 8628 42770
rect 8576 42706 8628 42712
rect 8588 41478 8616 42706
rect 8576 41472 8628 41478
rect 8576 41414 8628 41420
rect 8484 40928 8536 40934
rect 8484 40870 8536 40876
rect 8482 40760 8538 40769
rect 8482 40695 8484 40704
rect 8536 40695 8538 40704
rect 8484 40666 8536 40672
rect 8484 39908 8536 39914
rect 8484 39850 8536 39856
rect 8496 39642 8524 39850
rect 8484 39636 8536 39642
rect 8484 39578 8536 39584
rect 8576 38480 8628 38486
rect 8576 38422 8628 38428
rect 8484 38208 8536 38214
rect 8484 38150 8536 38156
rect 8496 36922 8524 38150
rect 8588 37466 8616 38422
rect 8680 37466 8708 44678
rect 8864 43246 8892 45494
rect 9220 45484 9272 45490
rect 9220 45426 9272 45432
rect 8944 44396 8996 44402
rect 8944 44338 8996 44344
rect 8852 43240 8904 43246
rect 8852 43182 8904 43188
rect 8864 42906 8892 43182
rect 8852 42900 8904 42906
rect 8852 42842 8904 42848
rect 8852 42560 8904 42566
rect 8852 42502 8904 42508
rect 8864 42242 8892 42502
rect 8772 42226 8892 42242
rect 8772 42220 8904 42226
rect 8772 42214 8852 42220
rect 8772 41750 8800 42214
rect 8852 42162 8904 42168
rect 8956 42106 8984 44338
rect 9232 42770 9260 45426
rect 9416 43994 9444 50254
rect 9496 46028 9548 46034
rect 9496 45970 9548 45976
rect 9404 43988 9456 43994
rect 9404 43930 9456 43936
rect 9404 43852 9456 43858
rect 9404 43794 9456 43800
rect 9312 42900 9364 42906
rect 9312 42842 9364 42848
rect 9220 42764 9272 42770
rect 9220 42706 9272 42712
rect 9232 42362 9260 42706
rect 9220 42356 9272 42362
rect 9220 42298 9272 42304
rect 9128 42220 9180 42226
rect 9128 42162 9180 42168
rect 8864 42078 8984 42106
rect 8760 41744 8812 41750
rect 8760 41686 8812 41692
rect 8760 40112 8812 40118
rect 8760 40054 8812 40060
rect 8576 37460 8628 37466
rect 8576 37402 8628 37408
rect 8668 37460 8720 37466
rect 8668 37402 8720 37408
rect 8668 37324 8720 37330
rect 8668 37266 8720 37272
rect 8484 36916 8536 36922
rect 8484 36858 8536 36864
rect 8680 36582 8708 37266
rect 8668 36576 8720 36582
rect 8668 36518 8720 36524
rect 8574 36136 8630 36145
rect 8404 36094 8574 36122
rect 8574 36071 8630 36080
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 8588 35834 8616 36071
rect 8680 35873 8708 36518
rect 8666 35864 8722 35873
rect 8576 35828 8628 35834
rect 8666 35799 8722 35808
rect 8576 35770 8628 35776
rect 8576 35488 8628 35494
rect 8576 35430 8628 35436
rect 8300 34944 8352 34950
rect 8300 34886 8352 34892
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 8312 34746 8340 34886
rect 8300 34740 8352 34746
rect 8300 34682 8352 34688
rect 8484 34672 8536 34678
rect 8484 34614 8536 34620
rect 7748 34196 7800 34202
rect 7748 34138 7800 34144
rect 7840 34196 7892 34202
rect 7840 34138 7892 34144
rect 7656 33924 7708 33930
rect 7656 33866 7708 33872
rect 7564 33040 7616 33046
rect 7564 32982 7616 32988
rect 7576 32298 7604 32982
rect 7564 32292 7616 32298
rect 7564 32234 7616 32240
rect 7668 31482 7696 33866
rect 7760 33862 7788 34138
rect 8496 34134 8524 34614
rect 8588 34610 8616 35430
rect 8680 35170 8708 35799
rect 8772 35290 8800 40054
rect 8864 38593 8892 42078
rect 9140 41546 9168 42162
rect 9232 41682 9260 42298
rect 9220 41676 9272 41682
rect 9220 41618 9272 41624
rect 9324 41562 9352 42842
rect 9416 42770 9444 43794
rect 9508 43314 9536 45970
rect 9692 44538 9720 51954
rect 9784 51950 9812 53536
rect 9772 51944 9824 51950
rect 9772 51886 9824 51892
rect 9968 51610 9996 54130
rect 10336 53038 10364 56200
rect 10324 53032 10376 53038
rect 10324 52974 10376 52980
rect 10704 52562 10732 56200
rect 11072 53650 11100 56200
rect 11440 54262 11468 56200
rect 11428 54256 11480 54262
rect 11428 54198 11480 54204
rect 11612 54188 11664 54194
rect 11612 54130 11664 54136
rect 11244 54120 11296 54126
rect 11244 54062 11296 54068
rect 11060 53644 11112 53650
rect 11060 53586 11112 53592
rect 10692 52556 10744 52562
rect 10692 52498 10744 52504
rect 10876 52012 10928 52018
rect 10876 51954 10928 51960
rect 10416 51876 10468 51882
rect 10416 51818 10468 51824
rect 9956 51604 10008 51610
rect 9956 51546 10008 51552
rect 9864 49972 9916 49978
rect 9864 49914 9916 49920
rect 9876 47258 9904 49914
rect 9864 47252 9916 47258
rect 9864 47194 9916 47200
rect 9876 45642 9904 47194
rect 10048 46912 10100 46918
rect 10048 46854 10100 46860
rect 9784 45614 9904 45642
rect 9784 45558 9812 45614
rect 9772 45552 9824 45558
rect 9772 45494 9824 45500
rect 9876 45422 9904 45614
rect 10060 45558 10088 46854
rect 10048 45552 10100 45558
rect 10048 45494 10100 45500
rect 9864 45416 9916 45422
rect 9864 45358 9916 45364
rect 10060 45286 10088 45494
rect 10048 45280 10100 45286
rect 10048 45222 10100 45228
rect 9772 44736 9824 44742
rect 9772 44678 9824 44684
rect 9680 44532 9732 44538
rect 9680 44474 9732 44480
rect 9588 43444 9640 43450
rect 9588 43386 9640 43392
rect 9496 43308 9548 43314
rect 9496 43250 9548 43256
rect 9508 42906 9536 43250
rect 9496 42900 9548 42906
rect 9496 42842 9548 42848
rect 9404 42764 9456 42770
rect 9404 42706 9456 42712
rect 9128 41540 9180 41546
rect 9128 41482 9180 41488
rect 9232 41534 9352 41562
rect 9128 41200 9180 41206
rect 9128 41142 9180 41148
rect 9036 40928 9088 40934
rect 9036 40870 9088 40876
rect 8850 38584 8906 38593
rect 8850 38519 8906 38528
rect 8852 37392 8904 37398
rect 8852 37334 8904 37340
rect 8760 35284 8812 35290
rect 8760 35226 8812 35232
rect 8680 35142 8800 35170
rect 8668 35012 8720 35018
rect 8668 34954 8720 34960
rect 8576 34604 8628 34610
rect 8576 34546 8628 34552
rect 8484 34128 8536 34134
rect 8484 34070 8536 34076
rect 7748 33856 7800 33862
rect 7748 33798 7800 33804
rect 8392 33856 8444 33862
rect 8392 33798 8444 33804
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 8300 33380 8352 33386
rect 8300 33322 8352 33328
rect 8312 32978 8340 33322
rect 8300 32972 8352 32978
rect 8300 32914 8352 32920
rect 7748 32836 7800 32842
rect 7748 32778 7800 32784
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 7760 29850 7788 32778
rect 7840 32768 7892 32774
rect 7840 32710 7892 32716
rect 7852 32570 7880 32710
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 7840 32564 7892 32570
rect 7840 32506 7892 32512
rect 8312 32026 8340 32914
rect 8404 32366 8432 33798
rect 8392 32360 8444 32366
rect 8392 32302 8444 32308
rect 8404 32026 8432 32302
rect 8300 32020 8352 32026
rect 8300 31962 8352 31968
rect 8392 32020 8444 32026
rect 8392 31962 8444 31968
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 8680 31482 8708 34954
rect 8668 31476 8720 31482
rect 8668 31418 8720 31424
rect 8772 31346 8800 35142
rect 7840 31340 7892 31346
rect 7840 31282 7892 31288
rect 8760 31340 8812 31346
rect 8760 31282 8812 31288
rect 7852 30802 7880 31282
rect 8668 31204 8720 31210
rect 8668 31146 8720 31152
rect 8760 31204 8812 31210
rect 8760 31146 8812 31152
rect 7840 30796 7892 30802
rect 7840 30738 7892 30744
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 7656 29844 7708 29850
rect 7656 29786 7708 29792
rect 7748 29844 7800 29850
rect 7748 29786 7800 29792
rect 7288 29640 7340 29646
rect 7288 29582 7340 29588
rect 5264 29572 5316 29578
rect 5264 29514 5316 29520
rect 7012 29572 7064 29578
rect 7012 29514 7064 29520
rect 5172 28620 5224 28626
rect 5172 28562 5224 28568
rect 5080 23180 5132 23186
rect 5080 23122 5132 23128
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4724 21554 4752 21830
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4724 17678 4752 21490
rect 5092 20058 5120 23122
rect 5080 20052 5132 20058
rect 5080 19994 5132 20000
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4066 16552 4122 16561
rect 4066 16487 4122 16496
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 3882 11656 3938 11665
rect 3882 11591 3938 11600
rect 4080 6497 4108 15982
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4066 6488 4122 6497
rect 4356 6458 4384 7754
rect 4066 6423 4122 6432
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 3790 5808 3846 5817
rect 3790 5743 3846 5752
rect 3804 5370 3832 5743
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3896 4162 3924 5510
rect 4172 4826 4200 5850
rect 4448 5370 4476 9454
rect 4908 9110 4936 18770
rect 5184 18766 5212 28562
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5276 18290 5304 29514
rect 6552 29096 6604 29102
rect 6552 29038 6604 29044
rect 6564 28626 6592 29038
rect 6552 28620 6604 28626
rect 6552 28562 6604 28568
rect 6564 27538 6592 28562
rect 6552 27532 6604 27538
rect 6552 27474 6604 27480
rect 6564 26994 6592 27474
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 6564 26466 6592 26930
rect 6472 26450 6592 26466
rect 6460 26444 6592 26450
rect 6512 26438 6592 26444
rect 6460 26386 6512 26392
rect 6184 25832 6236 25838
rect 6184 25774 6236 25780
rect 5448 25696 5500 25702
rect 5448 25638 5500 25644
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 4986 18184 5042 18193
rect 4986 18119 5042 18128
rect 5000 18086 5028 18119
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 5000 5846 5028 18022
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 4988 5840 5040 5846
rect 4988 5782 5040 5788
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3804 4134 3924 4162
rect 3698 4040 3754 4049
rect 3698 3975 3754 3984
rect 3804 2514 3832 4134
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 3896 800 3924 3946
rect 3988 2650 4016 4558
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4172 3194 4200 3470
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4632 3058 4660 3334
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4816 2922 4844 5510
rect 5184 5370 5212 16390
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3516 4936 3878
rect 5000 3738 5028 4558
rect 5368 4146 5396 4966
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4988 3528 5040 3534
rect 4908 3488 4988 3516
rect 4988 3470 5040 3476
rect 4804 2916 4856 2922
rect 4804 2858 4856 2864
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4724 2446 4752 2790
rect 4712 2440 4764 2446
rect 4632 2400 4712 2428
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 4080 2258 4108 2314
rect 4080 2230 4292 2258
rect 4264 800 4292 2230
rect 4632 800 4660 2400
rect 4712 2382 4764 2388
rect 5000 800 5028 3470
rect 5368 800 5396 4082
rect 5460 4010 5488 25638
rect 6000 24744 6052 24750
rect 6000 24686 6052 24692
rect 6012 23866 6040 24686
rect 6196 24410 6224 25774
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6368 24336 6420 24342
rect 6368 24278 6420 24284
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 5724 23520 5776 23526
rect 5724 23462 5776 23468
rect 5736 23186 5764 23462
rect 5724 23180 5776 23186
rect 5724 23122 5776 23128
rect 5736 20602 5764 23122
rect 6012 22574 6040 23802
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 5736 20466 5764 20538
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5736 19922 5764 20402
rect 5828 20262 5856 21286
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5828 13530 5856 20198
rect 5920 18834 5948 21286
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 6288 17882 6316 19314
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5920 4826 5948 5714
rect 6380 5574 6408 24278
rect 6472 23186 6500 26386
rect 6736 26036 6788 26042
rect 6736 25978 6788 25984
rect 6460 23180 6512 23186
rect 6460 23122 6512 23128
rect 6460 20528 6512 20534
rect 6460 20470 6512 20476
rect 6472 20262 6500 20470
rect 6460 20256 6512 20262
rect 6460 20198 6512 20204
rect 6472 19786 6500 20198
rect 6460 19780 6512 19786
rect 6460 19722 6512 19728
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6564 17134 6592 19314
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6564 16640 6592 17070
rect 6644 16652 6696 16658
rect 6564 16612 6644 16640
rect 6644 16594 6696 16600
rect 6656 16114 6684 16594
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6564 9450 6592 12786
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6656 8106 6684 12854
rect 6564 8090 6684 8106
rect 6552 8084 6684 8090
rect 6604 8078 6684 8084
rect 6552 8026 6604 8032
rect 6564 7886 6592 8026
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3058 5580 3878
rect 5736 3738 5764 4558
rect 6012 4146 6040 5170
rect 6748 4826 6776 25978
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6932 24070 6960 24550
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 6840 19310 6868 23802
rect 6932 23798 6960 24006
rect 6920 23792 6972 23798
rect 6920 23734 6972 23740
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6932 17864 6960 22374
rect 6840 17836 6960 17864
rect 6840 16674 6868 17836
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6932 17134 6960 17682
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6932 16794 6960 17070
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6840 16646 6960 16674
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6840 8090 6868 13262
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6564 4146 6592 4422
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5736 2310 5764 3470
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 5736 800 5764 2246
rect 6104 800 6132 2994
rect 6564 2774 6592 4082
rect 6932 4010 6960 16646
rect 7024 4826 7052 29514
rect 7668 29510 7696 29786
rect 7840 29640 7892 29646
rect 7840 29582 7892 29588
rect 7656 29504 7708 29510
rect 7656 29446 7708 29452
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 7116 25226 7144 26522
rect 7668 25514 7696 29446
rect 7748 29300 7800 29306
rect 7748 29242 7800 29248
rect 7760 26586 7788 29242
rect 7852 27606 7880 29582
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 8116 28756 8168 28762
rect 8116 28698 8168 28704
rect 8128 28490 8156 28698
rect 8116 28484 8168 28490
rect 8168 28444 8340 28472
rect 8116 28426 8168 28432
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 8312 27606 8340 28444
rect 8576 28008 8628 28014
rect 8576 27950 8628 27956
rect 7840 27600 7892 27606
rect 7840 27542 7892 27548
rect 8300 27600 8352 27606
rect 8300 27542 8352 27548
rect 7852 26926 7880 27542
rect 8312 27402 8340 27542
rect 8300 27396 8352 27402
rect 8300 27338 8352 27344
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 8312 27062 8340 27338
rect 8116 27056 8168 27062
rect 8116 26998 8168 27004
rect 8300 27056 8352 27062
rect 8300 26998 8352 27004
rect 7840 26920 7892 26926
rect 7840 26862 7892 26868
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7852 25922 7880 26862
rect 8128 26314 8156 26998
rect 8300 26852 8352 26858
rect 8300 26794 8352 26800
rect 8312 26450 8340 26794
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 8116 26308 8168 26314
rect 8116 26250 8168 26256
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 8496 25974 8524 26250
rect 7576 25486 7696 25514
rect 7760 25894 7880 25922
rect 8484 25968 8536 25974
rect 8484 25910 8536 25916
rect 7104 25220 7156 25226
rect 7104 25162 7156 25168
rect 7116 24886 7144 25162
rect 7104 24880 7156 24886
rect 7104 24822 7156 24828
rect 7576 24818 7604 25486
rect 7656 25356 7708 25362
rect 7656 25298 7708 25304
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7472 24608 7524 24614
rect 7472 24550 7524 24556
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7116 21690 7144 24142
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7300 21146 7328 22510
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7392 20618 7420 23122
rect 7484 22250 7512 24550
rect 7668 23662 7696 25298
rect 7760 24818 7788 25894
rect 7840 25832 7892 25838
rect 7840 25774 7892 25780
rect 7852 24954 7880 25774
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7840 24948 7892 24954
rect 7840 24890 7892 24896
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 8116 24744 8168 24750
rect 8168 24704 8340 24732
rect 8116 24686 8168 24692
rect 7840 24064 7892 24070
rect 7840 24006 7892 24012
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7576 23322 7604 23598
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7576 22574 7604 23258
rect 7852 23254 7880 24006
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7748 23044 7800 23050
rect 7748 22986 7800 22992
rect 7564 22568 7616 22574
rect 7616 22516 7696 22522
rect 7564 22510 7696 22516
rect 7576 22494 7696 22510
rect 7484 22222 7604 22250
rect 7472 22160 7524 22166
rect 7472 22102 7524 22108
rect 7484 21418 7512 22102
rect 7472 21412 7524 21418
rect 7472 21354 7524 21360
rect 7300 20590 7420 20618
rect 7300 20534 7328 20590
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 7300 20262 7328 20470
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7300 19854 7328 20198
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7300 19446 7328 19790
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7288 19440 7340 19446
rect 7288 19382 7340 19388
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7116 13258 7144 18158
rect 7392 17882 7420 19654
rect 7576 18426 7604 22222
rect 7668 21622 7696 22494
rect 7656 21616 7708 21622
rect 7656 21558 7708 21564
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7668 19786 7696 21422
rect 7760 21010 7788 22986
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7852 21418 7880 22578
rect 8312 22094 8340 24704
rect 8404 24682 8432 25230
rect 8392 24676 8444 24682
rect 8392 24618 8444 24624
rect 8496 24070 8524 25910
rect 8588 25770 8616 27950
rect 8680 26926 8708 31146
rect 8772 30598 8800 31146
rect 8760 30592 8812 30598
rect 8760 30534 8812 30540
rect 8668 26920 8720 26926
rect 8668 26862 8720 26868
rect 8680 26314 8708 26862
rect 8668 26308 8720 26314
rect 8668 26250 8720 26256
rect 8576 25764 8628 25770
rect 8576 25706 8628 25712
rect 8576 25152 8628 25158
rect 8576 25094 8628 25100
rect 8588 24342 8616 25094
rect 8576 24336 8628 24342
rect 8576 24278 8628 24284
rect 8484 24064 8536 24070
rect 8484 24006 8536 24012
rect 8496 23798 8524 24006
rect 8484 23792 8536 23798
rect 8484 23734 8536 23740
rect 8588 23662 8616 24278
rect 8576 23656 8628 23662
rect 8576 23598 8628 23604
rect 8312 22066 8432 22094
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7840 21412 7892 21418
rect 7840 21354 7892 21360
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7748 20868 7800 20874
rect 7748 20810 7800 20816
rect 7656 19780 7708 19786
rect 7656 19722 7708 19728
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7760 18290 7788 20810
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8312 19922 8340 20198
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8404 19378 8432 22066
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8588 20806 8616 21830
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8680 20466 8708 26250
rect 8772 25838 8800 30534
rect 8864 26042 8892 37334
rect 9048 36922 9076 40870
rect 9140 40390 9168 41142
rect 9232 40526 9260 41534
rect 9312 41472 9364 41478
rect 9312 41414 9364 41420
rect 9220 40520 9272 40526
rect 9220 40462 9272 40468
rect 9128 40384 9180 40390
rect 9128 40326 9180 40332
rect 9220 40384 9272 40390
rect 9220 40326 9272 40332
rect 9140 40186 9168 40326
rect 9128 40180 9180 40186
rect 9128 40122 9180 40128
rect 9232 39506 9260 40326
rect 9220 39500 9272 39506
rect 9220 39442 9272 39448
rect 9128 38752 9180 38758
rect 9128 38694 9180 38700
rect 9140 38418 9168 38694
rect 9128 38412 9180 38418
rect 9128 38354 9180 38360
rect 9220 38344 9272 38350
rect 9220 38286 9272 38292
rect 9128 38004 9180 38010
rect 9128 37946 9180 37952
rect 9036 36916 9088 36922
rect 9036 36858 9088 36864
rect 9140 36378 9168 37946
rect 9128 36372 9180 36378
rect 9128 36314 9180 36320
rect 9232 34066 9260 38286
rect 9324 37874 9352 41414
rect 9416 41274 9444 42706
rect 9600 42140 9628 43386
rect 9680 42628 9732 42634
rect 9680 42570 9732 42576
rect 9692 42362 9720 42570
rect 9680 42356 9732 42362
rect 9680 42298 9732 42304
rect 9508 42112 9628 42140
rect 9404 41268 9456 41274
rect 9404 41210 9456 41216
rect 9404 40588 9456 40594
rect 9404 40530 9456 40536
rect 9416 40186 9444 40530
rect 9508 40458 9536 42112
rect 9588 42016 9640 42022
rect 9640 41964 9720 41970
rect 9588 41958 9720 41964
rect 9600 41942 9720 41958
rect 9692 41750 9720 41942
rect 9680 41744 9732 41750
rect 9680 41686 9732 41692
rect 9588 40724 9640 40730
rect 9588 40666 9640 40672
rect 9600 40497 9628 40666
rect 9586 40488 9642 40497
rect 9496 40452 9548 40458
rect 9586 40423 9642 40432
rect 9496 40394 9548 40400
rect 9404 40180 9456 40186
rect 9404 40122 9456 40128
rect 9312 37868 9364 37874
rect 9312 37810 9364 37816
rect 9416 37330 9444 40122
rect 9508 39098 9536 40394
rect 9600 40390 9628 40423
rect 9588 40384 9640 40390
rect 9588 40326 9640 40332
rect 9496 39092 9548 39098
rect 9496 39034 9548 39040
rect 9680 38888 9732 38894
rect 9508 38836 9680 38842
rect 9508 38830 9732 38836
rect 9508 38826 9720 38830
rect 9496 38820 9720 38826
rect 9548 38814 9720 38820
rect 9496 38762 9548 38768
rect 9600 37942 9628 38814
rect 9588 37936 9640 37942
rect 9588 37878 9640 37884
rect 9404 37324 9456 37330
rect 9404 37266 9456 37272
rect 9784 36825 9812 44678
rect 10060 43722 10088 45222
rect 10048 43716 10100 43722
rect 10048 43658 10100 43664
rect 10060 43382 10088 43658
rect 10428 43450 10456 51818
rect 10692 49224 10744 49230
rect 10692 49166 10744 49172
rect 10508 46980 10560 46986
rect 10508 46922 10560 46928
rect 10520 45354 10548 46922
rect 10704 46170 10732 49166
rect 10784 49088 10836 49094
rect 10784 49030 10836 49036
rect 10796 46594 10824 49030
rect 10888 46714 10916 51954
rect 10876 46708 10928 46714
rect 10876 46650 10928 46656
rect 10796 46566 11008 46594
rect 10692 46164 10744 46170
rect 10692 46106 10744 46112
rect 10508 45348 10560 45354
rect 10508 45290 10560 45296
rect 10980 43654 11008 46566
rect 11060 46572 11112 46578
rect 11060 46514 11112 46520
rect 10968 43648 11020 43654
rect 10968 43590 11020 43596
rect 10416 43444 10468 43450
rect 10416 43386 10468 43392
rect 10048 43376 10100 43382
rect 10048 43318 10100 43324
rect 10060 41274 10088 43318
rect 10324 43308 10376 43314
rect 10324 43250 10376 43256
rect 10336 42566 10364 43250
rect 10324 42560 10376 42566
rect 10322 42528 10324 42537
rect 10876 42560 10928 42566
rect 10376 42528 10378 42537
rect 10876 42502 10928 42508
rect 10322 42463 10378 42472
rect 10140 42152 10192 42158
rect 10140 42094 10192 42100
rect 10048 41268 10100 41274
rect 10048 41210 10100 41216
rect 9864 38548 9916 38554
rect 9864 38490 9916 38496
rect 9770 36816 9826 36825
rect 9312 36780 9364 36786
rect 9770 36751 9826 36760
rect 9312 36722 9364 36728
rect 9220 34060 9272 34066
rect 9220 34002 9272 34008
rect 9324 33114 9352 36722
rect 9588 36712 9640 36718
rect 9588 36654 9640 36660
rect 9404 36644 9456 36650
rect 9404 36586 9456 36592
rect 9416 35290 9444 36586
rect 9600 35630 9628 36654
rect 9588 35624 9640 35630
rect 9588 35566 9640 35572
rect 9404 35284 9456 35290
rect 9404 35226 9456 35232
rect 9496 34740 9548 34746
rect 9600 34728 9628 35566
rect 9772 35488 9824 35494
rect 9772 35430 9824 35436
rect 9784 35154 9812 35430
rect 9876 35154 9904 38490
rect 10152 38486 10180 42094
rect 10508 42016 10560 42022
rect 10508 41958 10560 41964
rect 10520 41614 10548 41958
rect 10888 41750 10916 42502
rect 10876 41744 10928 41750
rect 10876 41686 10928 41692
rect 10600 41676 10652 41682
rect 10600 41618 10652 41624
rect 10784 41676 10836 41682
rect 10784 41618 10836 41624
rect 10508 41608 10560 41614
rect 10508 41550 10560 41556
rect 10520 41414 10548 41550
rect 10428 41386 10548 41414
rect 10232 41064 10284 41070
rect 10232 41006 10284 41012
rect 10140 38480 10192 38486
rect 10140 38422 10192 38428
rect 10244 38418 10272 41006
rect 10324 40928 10376 40934
rect 10324 40870 10376 40876
rect 10336 39982 10364 40870
rect 10324 39976 10376 39982
rect 10324 39918 10376 39924
rect 10324 39500 10376 39506
rect 10324 39442 10376 39448
rect 10336 38554 10364 39442
rect 10324 38548 10376 38554
rect 10324 38490 10376 38496
rect 10232 38412 10284 38418
rect 10232 38354 10284 38360
rect 10230 37768 10286 37777
rect 10230 37703 10286 37712
rect 10244 37670 10272 37703
rect 10048 37664 10100 37670
rect 10048 37606 10100 37612
rect 10232 37664 10284 37670
rect 10232 37606 10284 37612
rect 9954 36816 10010 36825
rect 9954 36751 10010 36760
rect 9772 35148 9824 35154
rect 9772 35090 9824 35096
rect 9864 35148 9916 35154
rect 9864 35090 9916 35096
rect 9548 34700 9628 34728
rect 9496 34682 9548 34688
rect 9588 34536 9640 34542
rect 9588 34478 9640 34484
rect 9600 33998 9628 34478
rect 9588 33992 9640 33998
rect 9588 33934 9640 33940
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9496 32768 9548 32774
rect 9496 32710 9548 32716
rect 9128 32496 9180 32502
rect 9128 32438 9180 32444
rect 9140 32026 9168 32438
rect 9404 32360 9456 32366
rect 9404 32302 9456 32308
rect 9312 32224 9364 32230
rect 9312 32166 9364 32172
rect 9128 32020 9180 32026
rect 9128 31962 9180 31968
rect 9324 31958 9352 32166
rect 9416 32026 9444 32302
rect 9404 32020 9456 32026
rect 9404 31962 9456 31968
rect 9312 31952 9364 31958
rect 9312 31894 9364 31900
rect 9324 31770 9352 31894
rect 9140 31742 9352 31770
rect 9140 31686 9168 31742
rect 9128 31680 9180 31686
rect 9128 31622 9180 31628
rect 9140 29714 9168 31622
rect 9508 29850 9536 32710
rect 9600 31754 9628 33934
rect 9772 33448 9824 33454
rect 9772 33390 9824 33396
rect 9784 32910 9812 33390
rect 9772 32904 9824 32910
rect 9772 32846 9824 32852
rect 9864 32360 9916 32366
rect 9864 32302 9916 32308
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 9588 31748 9640 31754
rect 9588 31690 9640 31696
rect 9600 31346 9628 31690
rect 9692 31414 9720 31962
rect 9770 31920 9826 31929
rect 9770 31855 9772 31864
rect 9824 31855 9826 31864
rect 9772 31826 9824 31832
rect 9876 31482 9904 32302
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 9680 31408 9732 31414
rect 9680 31350 9732 31356
rect 9588 31340 9640 31346
rect 9588 31282 9640 31288
rect 9600 30802 9628 31282
rect 9588 30796 9640 30802
rect 9588 30738 9640 30744
rect 9588 30320 9640 30326
rect 9588 30262 9640 30268
rect 9496 29844 9548 29850
rect 9496 29786 9548 29792
rect 9128 29708 9180 29714
rect 9128 29650 9180 29656
rect 9600 29578 9628 30262
rect 9312 29572 9364 29578
rect 9312 29514 9364 29520
rect 9588 29572 9640 29578
rect 9588 29514 9640 29520
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 9140 26450 9168 26930
rect 9220 26580 9272 26586
rect 9220 26522 9272 26528
rect 9128 26444 9180 26450
rect 9128 26386 9180 26392
rect 9232 26042 9260 26522
rect 8852 26036 8904 26042
rect 8852 25978 8904 25984
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 8760 25832 8812 25838
rect 8760 25774 8812 25780
rect 9324 24750 9352 29514
rect 9968 29458 9996 36751
rect 10060 30394 10088 37606
rect 10428 37466 10456 41386
rect 10508 41132 10560 41138
rect 10508 41074 10560 41080
rect 10520 38010 10548 41074
rect 10612 40730 10640 41618
rect 10796 41562 10824 41618
rect 10704 41534 10824 41562
rect 10704 40934 10732 41534
rect 10784 41472 10836 41478
rect 10784 41414 10836 41420
rect 10692 40928 10744 40934
rect 10692 40870 10744 40876
rect 10600 40724 10652 40730
rect 10600 40666 10652 40672
rect 10796 40202 10824 41414
rect 10704 40174 10824 40202
rect 10704 38570 10732 40174
rect 10888 38978 10916 41686
rect 10980 41478 11008 43590
rect 11072 41818 11100 46514
rect 11152 45824 11204 45830
rect 11152 45766 11204 45772
rect 11164 44538 11192 45766
rect 11256 45082 11284 54062
rect 11624 53242 11652 54130
rect 11612 53236 11664 53242
rect 11612 53178 11664 53184
rect 11808 53038 11836 56200
rect 12176 53650 12204 56200
rect 12348 54188 12400 54194
rect 12348 54130 12400 54136
rect 12164 53644 12216 53650
rect 12164 53586 12216 53592
rect 12072 53576 12124 53582
rect 12072 53518 12124 53524
rect 11888 53100 11940 53106
rect 11888 53042 11940 53048
rect 11796 53032 11848 53038
rect 11796 52974 11848 52980
rect 11900 52154 11928 53042
rect 11888 52148 11940 52154
rect 11888 52090 11940 52096
rect 11980 52012 12032 52018
rect 11980 51954 12032 51960
rect 11992 49434 12020 51954
rect 11980 49428 12032 49434
rect 11980 49370 12032 49376
rect 11336 48000 11388 48006
rect 11336 47942 11388 47948
rect 11244 45076 11296 45082
rect 11244 45018 11296 45024
rect 11152 44532 11204 44538
rect 11152 44474 11204 44480
rect 11348 43994 11376 47942
rect 11428 47660 11480 47666
rect 11428 47602 11480 47608
rect 11336 43988 11388 43994
rect 11336 43930 11388 43936
rect 11440 42362 11468 47602
rect 11888 46504 11940 46510
rect 11888 46446 11940 46452
rect 11900 46034 11928 46446
rect 11888 46028 11940 46034
rect 11888 45970 11940 45976
rect 11796 45960 11848 45966
rect 11796 45902 11848 45908
rect 11704 44328 11756 44334
rect 11610 44296 11666 44305
rect 11704 44270 11756 44276
rect 11610 44231 11612 44240
rect 11664 44231 11666 44240
rect 11612 44202 11664 44208
rect 11716 43178 11744 44270
rect 11704 43172 11756 43178
rect 11704 43114 11756 43120
rect 11428 42356 11480 42362
rect 11428 42298 11480 42304
rect 11152 42220 11204 42226
rect 11152 42162 11204 42168
rect 11060 41812 11112 41818
rect 11060 41754 11112 41760
rect 10968 41472 11020 41478
rect 10968 41414 11020 41420
rect 11060 41472 11112 41478
rect 11060 41414 11112 41420
rect 10968 39976 11020 39982
rect 10968 39918 11020 39924
rect 10980 39098 11008 39918
rect 10968 39092 11020 39098
rect 10968 39034 11020 39040
rect 10888 38950 11008 38978
rect 10980 38894 11008 38950
rect 10968 38888 11020 38894
rect 10968 38830 11020 38836
rect 10704 38542 10916 38570
rect 11072 38554 11100 41414
rect 11164 38826 11192 42162
rect 11808 41414 11836 45902
rect 12084 45082 12112 53518
rect 12360 52154 12388 54130
rect 12544 54126 12572 56200
rect 12912 54262 12940 56200
rect 13280 55214 13308 56200
rect 13280 55186 13400 55214
rect 12900 54256 12952 54262
rect 12900 54198 12952 54204
rect 12532 54120 12584 54126
rect 12532 54062 12584 54068
rect 12716 53984 12768 53990
rect 12716 53926 12768 53932
rect 12624 53576 12676 53582
rect 12624 53518 12676 53524
rect 12636 52698 12664 53518
rect 12624 52692 12676 52698
rect 12624 52634 12676 52640
rect 12348 52148 12400 52154
rect 12348 52090 12400 52096
rect 12532 48748 12584 48754
rect 12532 48690 12584 48696
rect 12164 46912 12216 46918
rect 12164 46854 12216 46860
rect 12176 46034 12204 46854
rect 12164 46028 12216 46034
rect 12164 45970 12216 45976
rect 12256 45348 12308 45354
rect 12256 45290 12308 45296
rect 12072 45076 12124 45082
rect 12072 45018 12124 45024
rect 12268 44266 12296 45290
rect 12440 45280 12492 45286
rect 12440 45222 12492 45228
rect 12452 44810 12480 45222
rect 12544 45082 12572 48690
rect 12624 46980 12676 46986
rect 12624 46922 12676 46928
rect 12636 46034 12664 46922
rect 12624 46028 12676 46034
rect 12624 45970 12676 45976
rect 12636 45898 12664 45970
rect 12624 45892 12676 45898
rect 12624 45834 12676 45840
rect 12532 45076 12584 45082
rect 12532 45018 12584 45024
rect 12624 44940 12676 44946
rect 12624 44882 12676 44888
rect 12440 44804 12492 44810
rect 12440 44746 12492 44752
rect 12348 44464 12400 44470
rect 12348 44406 12400 44412
rect 12256 44260 12308 44266
rect 12256 44202 12308 44208
rect 12072 43648 12124 43654
rect 12072 43590 12124 43596
rect 11716 41386 11836 41414
rect 11716 41274 11744 41386
rect 11520 41268 11572 41274
rect 11520 41210 11572 41216
rect 11704 41268 11756 41274
rect 11704 41210 11756 41216
rect 11242 40488 11298 40497
rect 11242 40423 11298 40432
rect 11152 38820 11204 38826
rect 11152 38762 11204 38768
rect 10692 38208 10744 38214
rect 10692 38150 10744 38156
rect 10784 38208 10836 38214
rect 10784 38150 10836 38156
rect 10508 38004 10560 38010
rect 10508 37946 10560 37952
rect 10508 37868 10560 37874
rect 10508 37810 10560 37816
rect 10520 37777 10548 37810
rect 10506 37768 10562 37777
rect 10506 37703 10562 37712
rect 10416 37460 10468 37466
rect 10416 37402 10468 37408
rect 10428 37194 10456 37402
rect 10704 37194 10732 38150
rect 10796 38010 10824 38150
rect 10784 38004 10836 38010
rect 10784 37946 10836 37952
rect 10888 37466 10916 38542
rect 11060 38548 11112 38554
rect 11060 38490 11112 38496
rect 11060 38208 11112 38214
rect 11060 38150 11112 38156
rect 10876 37460 10928 37466
rect 10876 37402 10928 37408
rect 10888 37330 10916 37402
rect 10876 37324 10928 37330
rect 10876 37266 10928 37272
rect 10416 37188 10468 37194
rect 10416 37130 10468 37136
rect 10692 37188 10744 37194
rect 10692 37130 10744 37136
rect 10428 36854 10456 37130
rect 10784 37120 10836 37126
rect 10784 37062 10836 37068
rect 10416 36848 10468 36854
rect 10416 36790 10468 36796
rect 10416 36100 10468 36106
rect 10416 36042 10468 36048
rect 10232 35828 10284 35834
rect 10232 35770 10284 35776
rect 10244 35494 10272 35770
rect 10232 35488 10284 35494
rect 10232 35430 10284 35436
rect 10140 34400 10192 34406
rect 10140 34342 10192 34348
rect 10152 32978 10180 34342
rect 10428 33658 10456 36042
rect 10796 35494 10824 37062
rect 10968 36712 11020 36718
rect 10968 36654 11020 36660
rect 10876 36576 10928 36582
rect 10876 36518 10928 36524
rect 10784 35488 10836 35494
rect 10784 35430 10836 35436
rect 10692 34944 10744 34950
rect 10692 34886 10744 34892
rect 10704 34746 10732 34886
rect 10692 34740 10744 34746
rect 10692 34682 10744 34688
rect 10796 34406 10824 35430
rect 10784 34400 10836 34406
rect 10784 34342 10836 34348
rect 10888 33658 10916 36518
rect 10980 35630 11008 36654
rect 10968 35624 11020 35630
rect 10968 35566 11020 35572
rect 10980 34542 11008 35566
rect 10968 34536 11020 34542
rect 10968 34478 11020 34484
rect 10968 33856 11020 33862
rect 10968 33798 11020 33804
rect 10416 33652 10468 33658
rect 10416 33594 10468 33600
rect 10876 33652 10928 33658
rect 10876 33594 10928 33600
rect 10980 33590 11008 33798
rect 10968 33584 11020 33590
rect 10968 33526 11020 33532
rect 10600 33312 10652 33318
rect 10600 33254 10652 33260
rect 10612 33114 10640 33254
rect 11072 33114 11100 38150
rect 11256 37942 11284 40423
rect 11532 40186 11560 41210
rect 11888 40520 11940 40526
rect 11980 40520 12032 40526
rect 11888 40462 11940 40468
rect 11978 40488 11980 40497
rect 12032 40488 12034 40497
rect 11520 40180 11572 40186
rect 11520 40122 11572 40128
rect 11532 39370 11560 40122
rect 11520 39364 11572 39370
rect 11520 39306 11572 39312
rect 11520 39024 11572 39030
rect 11520 38966 11572 38972
rect 11532 38758 11560 38966
rect 11520 38752 11572 38758
rect 11520 38694 11572 38700
rect 11704 38752 11756 38758
rect 11704 38694 11756 38700
rect 11244 37936 11296 37942
rect 11244 37878 11296 37884
rect 11532 37398 11560 38694
rect 11610 38312 11666 38321
rect 11610 38247 11666 38256
rect 11520 37392 11572 37398
rect 11520 37334 11572 37340
rect 11624 37210 11652 38247
rect 11532 37182 11652 37210
rect 11716 37194 11744 38694
rect 11704 37188 11756 37194
rect 11244 37120 11296 37126
rect 11244 37062 11296 37068
rect 11152 35148 11204 35154
rect 11152 35090 11204 35096
rect 11164 34474 11192 35090
rect 11152 34468 11204 34474
rect 11152 34410 11204 34416
rect 11152 34196 11204 34202
rect 11152 34138 11204 34144
rect 10600 33108 10652 33114
rect 10600 33050 10652 33056
rect 11060 33108 11112 33114
rect 11060 33050 11112 33056
rect 10140 32972 10192 32978
rect 10140 32914 10192 32920
rect 10152 32026 10180 32914
rect 10612 32910 10640 33050
rect 10600 32904 10652 32910
rect 10600 32846 10652 32852
rect 10968 32224 11020 32230
rect 10968 32166 11020 32172
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 10980 31754 11008 32166
rect 10968 31748 11020 31754
rect 10968 31690 11020 31696
rect 10876 30796 10928 30802
rect 11164 30784 11192 34138
rect 10928 30756 11192 30784
rect 10876 30738 10928 30744
rect 10048 30388 10100 30394
rect 10048 30330 10100 30336
rect 10324 30388 10376 30394
rect 10324 30330 10376 30336
rect 10048 29504 10100 29510
rect 9968 29452 10048 29458
rect 9968 29446 10100 29452
rect 9968 29430 10088 29446
rect 9496 29232 9548 29238
rect 9496 29174 9548 29180
rect 9404 29096 9456 29102
rect 9404 29038 9456 29044
rect 9416 28626 9444 29038
rect 9508 28762 9536 29174
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 9496 28756 9548 28762
rect 9496 28698 9548 28704
rect 9404 28620 9456 28626
rect 9404 28562 9456 28568
rect 9416 26926 9444 28562
rect 9692 27946 9720 28902
rect 9864 28688 9916 28694
rect 9864 28630 9916 28636
rect 9680 27940 9732 27946
rect 9680 27882 9732 27888
rect 9876 27674 9904 28630
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 9968 27878 9996 28494
rect 9956 27872 10008 27878
rect 9956 27814 10008 27820
rect 9864 27668 9916 27674
rect 9864 27610 9916 27616
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9680 26852 9732 26858
rect 9680 26794 9732 26800
rect 9588 26308 9640 26314
rect 9588 26250 9640 26256
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9416 25362 9444 25842
rect 9600 25770 9628 26250
rect 9588 25764 9640 25770
rect 9588 25706 9640 25712
rect 9692 25362 9720 26794
rect 9772 25968 9824 25974
rect 9772 25910 9824 25916
rect 9404 25356 9456 25362
rect 9404 25298 9456 25304
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 9784 25226 9812 25910
rect 9876 25838 9904 27610
rect 9968 27470 9996 27814
rect 9956 27464 10008 27470
rect 9956 27406 10008 27412
rect 9968 26382 9996 27406
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9864 25832 9916 25838
rect 9864 25774 9916 25780
rect 9772 25220 9824 25226
rect 9772 25162 9824 25168
rect 9496 24948 9548 24954
rect 9496 24890 9548 24896
rect 9312 24744 9364 24750
rect 9312 24686 9364 24692
rect 9324 24410 9352 24686
rect 8760 24404 8812 24410
rect 8760 24346 8812 24352
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 8772 21894 8800 24346
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 9324 23798 9352 24006
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9416 22778 9444 24006
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8680 19718 8708 20402
rect 8772 20330 8800 21422
rect 8864 20602 8892 22510
rect 9404 22500 9456 22506
rect 9404 22442 9456 22448
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8956 20602 8984 21490
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8864 19922 8892 20538
rect 9048 20534 9076 21422
rect 9036 20528 9088 20534
rect 9036 20470 9088 20476
rect 9048 20262 9076 20470
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8956 19718 8984 19790
rect 8668 19712 8720 19718
rect 8666 19680 8668 19689
rect 8944 19712 8996 19718
rect 8720 19680 8722 19689
rect 8944 19654 8996 19660
rect 8666 19615 8722 19624
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7852 18222 7880 19110
rect 8680 18630 8708 19314
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 8496 18154 8524 18566
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7208 16522 7236 16730
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 7208 16182 7236 16458
rect 7300 16250 7328 17478
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7196 16176 7248 16182
rect 7196 16118 7248 16124
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7116 9518 7144 13194
rect 7760 12986 7788 18022
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 8128 16794 8156 17206
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8404 16726 8432 17682
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8312 16046 8340 16526
rect 8404 16046 8432 16662
rect 8496 16658 8524 18090
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8588 16794 8616 17478
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8496 16454 8524 16594
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8496 15366 8524 16390
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8496 13394 8524 15302
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 8404 12918 8432 13262
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 8680 5710 8708 18566
rect 8772 17678 8800 19110
rect 8956 18970 8984 19654
rect 9324 19446 9352 20334
rect 9416 19514 9444 22442
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8772 17202 8800 17478
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8864 17134 8892 17274
rect 8956 17270 8984 18906
rect 8944 17264 8996 17270
rect 8944 17206 8996 17212
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8760 16720 8812 16726
rect 8760 16662 8812 16668
rect 8772 15706 8800 16662
rect 9048 16590 9076 19246
rect 9312 18624 9364 18630
rect 9232 18572 9312 18578
rect 9232 18566 9364 18572
rect 9232 18550 9352 18566
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8772 15162 8800 15642
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8772 12782 8800 13126
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 9232 7818 9260 18550
rect 9508 17864 9536 24890
rect 9680 24744 9732 24750
rect 9680 24686 9732 24692
rect 9692 23866 9720 24686
rect 9864 24268 9916 24274
rect 9864 24210 9916 24216
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 9784 23866 9812 24006
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9876 23730 9904 24210
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9968 23526 9996 26318
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 9772 23248 9824 23254
rect 9772 23190 9824 23196
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9600 19718 9628 20742
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 9600 18630 9628 19246
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9692 18426 9720 22578
rect 9784 21690 9812 23190
rect 9968 22982 9996 23462
rect 10060 23186 10088 29430
rect 10232 27328 10284 27334
rect 10232 27270 10284 27276
rect 10140 26852 10192 26858
rect 10140 26794 10192 26800
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 9956 22976 10008 22982
rect 9956 22918 10008 22924
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9968 20874 9996 22918
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9324 17836 9536 17864
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9324 5914 9352 17836
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9416 15094 9444 17682
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9508 17338 9536 17478
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 16561 9536 16934
rect 9600 16590 9628 17614
rect 9692 17610 9720 18362
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 9968 16726 9996 17002
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9588 16584 9640 16590
rect 9494 16552 9550 16561
rect 9588 16526 9640 16532
rect 9494 16487 9550 16496
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 15706 9996 16390
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9404 15088 9456 15094
rect 9404 15030 9456 15036
rect 9416 14056 9444 15030
rect 9416 14028 9536 14056
rect 9508 13870 9536 14028
rect 9600 14006 9628 15098
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9968 14482 9996 14758
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9588 14000 9640 14006
rect 9588 13942 9640 13948
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9600 13462 9628 13942
rect 9876 13734 9904 14214
rect 9968 14074 9996 14418
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9864 13388 9916 13394
rect 9968 13376 9996 14010
rect 9916 13348 9996 13376
rect 9864 13330 9916 13336
rect 9968 12918 9996 13348
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 9692 12306 9720 12854
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 8668 5704 8720 5710
rect 8482 5672 8538 5681
rect 8668 5646 8720 5652
rect 8482 5607 8538 5616
rect 9312 5636 9364 5642
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7208 4146 7236 4558
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6840 3534 6868 3878
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6472 2746 6592 2774
rect 6472 800 6500 2746
rect 6840 800 6868 3470
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7116 2310 7144 2518
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7208 800 7236 2994
rect 7392 2446 7420 4966
rect 8496 4826 8524 5607
rect 9312 5578 9364 5584
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7484 2650 7512 2790
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7668 2582 7696 4490
rect 7852 3534 7880 4490
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7300 2106 7328 2314
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7576 800 7604 2382
rect 7852 1986 7880 3470
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8312 3194 8340 4558
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8496 3058 8524 4422
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8588 3738 8616 4082
rect 8864 4010 8892 5510
rect 9036 4548 9088 4554
rect 9036 4490 9088 4496
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 9048 3058 9076 4490
rect 9324 3738 9352 5578
rect 9586 5128 9642 5137
rect 9586 5063 9642 5072
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8496 2774 8524 2994
rect 8496 2746 8708 2774
rect 8220 2378 8340 2394
rect 8208 2372 8340 2378
rect 8260 2366 8340 2372
rect 8208 2314 8260 2320
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 7852 1958 7972 1986
rect 7944 800 7972 1958
rect 8312 800 8340 2366
rect 8680 800 8708 2746
rect 9048 800 9076 2994
rect 9416 800 9444 4082
rect 9600 3058 9628 5063
rect 10060 4758 10088 22714
rect 10152 17626 10180 26794
rect 10244 26450 10272 27270
rect 10232 26444 10284 26450
rect 10232 26386 10284 26392
rect 10336 26330 10364 30330
rect 11164 30190 11192 30756
rect 11152 30184 11204 30190
rect 11152 30126 11204 30132
rect 10416 30048 10468 30054
rect 10416 29990 10468 29996
rect 10428 29646 10456 29990
rect 10416 29640 10468 29646
rect 10416 29582 10468 29588
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10600 27940 10652 27946
rect 10600 27882 10652 27888
rect 10612 26790 10640 27882
rect 10692 27872 10744 27878
rect 10692 27814 10744 27820
rect 10704 27130 10732 27814
rect 10692 27124 10744 27130
rect 10692 27066 10744 27072
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10244 26302 10364 26330
rect 10244 21894 10272 26302
rect 10520 26042 10548 26726
rect 10704 26314 10732 27066
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 10508 26036 10560 26042
rect 10508 25978 10560 25984
rect 10704 25974 10732 26250
rect 10692 25968 10744 25974
rect 10692 25910 10744 25916
rect 10796 25294 10824 29446
rect 10876 29028 10928 29034
rect 10876 28970 10928 28976
rect 10888 26042 10916 28970
rect 11256 27062 11284 37062
rect 11336 36032 11388 36038
rect 11336 35974 11388 35980
rect 11348 33658 11376 35974
rect 11336 33652 11388 33658
rect 11336 33594 11388 33600
rect 11336 31408 11388 31414
rect 11336 31350 11388 31356
rect 11348 30802 11376 31350
rect 11336 30796 11388 30802
rect 11336 30738 11388 30744
rect 11428 30728 11480 30734
rect 11426 30696 11428 30705
rect 11480 30696 11482 30705
rect 11426 30631 11482 30640
rect 11336 30592 11388 30598
rect 11336 30534 11388 30540
rect 11348 29782 11376 30534
rect 11336 29776 11388 29782
rect 11336 29718 11388 29724
rect 11348 28626 11376 29718
rect 11336 28620 11388 28626
rect 11336 28562 11388 28568
rect 11428 27396 11480 27402
rect 11428 27338 11480 27344
rect 11244 27056 11296 27062
rect 11244 26998 11296 27004
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 11440 25362 11468 27338
rect 11428 25356 11480 25362
rect 11428 25298 11480 25304
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 11152 25152 11204 25158
rect 11152 25094 11204 25100
rect 11164 24954 11192 25094
rect 11152 24948 11204 24954
rect 11152 24890 11204 24896
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 10324 24404 10376 24410
rect 10324 24346 10376 24352
rect 10232 21888 10284 21894
rect 10232 21830 10284 21836
rect 10244 18306 10272 21830
rect 10336 20874 10364 24346
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 10428 21010 10456 24210
rect 10784 24064 10836 24070
rect 11072 24041 11100 24210
rect 11164 24206 11192 24550
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 11532 24138 11560 37182
rect 11704 37130 11756 37136
rect 11900 36718 11928 40462
rect 11978 40423 12034 40432
rect 11980 38820 12032 38826
rect 11980 38762 12032 38768
rect 11992 38282 12020 38762
rect 11980 38276 12032 38282
rect 11980 38218 12032 38224
rect 12084 37890 12112 43590
rect 12164 42900 12216 42906
rect 12164 42842 12216 42848
rect 12176 42702 12204 42842
rect 12164 42696 12216 42702
rect 12164 42638 12216 42644
rect 12268 41070 12296 44202
rect 12360 43314 12388 44406
rect 12348 43308 12400 43314
rect 12348 43250 12400 43256
rect 12360 42770 12388 43250
rect 12348 42764 12400 42770
rect 12348 42706 12400 42712
rect 12360 41682 12388 42706
rect 12452 42702 12480 44746
rect 12532 44736 12584 44742
rect 12532 44678 12584 44684
rect 12440 42696 12492 42702
rect 12440 42638 12492 42644
rect 12440 42560 12492 42566
rect 12440 42502 12492 42508
rect 12452 42158 12480 42502
rect 12440 42152 12492 42158
rect 12440 42094 12492 42100
rect 12348 41676 12400 41682
rect 12348 41618 12400 41624
rect 12348 41472 12400 41478
rect 12348 41414 12400 41420
rect 12256 41064 12308 41070
rect 12256 41006 12308 41012
rect 12256 40452 12308 40458
rect 12256 40394 12308 40400
rect 12164 40384 12216 40390
rect 12164 40326 12216 40332
rect 12176 38418 12204 40326
rect 12268 40186 12296 40394
rect 12256 40180 12308 40186
rect 12256 40122 12308 40128
rect 12256 39636 12308 39642
rect 12256 39578 12308 39584
rect 12164 38412 12216 38418
rect 12164 38354 12216 38360
rect 12084 37862 12204 37890
rect 12072 37664 12124 37670
rect 12072 37606 12124 37612
rect 12084 37369 12112 37606
rect 12070 37360 12126 37369
rect 12070 37295 12126 37304
rect 12072 36780 12124 36786
rect 12072 36722 12124 36728
rect 11888 36712 11940 36718
rect 11888 36654 11940 36660
rect 11980 35624 12032 35630
rect 11980 35566 12032 35572
rect 11704 35488 11756 35494
rect 11704 35430 11756 35436
rect 11716 34066 11744 35430
rect 11992 35222 12020 35566
rect 11980 35216 12032 35222
rect 11980 35158 12032 35164
rect 12084 34678 12112 36722
rect 12072 34672 12124 34678
rect 12072 34614 12124 34620
rect 11796 34400 11848 34406
rect 11796 34342 11848 34348
rect 11704 34060 11756 34066
rect 11704 34002 11756 34008
rect 11808 33998 11836 34342
rect 11796 33992 11848 33998
rect 11796 33934 11848 33940
rect 11888 33516 11940 33522
rect 11888 33458 11940 33464
rect 11610 33008 11666 33017
rect 11610 32943 11612 32952
rect 11664 32943 11666 32952
rect 11612 32914 11664 32920
rect 11624 32774 11652 32914
rect 11612 32768 11664 32774
rect 11612 32710 11664 32716
rect 11900 32026 11928 33458
rect 11980 32904 12032 32910
rect 11980 32846 12032 32852
rect 11888 32020 11940 32026
rect 11888 31962 11940 31968
rect 11704 31680 11756 31686
rect 11704 31622 11756 31628
rect 11716 30870 11744 31622
rect 11704 30864 11756 30870
rect 11704 30806 11756 30812
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11900 29510 11928 29990
rect 11888 29504 11940 29510
rect 11888 29446 11940 29452
rect 11796 25832 11848 25838
rect 11796 25774 11848 25780
rect 11808 25294 11836 25774
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11520 24132 11572 24138
rect 11520 24074 11572 24080
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 10784 24006 10836 24012
rect 11058 24032 11114 24041
rect 10796 23866 10824 24006
rect 11058 23967 11114 23976
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 11808 23798 11836 24074
rect 11900 24041 11928 29446
rect 11992 25158 12020 32846
rect 12084 32298 12112 34614
rect 12072 32292 12124 32298
rect 12072 32234 12124 32240
rect 12176 31958 12204 37862
rect 12268 33114 12296 39578
rect 12360 38554 12388 41414
rect 12440 40044 12492 40050
rect 12440 39986 12492 39992
rect 12452 39506 12480 39986
rect 12440 39500 12492 39506
rect 12440 39442 12492 39448
rect 12452 39030 12480 39442
rect 12440 39024 12492 39030
rect 12440 38966 12492 38972
rect 12348 38548 12400 38554
rect 12348 38490 12400 38496
rect 12440 38004 12492 38010
rect 12440 37946 12492 37952
rect 12348 37664 12400 37670
rect 12348 37606 12400 37612
rect 12360 36174 12388 37606
rect 12348 36168 12400 36174
rect 12348 36110 12400 36116
rect 12452 35873 12480 37946
rect 12544 37913 12572 44678
rect 12636 43382 12664 44882
rect 12624 43376 12676 43382
rect 12624 43318 12676 43324
rect 12728 40526 12756 53926
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 13372 53174 13400 55186
rect 13648 54262 13676 56200
rect 14016 54330 14044 56200
rect 14384 56114 14412 56200
rect 14476 56114 14504 56222
rect 14384 56086 14504 56114
rect 14004 54324 14056 54330
rect 14004 54266 14056 54272
rect 13636 54256 13688 54262
rect 13636 54198 13688 54204
rect 13360 53168 13412 53174
rect 13360 53110 13412 53116
rect 13648 53106 13676 54198
rect 14016 53582 14044 54266
rect 14004 53576 14056 53582
rect 14004 53518 14056 53524
rect 14280 53440 14332 53446
rect 14280 53382 14332 53388
rect 13636 53100 13688 53106
rect 13636 53042 13688 53048
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 14292 52494 14320 53382
rect 14372 52896 14424 52902
rect 14372 52838 14424 52844
rect 14556 52896 14608 52902
rect 14556 52838 14608 52844
rect 12808 52488 12860 52494
rect 12808 52430 12860 52436
rect 13544 52488 13596 52494
rect 13544 52430 13596 52436
rect 14280 52488 14332 52494
rect 14280 52430 14332 52436
rect 12820 48890 12848 52430
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12808 48884 12860 48890
rect 12808 48826 12860 48832
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 13084 46980 13136 46986
rect 13084 46922 13136 46928
rect 13096 46646 13124 46922
rect 13084 46640 13136 46646
rect 13084 46582 13136 46588
rect 13360 46504 13412 46510
rect 13360 46446 13412 46452
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 13372 44470 13400 46446
rect 13452 44872 13504 44878
rect 13452 44814 13504 44820
rect 13360 44464 13412 44470
rect 13360 44406 13412 44412
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 13464 42362 13492 44814
rect 13452 42356 13504 42362
rect 13452 42298 13504 42304
rect 13360 42084 13412 42090
rect 13360 42026 13412 42032
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 12808 41676 12860 41682
rect 12808 41618 12860 41624
rect 12716 40520 12768 40526
rect 12716 40462 12768 40468
rect 12624 40384 12676 40390
rect 12624 40326 12676 40332
rect 12530 37904 12586 37913
rect 12530 37839 12586 37848
rect 12544 36378 12572 37839
rect 12532 36372 12584 36378
rect 12532 36314 12584 36320
rect 12438 35864 12494 35873
rect 12438 35799 12494 35808
rect 12348 33856 12400 33862
rect 12348 33798 12400 33804
rect 12256 33108 12308 33114
rect 12256 33050 12308 33056
rect 12256 32360 12308 32366
rect 12254 32328 12256 32337
rect 12308 32328 12310 32337
rect 12254 32263 12310 32272
rect 12360 32230 12388 33798
rect 12452 33114 12480 35799
rect 12544 33862 12572 36314
rect 12636 34066 12664 40326
rect 12820 40050 12848 41618
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12808 40044 12860 40050
rect 12808 39986 12860 39992
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 13084 39636 13136 39642
rect 13084 39578 13136 39584
rect 13096 39030 13124 39578
rect 13084 39024 13136 39030
rect 13084 38966 13136 38972
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 13266 38448 13322 38457
rect 13266 38383 13268 38392
rect 13320 38383 13322 38392
rect 13268 38354 13320 38360
rect 12716 38344 12768 38350
rect 12716 38286 12768 38292
rect 12728 37874 12756 38286
rect 12716 37868 12768 37874
rect 12716 37810 12768 37816
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 13084 37188 13136 37194
rect 13084 37130 13136 37136
rect 12716 37120 12768 37126
rect 12716 37062 12768 37068
rect 12728 36922 12756 37062
rect 12716 36916 12768 36922
rect 12716 36858 12768 36864
rect 13096 36854 13124 37130
rect 13084 36848 13136 36854
rect 13084 36790 13136 36796
rect 12808 36712 12860 36718
rect 12808 36654 12860 36660
rect 12716 36236 12768 36242
rect 12716 36178 12768 36184
rect 12728 36038 12756 36178
rect 12716 36032 12768 36038
rect 12716 35974 12768 35980
rect 12624 34060 12676 34066
rect 12624 34002 12676 34008
rect 12532 33856 12584 33862
rect 12532 33798 12584 33804
rect 12624 33584 12676 33590
rect 12624 33526 12676 33532
rect 12532 33516 12584 33522
rect 12532 33458 12584 33464
rect 12544 33318 12572 33458
rect 12532 33312 12584 33318
rect 12530 33280 12532 33289
rect 12584 33280 12586 33289
rect 12530 33215 12586 33224
rect 12440 33108 12492 33114
rect 12440 33050 12492 33056
rect 12532 32904 12584 32910
rect 12532 32846 12584 32852
rect 12348 32224 12400 32230
rect 12348 32166 12400 32172
rect 12164 31952 12216 31958
rect 12164 31894 12216 31900
rect 12440 31680 12492 31686
rect 12440 31622 12492 31628
rect 12452 30190 12480 31622
rect 12440 30184 12492 30190
rect 12440 30126 12492 30132
rect 12348 30048 12400 30054
rect 12348 29990 12400 29996
rect 12360 29578 12388 29990
rect 12348 29572 12400 29578
rect 12348 29514 12400 29520
rect 12544 28994 12572 32846
rect 12636 30938 12664 33526
rect 12728 31686 12756 35974
rect 12820 34746 12848 36654
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 13372 36378 13400 42026
rect 13452 39500 13504 39506
rect 13452 39442 13504 39448
rect 13464 38486 13492 39442
rect 13452 38480 13504 38486
rect 13452 38422 13504 38428
rect 13556 38010 13584 52430
rect 14384 52086 14412 52838
rect 14568 52426 14596 52838
rect 14556 52420 14608 52426
rect 14556 52362 14608 52368
rect 14464 52352 14516 52358
rect 14464 52294 14516 52300
rect 14372 52080 14424 52086
rect 14372 52022 14424 52028
rect 14096 51876 14148 51882
rect 14096 51818 14148 51824
rect 13728 46368 13780 46374
rect 13728 46310 13780 46316
rect 13636 45824 13688 45830
rect 13636 45766 13688 45772
rect 13648 44198 13676 45766
rect 13740 44946 13768 46310
rect 14004 46028 14056 46034
rect 14004 45970 14056 45976
rect 14016 45558 14044 45970
rect 14004 45552 14056 45558
rect 14004 45494 14056 45500
rect 13728 44940 13780 44946
rect 13728 44882 13780 44888
rect 14016 44470 14044 45494
rect 14004 44464 14056 44470
rect 14004 44406 14056 44412
rect 13636 44192 13688 44198
rect 13636 44134 13688 44140
rect 14016 43382 14044 44406
rect 14004 43376 14056 43382
rect 13924 43336 14004 43364
rect 13924 42906 13952 43336
rect 14004 43318 14056 43324
rect 14004 43104 14056 43110
rect 14004 43046 14056 43052
rect 13912 42900 13964 42906
rect 13912 42842 13964 42848
rect 13636 41676 13688 41682
rect 13636 41618 13688 41624
rect 13912 41676 13964 41682
rect 13912 41618 13964 41624
rect 13648 41138 13676 41618
rect 13636 41132 13688 41138
rect 13636 41074 13688 41080
rect 13924 41070 13952 41618
rect 13912 41064 13964 41070
rect 13912 41006 13964 41012
rect 13636 40588 13688 40594
rect 13636 40530 13688 40536
rect 13820 40588 13872 40594
rect 13820 40530 13872 40536
rect 13544 38004 13596 38010
rect 13544 37946 13596 37952
rect 13452 37800 13504 37806
rect 13452 37742 13504 37748
rect 13544 37800 13596 37806
rect 13544 37742 13596 37748
rect 13360 36372 13412 36378
rect 13360 36314 13412 36320
rect 13464 35834 13492 37742
rect 13556 37262 13584 37742
rect 13544 37256 13596 37262
rect 13544 37198 13596 37204
rect 13544 36916 13596 36922
rect 13544 36858 13596 36864
rect 13556 36378 13584 36858
rect 13544 36372 13596 36378
rect 13544 36314 13596 36320
rect 13544 36236 13596 36242
rect 13544 36178 13596 36184
rect 13556 35834 13584 36178
rect 13452 35828 13504 35834
rect 13452 35770 13504 35776
rect 13544 35828 13596 35834
rect 13544 35770 13596 35776
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 13360 34944 13412 34950
rect 13360 34886 13412 34892
rect 12808 34740 12860 34746
rect 12808 34682 12860 34688
rect 13372 34610 13400 34886
rect 13360 34604 13412 34610
rect 13360 34546 13412 34552
rect 13360 34468 13412 34474
rect 13360 34410 13412 34416
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12808 33856 12860 33862
rect 12808 33798 12860 33804
rect 13176 33856 13228 33862
rect 13176 33798 13228 33804
rect 12716 31680 12768 31686
rect 12716 31622 12768 31628
rect 12716 31476 12768 31482
rect 12716 31418 12768 31424
rect 12624 30932 12676 30938
rect 12624 30874 12676 30880
rect 12624 30184 12676 30190
rect 12624 30126 12676 30132
rect 12360 28966 12572 28994
rect 12360 28506 12388 28966
rect 12360 28478 12480 28506
rect 12072 27532 12124 27538
rect 12072 27474 12124 27480
rect 12084 27062 12112 27474
rect 12072 27056 12124 27062
rect 12072 26998 12124 27004
rect 12348 26784 12400 26790
rect 12348 26726 12400 26732
rect 12360 26518 12388 26726
rect 12256 26512 12308 26518
rect 12256 26454 12308 26460
rect 12348 26512 12400 26518
rect 12348 26454 12400 26460
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 12072 24608 12124 24614
rect 12072 24550 12124 24556
rect 11980 24064 12032 24070
rect 11886 24032 11942 24041
rect 11980 24006 12032 24012
rect 11886 23967 11942 23976
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 11888 23792 11940 23798
rect 11888 23734 11940 23740
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10784 23180 10836 23186
rect 10784 23122 10836 23128
rect 10796 23050 10824 23122
rect 10980 23118 11008 23462
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 10968 23112 11020 23118
rect 10968 23054 11020 23060
rect 10784 23044 10836 23050
rect 10784 22986 10836 22992
rect 10796 22438 10824 22986
rect 11520 22704 11572 22710
rect 11520 22646 11572 22652
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 11164 22030 11192 22510
rect 11532 22438 11560 22646
rect 11520 22432 11572 22438
rect 11520 22374 11572 22380
rect 11532 22166 11560 22374
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 11060 21412 11112 21418
rect 11060 21354 11112 21360
rect 10508 21140 10560 21146
rect 10508 21082 10560 21088
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10520 20874 10548 21082
rect 10324 20868 10376 20874
rect 10324 20810 10376 20816
rect 10508 20868 10560 20874
rect 10508 20810 10560 20816
rect 10336 19242 10364 20810
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10600 20392 10652 20398
rect 10600 20334 10652 20340
rect 10324 19236 10376 19242
rect 10324 19178 10376 19184
rect 10612 18970 10640 20334
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10704 18306 10732 20742
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10796 18970 10824 19110
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10244 18278 10364 18306
rect 10152 17598 10272 17626
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10152 16794 10180 17478
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10244 16522 10272 17598
rect 10336 16590 10364 18278
rect 10612 18278 10732 18306
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10520 17338 10548 17546
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 10520 16250 10548 17070
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10152 14226 10180 15642
rect 10244 14346 10272 15982
rect 10336 15366 10364 16050
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 10152 14198 10272 14226
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9784 800 9812 3470
rect 9876 2650 9904 4558
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3534 10088 3878
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10152 2990 10180 14010
rect 10244 10742 10272 14198
rect 10336 14074 10364 15302
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10336 5574 10364 13874
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 10244 2446 10272 4422
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10336 3058 10364 3946
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10232 2440 10284 2446
rect 10152 2400 10232 2428
rect 10152 800 10180 2400
rect 10232 2382 10284 2388
rect 10428 2310 10456 14554
rect 10612 13938 10640 18278
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10704 18086 10732 18158
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10704 14618 10732 18022
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10796 5778 10824 18906
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10888 16590 10916 18566
rect 10980 18222 11008 19178
rect 11072 18426 11100 21354
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11164 18766 11192 19110
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10980 17218 11008 18158
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 10980 17190 11100 17218
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10980 16658 11008 17070
rect 11072 17066 11100 17190
rect 11348 17134 11376 17546
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10888 14958 10916 15302
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10888 12442 10916 14894
rect 10980 14278 11008 16594
rect 11348 15570 11376 17070
rect 11440 16250 11468 21830
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11532 16250 11560 20470
rect 11624 20330 11652 23122
rect 11716 23118 11744 23598
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11900 22710 11928 23734
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11900 20942 11928 21966
rect 11992 21690 12020 24006
rect 12084 22778 12112 24550
rect 12164 23724 12216 23730
rect 12164 23666 12216 23672
rect 12176 23526 12204 23666
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 12176 23118 12204 23462
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 12164 22092 12216 22098
rect 12164 22034 12216 22040
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11612 20324 11664 20330
rect 11612 20266 11664 20272
rect 11624 19854 11652 20266
rect 11716 20058 11744 20402
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11624 18630 11652 19790
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11624 18086 11652 18566
rect 11900 18170 11928 20878
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11992 18290 12020 18566
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11900 18142 12020 18170
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 11440 15570 11468 15982
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11348 14550 11376 15506
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 11624 13530 11652 16934
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11716 15706 11744 16390
rect 11808 16182 11836 16390
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11532 12918 11560 13194
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10980 11762 11008 12242
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 11624 6458 11652 13466
rect 11808 12986 11836 13738
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11808 12306 11836 12922
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11256 3942 11284 4082
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 10888 3602 10916 3878
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 10520 800 10548 2994
rect 10888 800 10916 3538
rect 11256 800 11284 3878
rect 11624 800 11652 4558
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11716 3058 11744 3878
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11900 2774 11928 17818
rect 11992 17746 12020 18142
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 11992 15366 12020 17682
rect 12084 17270 12112 20198
rect 12176 19990 12204 22034
rect 12268 21622 12296 26454
rect 12348 25696 12400 25702
rect 12348 25638 12400 25644
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12268 21078 12296 21422
rect 12360 21078 12388 25638
rect 12452 24818 12480 28478
rect 12532 28484 12584 28490
rect 12532 28426 12584 28432
rect 12544 27674 12572 28426
rect 12532 27668 12584 27674
rect 12532 27610 12584 27616
rect 12544 27470 12572 27610
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12544 26858 12572 27406
rect 12532 26852 12584 26858
rect 12532 26794 12584 26800
rect 12544 26586 12572 26794
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12636 25294 12664 30126
rect 12624 25288 12676 25294
rect 12544 25236 12624 25242
rect 12544 25230 12676 25236
rect 12544 25214 12664 25230
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12452 23526 12480 24754
rect 12544 24750 12572 25214
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12636 24954 12664 25094
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12624 24812 12676 24818
rect 12624 24754 12676 24760
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12440 23248 12492 23254
rect 12440 23190 12492 23196
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 12348 21072 12400 21078
rect 12348 21014 12400 21020
rect 12164 19984 12216 19990
rect 12164 19926 12216 19932
rect 12162 19408 12218 19417
rect 12162 19343 12164 19352
rect 12216 19343 12218 19352
rect 12164 19314 12216 19320
rect 12176 18970 12204 19314
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12268 18222 12296 21014
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 12360 19310 12388 20878
rect 12452 19854 12480 23190
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 18358 12480 19110
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 12072 15972 12124 15978
rect 12072 15914 12124 15920
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11992 13530 12020 14350
rect 12084 13530 12112 15914
rect 12176 15162 12204 18158
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 12268 16046 12296 18022
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12268 15094 12296 15302
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12268 14550 12296 15030
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11992 13258 12020 13466
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 12360 4826 12388 18090
rect 12452 17066 12480 18158
rect 12544 18154 12572 24346
rect 12636 23662 12664 24754
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12636 23322 12664 23598
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12624 23180 12676 23186
rect 12624 23122 12676 23128
rect 12636 22982 12664 23122
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12636 20942 12664 22918
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12728 20482 12756 31418
rect 12820 29578 12848 33798
rect 13188 33318 13216 33798
rect 13372 33658 13400 34410
rect 13360 33652 13412 33658
rect 13360 33594 13412 33600
rect 13464 33454 13492 35770
rect 13648 35494 13676 40530
rect 13728 39840 13780 39846
rect 13728 39782 13780 39788
rect 13740 39098 13768 39782
rect 13832 39574 13860 40530
rect 13820 39568 13872 39574
rect 13820 39510 13872 39516
rect 13820 39296 13872 39302
rect 13820 39238 13872 39244
rect 13728 39092 13780 39098
rect 13728 39034 13780 39040
rect 13832 38321 13860 39238
rect 13818 38312 13874 38321
rect 13818 38247 13874 38256
rect 13728 38004 13780 38010
rect 13728 37946 13780 37952
rect 13636 35488 13688 35494
rect 13636 35430 13688 35436
rect 13740 35306 13768 37946
rect 13820 37392 13872 37398
rect 13820 37334 13872 37340
rect 13832 36768 13860 37334
rect 13924 37330 13952 41006
rect 14016 40594 14044 43046
rect 14004 40588 14056 40594
rect 14004 40530 14056 40536
rect 14004 38752 14056 38758
rect 14004 38694 14056 38700
rect 13912 37324 13964 37330
rect 13912 37266 13964 37272
rect 13912 36780 13964 36786
rect 13832 36740 13912 36768
rect 13912 36722 13964 36728
rect 13924 36530 13952 36722
rect 14016 36718 14044 38694
rect 14004 36712 14056 36718
rect 14004 36654 14056 36660
rect 13924 36502 14044 36530
rect 13820 36304 13872 36310
rect 13818 36272 13820 36281
rect 13872 36272 13874 36281
rect 13818 36207 13874 36216
rect 13912 35488 13964 35494
rect 13912 35430 13964 35436
rect 13648 35278 13768 35306
rect 13452 33448 13504 33454
rect 13452 33390 13504 33396
rect 13176 33312 13228 33318
rect 13176 33254 13228 33260
rect 13452 33312 13504 33318
rect 13452 33254 13504 33260
rect 13544 33312 13596 33318
rect 13544 33254 13596 33260
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 13464 32892 13492 33254
rect 13372 32864 13492 32892
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 13372 31482 13400 32864
rect 13452 32224 13504 32230
rect 13452 32166 13504 32172
rect 13360 31476 13412 31482
rect 13360 31418 13412 31424
rect 13268 31272 13320 31278
rect 13320 31232 13400 31260
rect 13268 31214 13320 31220
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 12808 29572 12860 29578
rect 12808 29514 12860 29520
rect 12900 29504 12952 29510
rect 12900 29446 12952 29452
rect 12912 29306 12940 29446
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 13372 28626 13400 31232
rect 13360 28620 13412 28626
rect 13360 28562 13412 28568
rect 13360 28484 13412 28490
rect 13360 28426 13412 28432
rect 12808 28416 12860 28422
rect 12808 28358 12860 28364
rect 13176 28416 13228 28422
rect 13176 28358 13228 28364
rect 13268 28416 13320 28422
rect 13268 28358 13320 28364
rect 12820 27538 12848 28358
rect 13188 28218 13216 28358
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 13280 28082 13308 28358
rect 13372 28218 13400 28426
rect 13360 28212 13412 28218
rect 13360 28154 13412 28160
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 13280 27962 13308 28018
rect 13280 27934 13400 27962
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 13268 27668 13320 27674
rect 13268 27610 13320 27616
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12820 27062 12848 27474
rect 12900 27328 12952 27334
rect 12900 27270 12952 27276
rect 12912 27130 12940 27270
rect 12900 27124 12952 27130
rect 12900 27066 12952 27072
rect 13280 27062 13308 27610
rect 12808 27056 12860 27062
rect 12808 26998 12860 27004
rect 13268 27056 13320 27062
rect 13268 26998 13320 27004
rect 12820 25362 12848 26998
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 13372 25480 13400 27934
rect 13280 25452 13400 25480
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12820 24274 12848 25094
rect 12992 24880 13044 24886
rect 12992 24822 13044 24828
rect 13004 24614 13032 24822
rect 13280 24818 13308 25452
rect 13464 25344 13492 32166
rect 13556 31278 13584 33254
rect 13648 32910 13676 35278
rect 13820 35216 13872 35222
rect 13820 35158 13872 35164
rect 13728 34740 13780 34746
rect 13728 34682 13780 34688
rect 13636 32904 13688 32910
rect 13636 32846 13688 32852
rect 13740 32502 13768 34682
rect 13832 34542 13860 35158
rect 13924 34678 13952 35430
rect 13912 34672 13964 34678
rect 13912 34614 13964 34620
rect 13820 34536 13872 34542
rect 13820 34478 13872 34484
rect 13924 34406 13952 34614
rect 13912 34400 13964 34406
rect 13912 34342 13964 34348
rect 13924 34202 13952 34342
rect 13912 34196 13964 34202
rect 13912 34138 13964 34144
rect 14016 34082 14044 36502
rect 13832 34054 14044 34082
rect 13728 32496 13780 32502
rect 13728 32438 13780 32444
rect 13832 32348 13860 34054
rect 13912 33108 13964 33114
rect 13912 33050 13964 33056
rect 14004 33108 14056 33114
rect 14004 33050 14056 33056
rect 13740 32320 13860 32348
rect 13544 31272 13596 31278
rect 13544 31214 13596 31220
rect 13544 29096 13596 29102
rect 13544 29038 13596 29044
rect 13372 25316 13492 25344
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13372 24410 13400 25316
rect 13452 25220 13504 25226
rect 13452 25162 13504 25168
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12820 22778 12848 23258
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 13096 22778 13124 22918
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 13096 22574 13124 22714
rect 13084 22568 13136 22574
rect 13084 22510 13136 22516
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12636 20454 12756 20482
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12530 17912 12586 17921
rect 12530 17847 12532 17856
rect 12584 17847 12586 17856
rect 12532 17818 12584 17824
rect 12544 17678 12572 17818
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12636 17354 12664 20454
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 13372 20346 13400 21830
rect 13464 20466 13492 25162
rect 13556 24206 13584 29038
rect 13636 29028 13688 29034
rect 13636 28970 13688 28976
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13648 22030 13676 28970
rect 13740 24614 13768 32320
rect 13924 31958 13952 33050
rect 14016 32774 14044 33050
rect 14004 32768 14056 32774
rect 14004 32710 14056 32716
rect 14016 32473 14044 32710
rect 14002 32464 14058 32473
rect 14002 32399 14058 32408
rect 13820 31952 13872 31958
rect 13820 31894 13872 31900
rect 13912 31952 13964 31958
rect 13912 31894 13964 31900
rect 13832 31686 13860 31894
rect 13820 31680 13872 31686
rect 13820 31622 13872 31628
rect 13832 25362 13860 31622
rect 14108 30598 14136 51818
rect 14188 46708 14240 46714
rect 14188 46650 14240 46656
rect 14200 44334 14228 46650
rect 14188 44328 14240 44334
rect 14240 44288 14320 44316
rect 14188 44270 14240 44276
rect 14188 43104 14240 43110
rect 14188 43046 14240 43052
rect 14200 36922 14228 43046
rect 14292 42158 14320 44288
rect 14372 42696 14424 42702
rect 14372 42638 14424 42644
rect 14280 42152 14332 42158
rect 14280 42094 14332 42100
rect 14280 39636 14332 39642
rect 14280 39578 14332 39584
rect 14292 38593 14320 39578
rect 14278 38584 14334 38593
rect 14278 38519 14334 38528
rect 14292 38418 14320 38519
rect 14280 38412 14332 38418
rect 14280 38354 14332 38360
rect 14384 38010 14412 42638
rect 14372 38004 14424 38010
rect 14372 37946 14424 37952
rect 14188 36916 14240 36922
rect 14188 36858 14240 36864
rect 14280 36576 14332 36582
rect 14280 36518 14332 36524
rect 14188 35012 14240 35018
rect 14188 34954 14240 34960
rect 14200 31958 14228 34954
rect 14292 32978 14320 36518
rect 14280 32972 14332 32978
rect 14280 32914 14332 32920
rect 14188 31952 14240 31958
rect 14188 31894 14240 31900
rect 14476 31754 14504 52294
rect 14660 52018 14688 56222
rect 14738 56200 14794 57000
rect 15106 56200 15162 57000
rect 15474 56200 15530 57000
rect 15842 56200 15898 57000
rect 16210 56200 16266 57000
rect 16578 56200 16634 57000
rect 16946 56200 17002 57000
rect 17314 56200 17370 57000
rect 17682 56200 17738 57000
rect 18050 56200 18106 57000
rect 18156 56222 18368 56250
rect 14752 54330 14780 56200
rect 14740 54324 14792 54330
rect 14740 54266 14792 54272
rect 15120 53582 15148 56200
rect 15488 55214 15516 56200
rect 15488 55186 15608 55214
rect 15580 54262 15608 55186
rect 15568 54256 15620 54262
rect 15568 54198 15620 54204
rect 15292 53984 15344 53990
rect 15292 53926 15344 53932
rect 15108 53576 15160 53582
rect 15108 53518 15160 53524
rect 14832 53100 14884 53106
rect 14832 53042 14884 53048
rect 14844 52698 14872 53042
rect 15120 52698 15148 53518
rect 14832 52692 14884 52698
rect 14832 52634 14884 52640
rect 15108 52692 15160 52698
rect 15108 52634 15160 52640
rect 14648 52012 14700 52018
rect 14648 51954 14700 51960
rect 15016 51876 15068 51882
rect 15016 51818 15068 51824
rect 14740 45892 14792 45898
rect 14740 45834 14792 45840
rect 14648 40656 14700 40662
rect 14648 40598 14700 40604
rect 14660 40186 14688 40598
rect 14648 40180 14700 40186
rect 14648 40122 14700 40128
rect 14556 40112 14608 40118
rect 14556 40054 14608 40060
rect 14568 39642 14596 40054
rect 14648 39840 14700 39846
rect 14648 39782 14700 39788
rect 14556 39636 14608 39642
rect 14556 39578 14608 39584
rect 14660 38894 14688 39782
rect 14752 39642 14780 45834
rect 14832 45280 14884 45286
rect 14832 45222 14884 45228
rect 14844 44878 14872 45222
rect 14832 44872 14884 44878
rect 14832 44814 14884 44820
rect 14844 42770 14872 44814
rect 15028 43450 15056 51818
rect 15108 46640 15160 46646
rect 15108 46582 15160 46588
rect 15120 45558 15148 46582
rect 15108 45552 15160 45558
rect 15108 45494 15160 45500
rect 15120 44470 15148 45494
rect 15200 44736 15252 44742
rect 15200 44678 15252 44684
rect 15108 44464 15160 44470
rect 15108 44406 15160 44412
rect 15016 43444 15068 43450
rect 15016 43386 15068 43392
rect 14924 43172 14976 43178
rect 14924 43114 14976 43120
rect 14832 42764 14884 42770
rect 14832 42706 14884 42712
rect 14936 41414 14964 43114
rect 15212 42362 15240 44678
rect 15200 42356 15252 42362
rect 15200 42298 15252 42304
rect 15108 42016 15160 42022
rect 15108 41958 15160 41964
rect 14844 41386 14964 41414
rect 14844 39846 14872 41386
rect 14924 41268 14976 41274
rect 14924 41210 14976 41216
rect 14832 39840 14884 39846
rect 14832 39782 14884 39788
rect 14740 39636 14792 39642
rect 14740 39578 14792 39584
rect 14740 39296 14792 39302
rect 14740 39238 14792 39244
rect 14752 39098 14780 39238
rect 14740 39092 14792 39098
rect 14740 39034 14792 39040
rect 14832 39092 14884 39098
rect 14832 39034 14884 39040
rect 14648 38888 14700 38894
rect 14648 38830 14700 38836
rect 14556 38208 14608 38214
rect 14608 38168 14780 38196
rect 14556 38150 14608 38156
rect 14556 37120 14608 37126
rect 14556 37062 14608 37068
rect 14568 36718 14596 37062
rect 14556 36712 14608 36718
rect 14556 36654 14608 36660
rect 14556 36576 14608 36582
rect 14556 36518 14608 36524
rect 14568 35086 14596 36518
rect 14648 36032 14700 36038
rect 14648 35974 14700 35980
rect 14660 35834 14688 35974
rect 14648 35828 14700 35834
rect 14648 35770 14700 35776
rect 14556 35080 14608 35086
rect 14556 35022 14608 35028
rect 14556 33652 14608 33658
rect 14556 33594 14608 33600
rect 14568 32434 14596 33594
rect 14648 32768 14700 32774
rect 14648 32710 14700 32716
rect 14660 32570 14688 32710
rect 14752 32570 14780 38168
rect 14844 37398 14872 39034
rect 14832 37392 14884 37398
rect 14832 37334 14884 37340
rect 14936 37126 14964 41210
rect 15016 41132 15068 41138
rect 15016 41074 15068 41080
rect 15028 40186 15056 41074
rect 15016 40180 15068 40186
rect 15016 40122 15068 40128
rect 15016 39364 15068 39370
rect 15016 39306 15068 39312
rect 15028 39098 15056 39306
rect 15016 39092 15068 39098
rect 15016 39034 15068 39040
rect 15120 38282 15148 41958
rect 15304 41256 15332 53926
rect 15568 53440 15620 53446
rect 15568 53382 15620 53388
rect 15580 52494 15608 53382
rect 15660 52624 15712 52630
rect 15660 52566 15712 52572
rect 15568 52488 15620 52494
rect 15568 52430 15620 52436
rect 15672 45554 15700 52566
rect 15752 52352 15804 52358
rect 15752 52294 15804 52300
rect 15580 45526 15700 45554
rect 15476 43784 15528 43790
rect 15476 43726 15528 43732
rect 15212 41228 15332 41256
rect 15212 41052 15240 41228
rect 15212 41024 15332 41052
rect 15200 40384 15252 40390
rect 15200 40326 15252 40332
rect 15212 38350 15240 40326
rect 15200 38344 15252 38350
rect 15200 38286 15252 38292
rect 15108 38276 15160 38282
rect 15108 38218 15160 38224
rect 15016 37664 15068 37670
rect 15016 37606 15068 37612
rect 15028 37330 15056 37606
rect 15120 37466 15148 38218
rect 15108 37460 15160 37466
rect 15108 37402 15160 37408
rect 15016 37324 15068 37330
rect 15016 37266 15068 37272
rect 14924 37120 14976 37126
rect 14924 37062 14976 37068
rect 15120 36922 15148 37402
rect 15198 37360 15254 37369
rect 15198 37295 15200 37304
rect 15252 37295 15254 37304
rect 15200 37266 15252 37272
rect 15212 36922 15240 37266
rect 15108 36916 15160 36922
rect 15108 36858 15160 36864
rect 15200 36916 15252 36922
rect 15200 36858 15252 36864
rect 15200 36712 15252 36718
rect 15200 36654 15252 36660
rect 15212 35630 15240 36654
rect 15200 35624 15252 35630
rect 15200 35566 15252 35572
rect 14832 34536 14884 34542
rect 14832 34478 14884 34484
rect 14844 32978 14872 34478
rect 14924 33040 14976 33046
rect 14924 32982 14976 32988
rect 14832 32972 14884 32978
rect 14832 32914 14884 32920
rect 14648 32564 14700 32570
rect 14648 32506 14700 32512
rect 14740 32564 14792 32570
rect 14740 32506 14792 32512
rect 14556 32428 14608 32434
rect 14556 32370 14608 32376
rect 14568 32230 14596 32370
rect 14832 32360 14884 32366
rect 14832 32302 14884 32308
rect 14556 32224 14608 32230
rect 14556 32166 14608 32172
rect 14384 31726 14504 31754
rect 14280 31340 14332 31346
rect 14280 31282 14332 31288
rect 14292 30870 14320 31282
rect 14280 30864 14332 30870
rect 14280 30806 14332 30812
rect 14096 30592 14148 30598
rect 14096 30534 14148 30540
rect 14384 30326 14412 31726
rect 14648 31476 14700 31482
rect 14648 31418 14700 31424
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14372 30320 14424 30326
rect 14372 30262 14424 30268
rect 14476 30258 14504 31078
rect 14464 30252 14516 30258
rect 14464 30194 14516 30200
rect 14464 30048 14516 30054
rect 14464 29990 14516 29996
rect 14476 29850 14504 29990
rect 14464 29844 14516 29850
rect 14464 29786 14516 29792
rect 14556 29776 14608 29782
rect 14556 29718 14608 29724
rect 14464 29708 14516 29714
rect 14464 29650 14516 29656
rect 14004 29640 14056 29646
rect 14004 29582 14056 29588
rect 14016 29170 14044 29582
rect 14004 29164 14056 29170
rect 14004 29106 14056 29112
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14016 28422 14044 29106
rect 14108 28762 14136 29106
rect 14096 28756 14148 28762
rect 14096 28698 14148 28704
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 14016 25786 14044 28358
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14016 25758 14136 25786
rect 13820 25356 13872 25362
rect 13820 25298 13872 25304
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13740 23730 13768 24550
rect 13832 24274 13860 24754
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 13636 22024 13688 22030
rect 13542 21992 13598 22001
rect 13636 21966 13688 21972
rect 13542 21927 13544 21936
rect 13596 21927 13598 21936
rect 13544 21898 13596 21904
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 12728 18834 12756 20334
rect 13372 20318 13492 20346
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13372 18902 13400 20198
rect 13464 19514 13492 20318
rect 13648 20058 13676 21490
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12728 17882 12756 18226
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12544 17326 12664 17354
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12452 15026 12480 17002
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12544 14498 12572 17326
rect 12728 16590 12756 17478
rect 12820 17270 12848 18702
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13372 18426 13400 18566
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 12912 18329 12940 18362
rect 12898 18320 12954 18329
rect 12898 18255 12954 18264
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12912 17134 12940 17818
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 13372 17134 13400 17206
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12820 16658 12848 16730
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12452 14470 12572 14498
rect 12452 14074 12480 14470
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12452 13530 12480 14010
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12544 12434 12572 14282
rect 12636 13852 12664 15370
rect 12728 14618 12756 16050
rect 12820 15366 12848 16594
rect 13372 16182 13400 17070
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13372 15502 13400 16118
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12636 13824 12756 13852
rect 12544 12406 12664 12434
rect 12440 10532 12492 10538
rect 12440 10474 12492 10480
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11808 2746 11928 2774
rect 11808 2106 11836 2746
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 11992 800 12020 2450
rect 12360 800 12388 2518
rect 12452 2446 12480 10474
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12544 3534 12572 3674
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12636 2378 12664 12406
rect 12728 3738 12756 13824
rect 12820 13394 12848 15302
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12820 12170 12848 12854
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12820 11812 12848 12106
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13280 11898 13308 12038
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13176 11824 13228 11830
rect 12820 11784 13176 11812
rect 13176 11766 13228 11772
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 12728 800 12756 3538
rect 13372 3194 13400 12650
rect 13464 10062 13492 19450
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 13648 18154 13676 18634
rect 13636 18148 13688 18154
rect 13636 18090 13688 18096
rect 13544 18080 13596 18086
rect 13596 18028 13676 18034
rect 13544 18022 13676 18028
rect 13556 18006 13676 18022
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13556 16250 13584 17478
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13648 15314 13676 18006
rect 13740 16250 13768 23462
rect 13924 23118 13952 23462
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13832 21690 13860 22578
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13924 21690 13952 22510
rect 14004 22500 14056 22506
rect 14004 22442 14056 22448
rect 14016 21690 14044 22442
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 14108 21570 14136 25758
rect 14200 25498 14228 26930
rect 14292 26382 14320 28358
rect 14372 26784 14424 26790
rect 14372 26726 14424 26732
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14384 25838 14412 26726
rect 14476 25838 14504 29650
rect 14372 25832 14424 25838
rect 14372 25774 14424 25780
rect 14464 25832 14516 25838
rect 14464 25774 14516 25780
rect 14188 25492 14240 25498
rect 14188 25434 14240 25440
rect 14188 25356 14240 25362
rect 14188 25298 14240 25304
rect 14016 21542 14136 21570
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13832 18766 13860 21286
rect 14016 20262 14044 21542
rect 14200 21146 14228 25298
rect 14384 24750 14412 25774
rect 14476 25430 14504 25774
rect 14464 25424 14516 25430
rect 14464 25366 14516 25372
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14568 24138 14596 29718
rect 14660 29102 14688 31418
rect 14844 30190 14872 32302
rect 14936 31686 14964 32982
rect 15108 32496 15160 32502
rect 15108 32438 15160 32444
rect 15120 31890 15148 32438
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15108 31884 15160 31890
rect 15108 31826 15160 31832
rect 14924 31680 14976 31686
rect 14924 31622 14976 31628
rect 15212 30802 15240 32166
rect 15304 31142 15332 41024
rect 15384 40996 15436 41002
rect 15384 40938 15436 40944
rect 15396 39982 15424 40938
rect 15384 39976 15436 39982
rect 15384 39918 15436 39924
rect 15384 39296 15436 39302
rect 15384 39238 15436 39244
rect 15396 36378 15424 39238
rect 15488 38876 15516 43726
rect 15580 43110 15608 45526
rect 15660 44804 15712 44810
rect 15660 44746 15712 44752
rect 15672 43246 15700 44746
rect 15660 43240 15712 43246
rect 15660 43182 15712 43188
rect 15568 43104 15620 43110
rect 15568 43046 15620 43052
rect 15568 42900 15620 42906
rect 15568 42842 15620 42848
rect 15580 42634 15608 42842
rect 15568 42628 15620 42634
rect 15568 42570 15620 42576
rect 15568 42288 15620 42294
rect 15568 42230 15620 42236
rect 15580 40186 15608 42230
rect 15568 40180 15620 40186
rect 15568 40122 15620 40128
rect 15672 39506 15700 43182
rect 15660 39500 15712 39506
rect 15660 39442 15712 39448
rect 15568 38888 15620 38894
rect 15488 38848 15568 38876
rect 15568 38830 15620 38836
rect 15476 38004 15528 38010
rect 15476 37946 15528 37952
rect 15488 37126 15516 37946
rect 15580 37806 15608 38830
rect 15660 38276 15712 38282
rect 15660 38218 15712 38224
rect 15568 37800 15620 37806
rect 15568 37742 15620 37748
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 15488 36961 15516 37062
rect 15474 36952 15530 36961
rect 15474 36887 15530 36896
rect 15384 36372 15436 36378
rect 15384 36314 15436 36320
rect 15672 36242 15700 38218
rect 15660 36236 15712 36242
rect 15660 36178 15712 36184
rect 15658 36136 15714 36145
rect 15658 36071 15660 36080
rect 15712 36071 15714 36080
rect 15660 36042 15712 36048
rect 15764 35306 15792 52294
rect 15856 52018 15884 56200
rect 16224 53582 16252 56200
rect 16592 53786 16620 56200
rect 16580 53780 16632 53786
rect 16580 53722 16632 53728
rect 16960 53582 16988 56200
rect 16212 53576 16264 53582
rect 16212 53518 16264 53524
rect 16948 53576 17000 53582
rect 16948 53518 17000 53524
rect 16224 52698 16252 53518
rect 16856 53440 16908 53446
rect 16856 53382 16908 53388
rect 16396 52964 16448 52970
rect 16396 52906 16448 52912
rect 16212 52692 16264 52698
rect 16212 52634 16264 52640
rect 16408 52601 16436 52906
rect 16394 52592 16450 52601
rect 16394 52527 16450 52536
rect 16868 52494 16896 53382
rect 17040 52896 17092 52902
rect 17040 52838 17092 52844
rect 16856 52488 16908 52494
rect 16856 52430 16908 52436
rect 15844 52012 15896 52018
rect 15844 51954 15896 51960
rect 16304 47524 16356 47530
rect 16304 47466 16356 47472
rect 16316 46374 16344 47466
rect 16580 47456 16632 47462
rect 16580 47398 16632 47404
rect 16396 46980 16448 46986
rect 16396 46922 16448 46928
rect 16408 46646 16436 46922
rect 16396 46640 16448 46646
rect 16396 46582 16448 46588
rect 16304 46368 16356 46374
rect 16304 46310 16356 46316
rect 16316 45422 16344 46310
rect 16408 45830 16436 46582
rect 16396 45824 16448 45830
rect 16396 45766 16448 45772
rect 16304 45416 16356 45422
rect 16304 45358 16356 45364
rect 16408 45354 16436 45766
rect 15844 45348 15896 45354
rect 15844 45290 15896 45296
rect 16396 45348 16448 45354
rect 16396 45290 16448 45296
rect 15856 44810 15884 45290
rect 16120 45280 16172 45286
rect 16120 45222 16172 45228
rect 15844 44804 15896 44810
rect 15844 44746 15896 44752
rect 15856 44470 15884 44746
rect 15844 44464 15896 44470
rect 15844 44406 15896 44412
rect 15844 43104 15896 43110
rect 15842 43072 15844 43081
rect 15896 43072 15898 43081
rect 15842 43007 15898 43016
rect 15844 42900 15896 42906
rect 15844 42842 15896 42848
rect 15856 41274 15884 42842
rect 16132 41682 16160 45222
rect 16408 45082 16436 45290
rect 16396 45076 16448 45082
rect 16396 45018 16448 45024
rect 16396 44532 16448 44538
rect 16396 44474 16448 44480
rect 16408 42634 16436 44474
rect 16488 44192 16540 44198
rect 16488 44134 16540 44140
rect 16396 42628 16448 42634
rect 16396 42570 16448 42576
rect 16500 42090 16528 44134
rect 16488 42084 16540 42090
rect 16488 42026 16540 42032
rect 16120 41676 16172 41682
rect 16120 41618 16172 41624
rect 16212 41472 16264 41478
rect 16212 41414 16264 41420
rect 15844 41268 15896 41274
rect 15844 41210 15896 41216
rect 15844 40452 15896 40458
rect 15844 40394 15896 40400
rect 15856 39574 15884 40394
rect 16028 39976 16080 39982
rect 16028 39918 16080 39924
rect 16040 39574 16068 39918
rect 15844 39568 15896 39574
rect 15844 39510 15896 39516
rect 16028 39568 16080 39574
rect 16028 39510 16080 39516
rect 15844 39432 15896 39438
rect 16040 39386 16068 39510
rect 15844 39374 15896 39380
rect 15856 38554 15884 39374
rect 15948 39358 16068 39386
rect 15948 39098 15976 39358
rect 16028 39296 16080 39302
rect 16028 39238 16080 39244
rect 16040 39098 16068 39238
rect 15936 39092 15988 39098
rect 15936 39034 15988 39040
rect 16028 39092 16080 39098
rect 16028 39034 16080 39040
rect 16028 38752 16080 38758
rect 16026 38720 16028 38729
rect 16080 38720 16082 38729
rect 16026 38655 16082 38664
rect 15844 38548 15896 38554
rect 15844 38490 15896 38496
rect 15936 38344 15988 38350
rect 15936 38286 15988 38292
rect 15844 36712 15896 36718
rect 15842 36680 15844 36689
rect 15896 36680 15898 36689
rect 15842 36615 15898 36624
rect 15948 35494 15976 38286
rect 16118 38040 16174 38049
rect 16118 37975 16120 37984
rect 16172 37975 16174 37984
rect 16120 37946 16172 37952
rect 16120 37800 16172 37806
rect 16120 37742 16172 37748
rect 16028 36644 16080 36650
rect 16028 36586 16080 36592
rect 15936 35488 15988 35494
rect 15936 35430 15988 35436
rect 15672 35278 15792 35306
rect 15672 35034 15700 35278
rect 15948 35170 15976 35430
rect 15764 35154 15976 35170
rect 15752 35148 15976 35154
rect 15804 35142 15976 35148
rect 15752 35090 15804 35096
rect 15672 35006 15792 35034
rect 15476 34400 15528 34406
rect 15476 34342 15528 34348
rect 15568 34400 15620 34406
rect 15568 34342 15620 34348
rect 15488 33522 15516 34342
rect 15476 33516 15528 33522
rect 15476 33458 15528 33464
rect 15488 33386 15516 33458
rect 15476 33380 15528 33386
rect 15476 33322 15528 33328
rect 15384 31408 15436 31414
rect 15384 31350 15436 31356
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15200 30796 15252 30802
rect 15200 30738 15252 30744
rect 14832 30184 14884 30190
rect 14832 30126 14884 30132
rect 15304 29646 15332 31078
rect 15396 30598 15424 31350
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15384 30592 15436 30598
rect 15384 30534 15436 30540
rect 15292 29640 15344 29646
rect 15292 29582 15344 29588
rect 14740 29572 14792 29578
rect 14740 29514 14792 29520
rect 14648 29096 14700 29102
rect 14648 29038 14700 29044
rect 14752 28393 14780 29514
rect 15108 29504 15160 29510
rect 15108 29446 15160 29452
rect 14832 28620 14884 28626
rect 14832 28562 14884 28568
rect 14738 28384 14794 28393
rect 14738 28319 14794 28328
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 14648 26580 14700 26586
rect 14648 26522 14700 26528
rect 14660 26246 14688 26522
rect 14648 26240 14700 26246
rect 14648 26182 14700 26188
rect 14660 25974 14688 26182
rect 14648 25968 14700 25974
rect 14648 25910 14700 25916
rect 14660 25226 14688 25910
rect 14648 25220 14700 25226
rect 14648 25162 14700 25168
rect 14648 24812 14700 24818
rect 14648 24754 14700 24760
rect 14660 24614 14688 24754
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14660 24342 14688 24550
rect 14648 24336 14700 24342
rect 14648 24278 14700 24284
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 14292 22098 14320 23122
rect 14280 22092 14332 22098
rect 14280 22034 14332 22040
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14200 20942 14228 21082
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 14004 20256 14056 20262
rect 14004 20198 14056 20204
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 14004 19440 14056 19446
rect 14004 19382 14056 19388
rect 14016 19310 14044 19382
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13740 15502 13768 16186
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13648 15286 13768 15314
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13648 14346 13676 14826
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13542 14104 13598 14113
rect 13542 14039 13598 14048
rect 13556 14006 13584 14039
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13544 13796 13596 13802
rect 13544 13738 13596 13744
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13096 870 13216 898
rect 13096 800 13124 870
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13188 762 13216 870
rect 13372 762 13400 2926
rect 13464 800 13492 4014
rect 13556 3058 13584 13738
rect 13648 4146 13676 13806
rect 13740 12714 13768 15286
rect 13924 12918 13952 18838
rect 14016 18086 14044 19246
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13924 12442 13952 12854
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13740 3126 13768 12038
rect 14016 11354 14044 13194
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14108 5574 14136 20198
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14200 18970 14228 19722
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14200 17066 14228 18770
rect 14188 17060 14240 17066
rect 14188 17002 14240 17008
rect 14200 15570 14228 17002
rect 14292 16726 14320 20742
rect 14280 16720 14332 16726
rect 14280 16662 14332 16668
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14292 13802 14320 15846
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14384 12918 14412 23598
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14568 21962 14596 23258
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14568 21486 14596 21898
rect 14646 21720 14702 21729
rect 14752 21690 14780 26726
rect 14844 26314 14872 28562
rect 14924 28416 14976 28422
rect 14924 28358 14976 28364
rect 14936 27878 14964 28358
rect 14924 27872 14976 27878
rect 14924 27814 14976 27820
rect 14832 26308 14884 26314
rect 14832 26250 14884 26256
rect 14936 26194 14964 27814
rect 15016 27328 15068 27334
rect 15016 27270 15068 27276
rect 14844 26166 14964 26194
rect 14844 24562 14872 26166
rect 14924 25152 14976 25158
rect 14924 25094 14976 25100
rect 14936 24682 14964 25094
rect 15028 24818 15056 27270
rect 15120 27130 15148 29446
rect 15396 29102 15424 30534
rect 15488 30326 15516 30670
rect 15476 30320 15528 30326
rect 15476 30262 15528 30268
rect 15384 29096 15436 29102
rect 15304 29056 15384 29084
rect 15200 28960 15252 28966
rect 15200 28902 15252 28908
rect 15212 28558 15240 28902
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 15304 28422 15332 29056
rect 15384 29038 15436 29044
rect 15488 28490 15516 30262
rect 15580 29306 15608 34342
rect 15660 31816 15712 31822
rect 15660 31758 15712 31764
rect 15568 29300 15620 29306
rect 15568 29242 15620 29248
rect 15476 28484 15528 28490
rect 15476 28426 15528 28432
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15304 28257 15332 28358
rect 15290 28248 15346 28257
rect 15290 28183 15346 28192
rect 15476 28212 15528 28218
rect 15476 28154 15528 28160
rect 15384 27396 15436 27402
rect 15384 27338 15436 27344
rect 15396 27305 15424 27338
rect 15382 27296 15438 27305
rect 15382 27231 15438 27240
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 15384 26376 15436 26382
rect 15384 26318 15436 26324
rect 15396 26042 15424 26318
rect 15384 26036 15436 26042
rect 15384 25978 15436 25984
rect 15108 25696 15160 25702
rect 15108 25638 15160 25644
rect 15016 24812 15068 24818
rect 15016 24754 15068 24760
rect 14924 24676 14976 24682
rect 14924 24618 14976 24624
rect 14844 24534 14964 24562
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 14646 21655 14702 21664
rect 14740 21684 14792 21690
rect 14660 21486 14688 21655
rect 14740 21626 14792 21632
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14660 20262 14688 21422
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14648 19984 14700 19990
rect 14648 19926 14700 19932
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14476 19310 14504 19858
rect 14660 19786 14688 19926
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 14740 19712 14792 19718
rect 14738 19680 14740 19689
rect 14792 19680 14794 19689
rect 14738 19615 14794 19624
rect 14844 19378 14872 23802
rect 14936 23662 14964 24534
rect 14924 23656 14976 23662
rect 14924 23598 14976 23604
rect 15120 22778 15148 25638
rect 15396 25362 15424 25978
rect 15384 25356 15436 25362
rect 15304 25316 15384 25344
rect 15200 24404 15252 24410
rect 15200 24346 15252 24352
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15212 20874 15240 24346
rect 15304 23186 15332 25316
rect 15384 25298 15436 25304
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15488 23066 15516 28154
rect 15568 27872 15620 27878
rect 15568 27814 15620 27820
rect 15580 26042 15608 27814
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 15672 24410 15700 31758
rect 15764 28506 15792 35006
rect 15844 34468 15896 34474
rect 15844 34410 15896 34416
rect 15856 33318 15884 34410
rect 15948 34066 15976 35142
rect 15936 34060 15988 34066
rect 15936 34002 15988 34008
rect 15948 33658 15976 34002
rect 15936 33652 15988 33658
rect 15936 33594 15988 33600
rect 15936 33516 15988 33522
rect 15936 33458 15988 33464
rect 15948 33386 15976 33458
rect 15936 33380 15988 33386
rect 15936 33322 15988 33328
rect 15844 33312 15896 33318
rect 15844 33254 15896 33260
rect 15844 32836 15896 32842
rect 15844 32778 15896 32784
rect 15856 30122 15884 32778
rect 15948 32434 15976 33322
rect 15936 32428 15988 32434
rect 15936 32370 15988 32376
rect 15948 31346 15976 32370
rect 15936 31340 15988 31346
rect 15936 31282 15988 31288
rect 15948 30870 15976 31282
rect 15936 30864 15988 30870
rect 15936 30806 15988 30812
rect 15948 30734 15976 30806
rect 15936 30728 15988 30734
rect 15936 30670 15988 30676
rect 15844 30116 15896 30122
rect 15844 30058 15896 30064
rect 16040 29850 16068 36586
rect 16132 35290 16160 37742
rect 16224 37330 16252 41414
rect 16396 40996 16448 41002
rect 16396 40938 16448 40944
rect 16304 40384 16356 40390
rect 16304 40326 16356 40332
rect 16316 40186 16344 40326
rect 16304 40180 16356 40186
rect 16304 40122 16356 40128
rect 16304 40044 16356 40050
rect 16304 39986 16356 39992
rect 16316 39846 16344 39986
rect 16304 39840 16356 39846
rect 16304 39782 16356 39788
rect 16316 37874 16344 39782
rect 16304 37868 16356 37874
rect 16304 37810 16356 37816
rect 16316 37670 16344 37810
rect 16304 37664 16356 37670
rect 16304 37606 16356 37612
rect 16316 37466 16344 37606
rect 16304 37460 16356 37466
rect 16304 37402 16356 37408
rect 16408 37398 16436 40938
rect 16500 37874 16528 42026
rect 16592 41614 16620 47398
rect 16672 47116 16724 47122
rect 16672 47058 16724 47064
rect 16948 47116 17000 47122
rect 16948 47058 17000 47064
rect 16684 47002 16712 47058
rect 16684 46974 16896 47002
rect 16868 46510 16896 46974
rect 16856 46504 16908 46510
rect 16856 46446 16908 46452
rect 16868 44946 16896 46446
rect 16856 44940 16908 44946
rect 16856 44882 16908 44888
rect 16764 44872 16816 44878
rect 16764 44814 16816 44820
rect 16672 43104 16724 43110
rect 16672 43046 16724 43052
rect 16684 42906 16712 43046
rect 16672 42900 16724 42906
rect 16672 42842 16724 42848
rect 16672 42560 16724 42566
rect 16672 42502 16724 42508
rect 16580 41608 16632 41614
rect 16580 41550 16632 41556
rect 16684 41070 16712 42502
rect 16672 41064 16724 41070
rect 16672 41006 16724 41012
rect 16580 38752 16632 38758
rect 16580 38694 16632 38700
rect 16488 37868 16540 37874
rect 16488 37810 16540 37816
rect 16396 37392 16448 37398
rect 16396 37334 16448 37340
rect 16212 37324 16264 37330
rect 16212 37266 16264 37272
rect 16396 37120 16448 37126
rect 16396 37062 16448 37068
rect 16120 35284 16172 35290
rect 16120 35226 16172 35232
rect 16212 33924 16264 33930
rect 16212 33866 16264 33872
rect 16120 32768 16172 32774
rect 16120 32710 16172 32716
rect 16132 32298 16160 32710
rect 16120 32292 16172 32298
rect 16120 32234 16172 32240
rect 16224 31482 16252 33866
rect 16304 33856 16356 33862
rect 16304 33798 16356 33804
rect 16316 33454 16344 33798
rect 16304 33448 16356 33454
rect 16304 33390 16356 33396
rect 16316 32366 16344 33390
rect 16304 32360 16356 32366
rect 16304 32302 16356 32308
rect 16408 31754 16436 37062
rect 16592 34678 16620 38694
rect 16672 38004 16724 38010
rect 16672 37946 16724 37952
rect 16684 37806 16712 37946
rect 16672 37800 16724 37806
rect 16672 37742 16724 37748
rect 16670 36816 16726 36825
rect 16670 36751 16672 36760
rect 16724 36751 16726 36760
rect 16672 36722 16724 36728
rect 16580 34672 16632 34678
rect 16580 34614 16632 34620
rect 16488 32972 16540 32978
rect 16488 32914 16540 32920
rect 16316 31726 16436 31754
rect 16212 31476 16264 31482
rect 16212 31418 16264 31424
rect 16120 30660 16172 30666
rect 16120 30602 16172 30608
rect 16132 30394 16160 30602
rect 16120 30388 16172 30394
rect 16120 30330 16172 30336
rect 16316 30326 16344 31726
rect 16500 30802 16528 32914
rect 16776 32910 16804 44814
rect 16868 44334 16896 44882
rect 16960 44878 16988 47058
rect 16948 44872 17000 44878
rect 16948 44814 17000 44820
rect 16856 44328 16908 44334
rect 16856 44270 16908 44276
rect 17052 43194 17080 52838
rect 17132 52692 17184 52698
rect 17132 52634 17184 52640
rect 17144 52601 17172 52634
rect 17130 52592 17186 52601
rect 17130 52527 17186 52536
rect 17328 52018 17356 56200
rect 17408 54188 17460 54194
rect 17408 54130 17460 54136
rect 17420 53242 17448 54130
rect 17500 53984 17552 53990
rect 17500 53926 17552 53932
rect 17408 53236 17460 53242
rect 17408 53178 17460 53184
rect 17512 53174 17540 53926
rect 17696 53718 17724 56200
rect 18064 56114 18092 56200
rect 18156 56114 18184 56222
rect 18064 56086 18184 56114
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 17960 54188 18012 54194
rect 17960 54130 18012 54136
rect 17972 53786 18000 54130
rect 17960 53780 18012 53786
rect 17960 53722 18012 53728
rect 17684 53712 17736 53718
rect 17684 53654 17736 53660
rect 17684 53576 17736 53582
rect 17684 53518 17736 53524
rect 17592 53440 17644 53446
rect 17592 53382 17644 53388
rect 17500 53168 17552 53174
rect 17500 53110 17552 53116
rect 17604 52494 17632 53382
rect 17696 53242 17724 53518
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17684 53236 17736 53242
rect 17684 53178 17736 53184
rect 18340 53106 18368 56222
rect 18418 56200 18474 57000
rect 18786 56200 18842 57000
rect 19154 56200 19210 57000
rect 19522 56200 19578 57000
rect 19890 56200 19946 57000
rect 20258 56200 20314 57000
rect 20626 56200 20682 57000
rect 20994 56200 21050 57000
rect 21362 56200 21418 57000
rect 21730 56200 21786 57000
rect 22098 56200 22154 57000
rect 22466 56200 22522 57000
rect 22834 56200 22890 57000
rect 23202 56200 23258 57000
rect 23570 56200 23626 57000
rect 24582 56264 24638 56273
rect 18432 53786 18460 56200
rect 18800 55214 18828 56200
rect 18800 55186 18920 55214
rect 18696 54120 18748 54126
rect 18696 54062 18748 54068
rect 18604 53984 18656 53990
rect 18604 53926 18656 53932
rect 18420 53780 18472 53786
rect 18420 53722 18472 53728
rect 18616 53174 18644 53926
rect 18708 53650 18736 54062
rect 18696 53644 18748 53650
rect 18696 53586 18748 53592
rect 18604 53168 18656 53174
rect 18604 53110 18656 53116
rect 18328 53100 18380 53106
rect 18328 53042 18380 53048
rect 18788 52896 18840 52902
rect 18788 52838 18840 52844
rect 18800 52494 18828 52838
rect 17592 52488 17644 52494
rect 17592 52430 17644 52436
rect 18788 52488 18840 52494
rect 18788 52430 18840 52436
rect 18512 52352 18564 52358
rect 18512 52294 18564 52300
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17316 52012 17368 52018
rect 17316 51954 17368 51960
rect 17224 51876 17276 51882
rect 17224 51818 17276 51824
rect 18420 51876 18472 51882
rect 18420 51818 18472 51824
rect 17236 47802 17264 51818
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 18328 49088 18380 49094
rect 18328 49030 18380 49036
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17316 48272 17368 48278
rect 17316 48214 17368 48220
rect 17328 47802 17356 48214
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17224 47796 17276 47802
rect 17224 47738 17276 47744
rect 17316 47796 17368 47802
rect 17316 47738 17368 47744
rect 17328 47410 17356 47738
rect 16868 43166 17080 43194
rect 17144 47382 17356 47410
rect 17500 47456 17552 47462
rect 17500 47398 17552 47404
rect 16868 40526 16896 43166
rect 17040 43104 17092 43110
rect 17040 43046 17092 43052
rect 17052 40594 17080 43046
rect 16948 40588 17000 40594
rect 16948 40530 17000 40536
rect 17040 40588 17092 40594
rect 17040 40530 17092 40536
rect 16856 40520 16908 40526
rect 16856 40462 16908 40468
rect 16868 40089 16896 40462
rect 16854 40080 16910 40089
rect 16854 40015 16910 40024
rect 16856 38888 16908 38894
rect 16856 38830 16908 38836
rect 16868 38010 16896 38830
rect 16856 38004 16908 38010
rect 16856 37946 16908 37952
rect 16960 36310 16988 40530
rect 17144 39953 17172 47382
rect 17316 47116 17368 47122
rect 17316 47058 17368 47064
rect 17224 46368 17276 46374
rect 17224 46310 17276 46316
rect 17236 44742 17264 46310
rect 17224 44736 17276 44742
rect 17224 44678 17276 44684
rect 17236 40594 17264 44678
rect 17328 43246 17356 47058
rect 17408 43648 17460 43654
rect 17408 43590 17460 43596
rect 17420 43450 17448 43590
rect 17512 43450 17540 47398
rect 17592 46912 17644 46918
rect 17592 46854 17644 46860
rect 17604 46646 17632 46854
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17592 46640 17644 46646
rect 17592 46582 17644 46588
rect 17604 46170 17632 46582
rect 17592 46164 17644 46170
rect 17592 46106 17644 46112
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 18340 45554 18368 49030
rect 18432 47802 18460 51818
rect 18524 47802 18552 52294
rect 18892 52018 18920 55186
rect 19168 54126 19196 56200
rect 19432 54188 19484 54194
rect 19432 54130 19484 54136
rect 19156 54120 19208 54126
rect 19156 54062 19208 54068
rect 19340 53984 19392 53990
rect 19340 53926 19392 53932
rect 19352 53174 19380 53926
rect 19444 53446 19472 54130
rect 19536 53582 19564 56200
rect 19524 53576 19576 53582
rect 19524 53518 19576 53524
rect 19432 53440 19484 53446
rect 19432 53382 19484 53388
rect 19340 53168 19392 53174
rect 19340 53110 19392 53116
rect 19904 53106 19932 56200
rect 20168 53440 20220 53446
rect 20168 53382 20220 53388
rect 19892 53100 19944 53106
rect 19892 53042 19944 53048
rect 19432 52896 19484 52902
rect 19432 52838 19484 52844
rect 18880 52012 18932 52018
rect 18880 51954 18932 51960
rect 18604 51808 18656 51814
rect 18604 51750 18656 51756
rect 18420 47796 18472 47802
rect 18420 47738 18472 47744
rect 18512 47796 18564 47802
rect 18512 47738 18564 47744
rect 18524 47705 18552 47738
rect 18510 47696 18566 47705
rect 18510 47631 18566 47640
rect 18420 47592 18472 47598
rect 18420 47534 18472 47540
rect 18432 47258 18460 47534
rect 18420 47252 18472 47258
rect 18420 47194 18472 47200
rect 18432 46714 18460 47194
rect 18512 47184 18564 47190
rect 18512 47126 18564 47132
rect 18420 46708 18472 46714
rect 18420 46650 18472 46656
rect 18340 45526 18460 45554
rect 18328 45416 18380 45422
rect 18328 45358 18380 45364
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 18340 44198 18368 45358
rect 18328 44192 18380 44198
rect 18328 44134 18380 44140
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17408 43444 17460 43450
rect 17408 43386 17460 43392
rect 17500 43444 17552 43450
rect 17500 43386 17552 43392
rect 18340 43246 18368 44134
rect 17316 43240 17368 43246
rect 17316 43182 17368 43188
rect 18328 43240 18380 43246
rect 18328 43182 18380 43188
rect 18144 43172 18196 43178
rect 18144 43114 18196 43120
rect 18156 42770 18184 43114
rect 18432 42770 18460 45526
rect 18144 42764 18196 42770
rect 18144 42706 18196 42712
rect 18420 42764 18472 42770
rect 18420 42706 18472 42712
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 17868 42288 17920 42294
rect 17868 42230 17920 42236
rect 17684 40724 17736 40730
rect 17684 40666 17736 40672
rect 17224 40588 17276 40594
rect 17224 40530 17276 40536
rect 17500 40384 17552 40390
rect 17500 40326 17552 40332
rect 17130 39944 17186 39953
rect 17130 39879 17186 39888
rect 17132 39840 17184 39846
rect 17132 39782 17184 39788
rect 17040 39364 17092 39370
rect 17040 39306 17092 39312
rect 17052 36922 17080 39306
rect 17040 36916 17092 36922
rect 17040 36858 17092 36864
rect 16948 36304 17000 36310
rect 16948 36246 17000 36252
rect 17144 36156 17172 39782
rect 17314 38584 17370 38593
rect 17314 38519 17370 38528
rect 17328 38350 17356 38519
rect 17316 38344 17368 38350
rect 17316 38286 17368 38292
rect 17328 38010 17356 38286
rect 17316 38004 17368 38010
rect 17316 37946 17368 37952
rect 17408 37868 17460 37874
rect 17408 37810 17460 37816
rect 17316 37120 17368 37126
rect 17316 37062 17368 37068
rect 17328 36854 17356 37062
rect 17316 36848 17368 36854
rect 17316 36790 17368 36796
rect 17224 36576 17276 36582
rect 17224 36518 17276 36524
rect 16960 36128 17172 36156
rect 16960 34202 16988 36128
rect 16948 34196 17000 34202
rect 16948 34138 17000 34144
rect 16764 32904 16816 32910
rect 16764 32846 16816 32852
rect 16578 32464 16634 32473
rect 16578 32399 16634 32408
rect 16488 30796 16540 30802
rect 16488 30738 16540 30744
rect 16592 30410 16620 32399
rect 16672 32224 16724 32230
rect 16672 32166 16724 32172
rect 16408 30382 16620 30410
rect 16304 30320 16356 30326
rect 16304 30262 16356 30268
rect 16212 30184 16264 30190
rect 16212 30126 16264 30132
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 16118 29200 16174 29209
rect 16118 29135 16174 29144
rect 16028 28960 16080 28966
rect 16028 28902 16080 28908
rect 15764 28478 15884 28506
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15304 23038 15516 23066
rect 15304 22710 15332 23038
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15396 22778 15424 22918
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15200 20868 15252 20874
rect 15200 20810 15252 20816
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14476 18222 14504 19246
rect 14660 19174 14688 19314
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14476 16998 14504 17682
rect 14660 17678 14688 19110
rect 14844 18834 14872 19110
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14752 17542 14780 18022
rect 14844 17746 14872 18770
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 15028 17066 15056 18226
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15120 17678 15148 17818
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15120 17270 15148 17614
rect 15108 17264 15160 17270
rect 15108 17206 15160 17212
rect 15016 17060 15068 17066
rect 15016 17002 15068 17008
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14476 14482 14504 16934
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14738 16280 14794 16289
rect 14738 16215 14740 16224
rect 14792 16215 14794 16224
rect 14740 16186 14792 16192
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14568 14550 14596 14962
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 14292 3058 14320 12650
rect 14476 12442 14504 13262
rect 14844 13258 14872 14894
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14568 11626 14596 13194
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13832 800 13860 2314
rect 14200 800 14228 2926
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14568 800 14596 2450
rect 14660 2446 14688 12650
rect 14844 10674 14872 12718
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14936 3754 14964 16594
rect 14844 3726 14964 3754
rect 14844 3534 14872 3726
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14936 800 14964 3538
rect 15028 2310 15056 17002
rect 15304 16538 15332 22646
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15396 21486 15424 21830
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 15396 18222 15424 21422
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15212 16510 15332 16538
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15120 11898 15148 13670
rect 15212 12918 15240 16510
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15304 15502 15332 16390
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15396 15094 15424 17478
rect 15488 15434 15516 22918
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15580 17678 15608 22374
rect 15764 20942 15792 28358
rect 15856 27878 15884 28478
rect 15934 28248 15990 28257
rect 15934 28183 15936 28192
rect 15988 28183 15990 28192
rect 15936 28154 15988 28160
rect 16040 28098 16068 28902
rect 16132 28506 16160 29135
rect 16224 28626 16252 30126
rect 16304 29640 16356 29646
rect 16304 29582 16356 29588
rect 16316 29050 16344 29582
rect 16408 29306 16436 30382
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16580 29844 16632 29850
rect 16580 29786 16632 29792
rect 16396 29300 16448 29306
rect 16396 29242 16448 29248
rect 16394 29064 16450 29073
rect 16316 29022 16394 29050
rect 16394 28999 16396 29008
rect 16448 28999 16450 29008
rect 16396 28970 16448 28976
rect 16396 28688 16448 28694
rect 16396 28630 16448 28636
rect 16212 28620 16264 28626
rect 16212 28562 16264 28568
rect 16132 28478 16344 28506
rect 15936 28076 15988 28082
rect 16040 28070 16252 28098
rect 15936 28018 15988 28024
rect 15844 27872 15896 27878
rect 15844 27814 15896 27820
rect 15844 27464 15896 27470
rect 15844 27406 15896 27412
rect 15856 22982 15884 27406
rect 15948 23202 15976 28018
rect 16028 28008 16080 28014
rect 16026 27976 16028 27985
rect 16080 27976 16082 27985
rect 16026 27911 16082 27920
rect 16028 25832 16080 25838
rect 16028 25774 16080 25780
rect 16040 23322 16068 25774
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 15948 23174 16068 23202
rect 15936 23044 15988 23050
rect 15936 22986 15988 22992
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15948 22574 15976 22986
rect 16040 22778 16068 23174
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 16132 22710 16160 23054
rect 16224 22982 16252 28070
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 16120 22704 16172 22710
rect 16316 22692 16344 28478
rect 16408 28150 16436 28630
rect 16396 28144 16448 28150
rect 16396 28086 16448 28092
rect 16500 23594 16528 29786
rect 16592 29578 16620 29786
rect 16580 29572 16632 29578
rect 16580 29514 16632 29520
rect 16592 25106 16620 29514
rect 16684 28490 16712 32166
rect 16776 31822 16804 32846
rect 17236 32502 17264 36518
rect 17420 35766 17448 37810
rect 17408 35760 17460 35766
rect 17408 35702 17460 35708
rect 17408 35624 17460 35630
rect 17408 35566 17460 35572
rect 17316 34604 17368 34610
rect 17316 34546 17368 34552
rect 17224 32496 17276 32502
rect 17224 32438 17276 32444
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 17224 31680 17276 31686
rect 17224 31622 17276 31628
rect 17040 31272 17092 31278
rect 17040 31214 17092 31220
rect 16764 29776 16816 29782
rect 16764 29718 16816 29724
rect 16776 29170 16804 29718
rect 16764 29164 16816 29170
rect 16764 29106 16816 29112
rect 16856 28960 16908 28966
rect 16856 28902 16908 28908
rect 16868 28558 16896 28902
rect 16856 28552 16908 28558
rect 16856 28494 16908 28500
rect 16672 28484 16724 28490
rect 16672 28426 16724 28432
rect 16764 28416 16816 28422
rect 16762 28384 16764 28393
rect 16948 28416 17000 28422
rect 16816 28384 16818 28393
rect 16948 28358 17000 28364
rect 16762 28319 16818 28328
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16684 25362 16712 26522
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16592 25078 16712 25106
rect 16488 23588 16540 23594
rect 16488 23530 16540 23536
rect 16500 23474 16528 23530
rect 16500 23446 16620 23474
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16408 23118 16436 23258
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16488 22976 16540 22982
rect 16488 22918 16540 22924
rect 16316 22664 16436 22692
rect 16120 22646 16172 22652
rect 15936 22568 15988 22574
rect 15936 22510 15988 22516
rect 15948 22094 15976 22510
rect 16132 22234 16160 22646
rect 16408 22386 16436 22664
rect 16316 22358 16436 22386
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 16120 22094 16172 22098
rect 15948 22092 16172 22094
rect 15948 22066 16120 22092
rect 16120 22034 16172 22040
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15948 21418 15976 21830
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16212 21548 16264 21554
rect 16212 21490 16264 21496
rect 15936 21412 15988 21418
rect 15936 21354 15988 21360
rect 16132 20942 16160 21490
rect 16224 21078 16252 21490
rect 16212 21072 16264 21078
rect 16212 21014 16264 21020
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 16118 20768 16174 20777
rect 15672 17678 15700 20742
rect 16118 20703 16174 20712
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 16040 16658 16068 18158
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 15934 16280 15990 16289
rect 15934 16215 15990 16224
rect 15948 16182 15976 16215
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15396 14618 15424 15030
rect 15488 15026 15516 15370
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15396 13394 15424 14418
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15304 12986 15332 13194
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15120 11218 15148 11698
rect 15304 11218 15332 12242
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15212 10470 15240 11018
rect 15304 10810 15332 11154
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 4758 15240 10406
rect 15200 4752 15252 4758
rect 15200 4694 15252 4700
rect 15488 3466 15516 12582
rect 15580 3534 15608 15846
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15672 12442 15700 15302
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15764 12986 15792 14214
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15764 11898 15792 12922
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15856 6798 15884 14554
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15948 13530 15976 14282
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 15948 12850 15976 13466
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 15948 12374 15976 12650
rect 16040 12442 16068 16594
rect 16132 15094 16160 20703
rect 16316 19446 16344 22358
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16408 21962 16436 22170
rect 16396 21956 16448 21962
rect 16396 21898 16448 21904
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16224 18222 16252 18702
rect 16500 18306 16528 22918
rect 16592 22778 16620 23446
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 16684 22094 16712 25078
rect 16776 24206 16804 25434
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 16868 24954 16896 25094
rect 16856 24948 16908 24954
rect 16856 24890 16908 24896
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16868 24614 16896 24754
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16592 22066 16712 22094
rect 16868 22094 16896 24550
rect 16960 24274 16988 28358
rect 17052 26450 17080 31214
rect 17132 31136 17184 31142
rect 17132 31078 17184 31084
rect 17144 28626 17172 31078
rect 17236 30274 17264 31622
rect 17328 31482 17356 34546
rect 17420 31929 17448 35566
rect 17512 32450 17540 40326
rect 17592 37188 17644 37194
rect 17592 37130 17644 37136
rect 17604 35834 17632 37130
rect 17696 36718 17724 40666
rect 17776 39500 17828 39506
rect 17776 39442 17828 39448
rect 17788 38214 17816 39442
rect 17880 38554 17908 42230
rect 18432 41562 18460 42706
rect 18524 41682 18552 47126
rect 18616 47122 18644 51750
rect 19444 48278 19472 52838
rect 19616 52352 19668 52358
rect 19616 52294 19668 52300
rect 19432 48272 19484 48278
rect 19432 48214 19484 48220
rect 18604 47116 18656 47122
rect 18604 47058 18656 47064
rect 19340 47116 19392 47122
rect 19340 47058 19392 47064
rect 18972 46708 19024 46714
rect 18972 46650 19024 46656
rect 18604 46504 18656 46510
rect 18604 46446 18656 46452
rect 18616 44198 18644 46446
rect 18880 45280 18932 45286
rect 18880 45222 18932 45228
rect 18892 44538 18920 45222
rect 18880 44532 18932 44538
rect 18880 44474 18932 44480
rect 18604 44192 18656 44198
rect 18604 44134 18656 44140
rect 18788 44192 18840 44198
rect 18788 44134 18840 44140
rect 18512 41676 18564 41682
rect 18512 41618 18564 41624
rect 18432 41534 18552 41562
rect 18420 41472 18472 41478
rect 18420 41414 18472 41420
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 18328 40928 18380 40934
rect 18328 40870 18380 40876
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 18234 40080 18290 40089
rect 18234 40015 18290 40024
rect 18248 39914 18276 40015
rect 18236 39908 18288 39914
rect 18236 39850 18288 39856
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 18340 38826 18368 40870
rect 18432 39982 18460 41414
rect 18420 39976 18472 39982
rect 18420 39918 18472 39924
rect 18524 39642 18552 41534
rect 18696 40656 18748 40662
rect 18696 40598 18748 40604
rect 18604 40112 18656 40118
rect 18604 40054 18656 40060
rect 18512 39636 18564 39642
rect 18512 39578 18564 39584
rect 18420 39296 18472 39302
rect 18420 39238 18472 39244
rect 18432 38894 18460 39238
rect 18524 39030 18552 39578
rect 18512 39024 18564 39030
rect 18512 38966 18564 38972
rect 18420 38888 18472 38894
rect 18418 38856 18420 38865
rect 18472 38856 18474 38865
rect 18328 38820 18380 38826
rect 18418 38791 18474 38800
rect 18328 38762 18380 38768
rect 17868 38548 17920 38554
rect 17868 38490 17920 38496
rect 18340 38418 18368 38762
rect 18512 38752 18564 38758
rect 18512 38694 18564 38700
rect 18328 38412 18380 38418
rect 18328 38354 18380 38360
rect 17776 38208 17828 38214
rect 17776 38150 17828 38156
rect 17684 36712 17736 36718
rect 17684 36654 17736 36660
rect 17592 35828 17644 35834
rect 17592 35770 17644 35776
rect 17788 35766 17816 38150
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 18236 38004 18288 38010
rect 18288 37964 18368 37992
rect 18236 37946 18288 37952
rect 17868 37732 17920 37738
rect 17868 37674 17920 37680
rect 17880 37330 17908 37674
rect 17868 37324 17920 37330
rect 17868 37266 17920 37272
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 18340 35766 18368 37964
rect 18524 37210 18552 38694
rect 18616 37738 18644 40054
rect 18708 38758 18736 40598
rect 18800 39982 18828 44134
rect 18892 41206 18920 44474
rect 18984 44334 19012 46650
rect 19352 46510 19380 47058
rect 19340 46504 19392 46510
rect 19340 46446 19392 46452
rect 19444 46458 19472 48214
rect 19352 45626 19380 46446
rect 19444 46430 19564 46458
rect 19432 46368 19484 46374
rect 19432 46310 19484 46316
rect 19340 45620 19392 45626
rect 19340 45562 19392 45568
rect 19444 44962 19472 46310
rect 19536 45554 19564 46430
rect 19628 46170 19656 52294
rect 19904 52154 19932 53042
rect 20180 52494 20208 53382
rect 20168 52488 20220 52494
rect 20168 52430 20220 52436
rect 19892 52148 19944 52154
rect 19892 52090 19944 52096
rect 20272 52018 20300 56200
rect 20640 55214 20668 56200
rect 20640 55186 20760 55214
rect 20732 54194 20760 55186
rect 20720 54188 20772 54194
rect 20720 54130 20772 54136
rect 20536 54052 20588 54058
rect 20536 53994 20588 54000
rect 20548 53582 20576 53994
rect 21008 53582 21036 56200
rect 21376 54126 21404 56200
rect 21364 54120 21416 54126
rect 21364 54062 21416 54068
rect 21180 53984 21232 53990
rect 21180 53926 21232 53932
rect 20536 53576 20588 53582
rect 20536 53518 20588 53524
rect 20996 53576 21048 53582
rect 20996 53518 21048 53524
rect 20904 53440 20956 53446
rect 20904 53382 20956 53388
rect 20916 52494 20944 53382
rect 21192 52562 21220 53926
rect 21456 53576 21508 53582
rect 21456 53518 21508 53524
rect 21364 52692 21416 52698
rect 21364 52634 21416 52640
rect 21180 52556 21232 52562
rect 21180 52498 21232 52504
rect 20904 52488 20956 52494
rect 20904 52430 20956 52436
rect 20352 52352 20404 52358
rect 20352 52294 20404 52300
rect 21088 52352 21140 52358
rect 21088 52294 21140 52300
rect 20260 52012 20312 52018
rect 20260 51954 20312 51960
rect 20168 51808 20220 51814
rect 20168 51750 20220 51756
rect 19616 46164 19668 46170
rect 19616 46106 19668 46112
rect 19628 45966 19656 46106
rect 20180 46034 20208 51750
rect 20260 48000 20312 48006
rect 20260 47942 20312 47948
rect 20168 46028 20220 46034
rect 20168 45970 20220 45976
rect 19616 45960 19668 45966
rect 20076 45960 20128 45966
rect 19616 45902 19668 45908
rect 20074 45928 20076 45937
rect 20128 45928 20130 45937
rect 20074 45863 20130 45872
rect 19892 45824 19944 45830
rect 19892 45766 19944 45772
rect 19536 45526 19656 45554
rect 19444 44934 19564 44962
rect 19536 44878 19564 44934
rect 19524 44872 19576 44878
rect 19524 44814 19576 44820
rect 19536 44334 19564 44814
rect 18972 44328 19024 44334
rect 18972 44270 19024 44276
rect 19524 44328 19576 44334
rect 19524 44270 19576 44276
rect 18984 41682 19012 44270
rect 19248 43104 19300 43110
rect 19248 43046 19300 43052
rect 19260 42158 19288 43046
rect 19340 42560 19392 42566
rect 19340 42502 19392 42508
rect 19248 42152 19300 42158
rect 19248 42094 19300 42100
rect 19260 41682 19288 42094
rect 18972 41676 19024 41682
rect 18972 41618 19024 41624
rect 19248 41676 19300 41682
rect 19248 41618 19300 41624
rect 18880 41200 18932 41206
rect 18880 41142 18932 41148
rect 18788 39976 18840 39982
rect 18788 39918 18840 39924
rect 18696 38752 18748 38758
rect 18696 38694 18748 38700
rect 18696 38412 18748 38418
rect 18696 38354 18748 38360
rect 18880 38412 18932 38418
rect 18880 38354 18932 38360
rect 18708 38010 18736 38354
rect 18788 38208 18840 38214
rect 18788 38150 18840 38156
rect 18696 38004 18748 38010
rect 18696 37946 18748 37952
rect 18696 37868 18748 37874
rect 18696 37810 18748 37816
rect 18604 37732 18656 37738
rect 18604 37674 18656 37680
rect 18708 37670 18736 37810
rect 18696 37664 18748 37670
rect 18696 37606 18748 37612
rect 18524 37182 18644 37210
rect 18512 37120 18564 37126
rect 18512 37062 18564 37068
rect 18524 36922 18552 37062
rect 18512 36916 18564 36922
rect 18512 36858 18564 36864
rect 18512 36712 18564 36718
rect 18512 36654 18564 36660
rect 17776 35760 17828 35766
rect 17776 35702 17828 35708
rect 18328 35760 18380 35766
rect 18328 35702 18380 35708
rect 17960 35488 18012 35494
rect 17960 35430 18012 35436
rect 17972 35154 18000 35430
rect 18340 35290 18368 35702
rect 18328 35284 18380 35290
rect 18380 35244 18460 35272
rect 18328 35226 18380 35232
rect 17960 35148 18012 35154
rect 17960 35090 18012 35096
rect 18328 35148 18380 35154
rect 18328 35090 18380 35096
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17960 34672 18012 34678
rect 17960 34614 18012 34620
rect 17972 34202 18000 34614
rect 17960 34196 18012 34202
rect 17960 34138 18012 34144
rect 18052 34196 18104 34202
rect 18052 34138 18104 34144
rect 17868 34128 17920 34134
rect 17868 34070 17920 34076
rect 17592 33924 17644 33930
rect 17592 33866 17644 33872
rect 17604 33658 17632 33866
rect 17592 33652 17644 33658
rect 17592 33594 17644 33600
rect 17604 32842 17632 33594
rect 17592 32836 17644 32842
rect 17644 32796 17724 32824
rect 17592 32778 17644 32784
rect 17512 32422 17632 32450
rect 17500 32360 17552 32366
rect 17500 32302 17552 32308
rect 17406 31920 17462 31929
rect 17406 31855 17462 31864
rect 17420 31754 17448 31855
rect 17408 31748 17460 31754
rect 17408 31690 17460 31696
rect 17316 31476 17368 31482
rect 17316 31418 17368 31424
rect 17512 30598 17540 32302
rect 17604 32298 17632 32422
rect 17592 32292 17644 32298
rect 17592 32234 17644 32240
rect 17592 32020 17644 32026
rect 17592 31962 17644 31968
rect 17604 31210 17632 31962
rect 17592 31204 17644 31210
rect 17592 31146 17644 31152
rect 17696 30870 17724 32796
rect 17684 30864 17736 30870
rect 17684 30806 17736 30812
rect 17500 30592 17552 30598
rect 17500 30534 17552 30540
rect 17236 30246 17356 30274
rect 17224 30184 17276 30190
rect 17224 30126 17276 30132
rect 17236 29306 17264 30126
rect 17224 29300 17276 29306
rect 17224 29242 17276 29248
rect 17132 28620 17184 28626
rect 17132 28562 17184 28568
rect 17130 27432 17186 27441
rect 17130 27367 17186 27376
rect 17224 27396 17276 27402
rect 17144 27334 17172 27367
rect 17224 27338 17276 27344
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17040 26444 17092 26450
rect 17040 26386 17092 26392
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 17052 24274 17080 25094
rect 17236 24886 17264 27338
rect 17224 24880 17276 24886
rect 17224 24822 17276 24828
rect 17328 24834 17356 30246
rect 17512 30054 17540 30534
rect 17684 30116 17736 30122
rect 17684 30058 17736 30064
rect 17500 30048 17552 30054
rect 17500 29990 17552 29996
rect 17592 30048 17644 30054
rect 17592 29990 17644 29996
rect 17512 29696 17540 29990
rect 17604 29782 17632 29990
rect 17592 29776 17644 29782
rect 17592 29718 17644 29724
rect 17420 29668 17540 29696
rect 17420 29102 17448 29668
rect 17592 29572 17644 29578
rect 17592 29514 17644 29520
rect 17500 29504 17552 29510
rect 17500 29446 17552 29452
rect 17512 29306 17540 29446
rect 17604 29306 17632 29514
rect 17500 29300 17552 29306
rect 17500 29242 17552 29248
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17408 29096 17460 29102
rect 17408 29038 17460 29044
rect 17696 27470 17724 30058
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 17788 26586 17816 28562
rect 17880 28558 17908 34070
rect 18064 33930 18092 34138
rect 18052 33924 18104 33930
rect 18052 33866 18104 33872
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 18340 33590 18368 35090
rect 18432 34202 18460 35244
rect 18420 34196 18472 34202
rect 18420 34138 18472 34144
rect 18420 34060 18472 34066
rect 18420 34002 18472 34008
rect 18328 33584 18380 33590
rect 18328 33526 18380 33532
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 18432 32450 18460 34002
rect 18524 32978 18552 36654
rect 18512 32972 18564 32978
rect 18512 32914 18564 32920
rect 18616 32858 18644 37182
rect 18524 32830 18644 32858
rect 18524 32570 18552 32830
rect 18604 32768 18656 32774
rect 18604 32710 18656 32716
rect 18512 32564 18564 32570
rect 18512 32506 18564 32512
rect 18248 32422 18460 32450
rect 18248 32026 18276 32422
rect 18616 32366 18644 32710
rect 18604 32360 18656 32366
rect 18432 32320 18604 32348
rect 18328 32224 18380 32230
rect 18328 32166 18380 32172
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 18234 31784 18290 31793
rect 18234 31719 18290 31728
rect 18248 31686 18276 31719
rect 18236 31680 18288 31686
rect 18236 31622 18288 31628
rect 18340 31634 18368 32166
rect 18432 31754 18460 32320
rect 18604 32302 18656 32308
rect 18604 32020 18656 32026
rect 18604 31962 18656 31968
rect 18432 31726 18552 31754
rect 18340 31606 18460 31634
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 17960 30388 18012 30394
rect 17960 30330 18012 30336
rect 17972 30122 18000 30330
rect 18050 30288 18106 30297
rect 18050 30223 18106 30232
rect 18064 30190 18092 30223
rect 18052 30184 18104 30190
rect 18052 30126 18104 30132
rect 17960 30116 18012 30122
rect 17960 30058 18012 30064
rect 18064 29646 18092 30126
rect 18432 29696 18460 31606
rect 18248 29668 18460 29696
rect 18052 29640 18104 29646
rect 18052 29582 18104 29588
rect 18248 29510 18276 29668
rect 18524 29594 18552 31726
rect 18340 29566 18552 29594
rect 18236 29504 18288 29510
rect 18236 29446 18288 29452
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 18340 28694 18368 29566
rect 18420 29504 18472 29510
rect 18420 29446 18472 29452
rect 18512 29504 18564 29510
rect 18512 29446 18564 29452
rect 18328 28688 18380 28694
rect 18328 28630 18380 28636
rect 17868 28552 17920 28558
rect 17868 28494 17920 28500
rect 18326 28520 18382 28529
rect 18326 28455 18382 28464
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 18340 28218 18368 28455
rect 18328 28212 18380 28218
rect 18328 28154 18380 28160
rect 17868 27872 17920 27878
rect 17868 27814 17920 27820
rect 17776 26580 17828 26586
rect 17776 26522 17828 26528
rect 17880 26450 17908 27814
rect 18340 27674 18368 28154
rect 18328 27668 18380 27674
rect 18328 27610 18380 27616
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 18328 26784 18380 26790
rect 18328 26726 18380 26732
rect 17868 26444 17920 26450
rect 17868 26386 17920 26392
rect 17684 26308 17736 26314
rect 17684 26250 17736 26256
rect 17592 26240 17644 26246
rect 17592 26182 17644 26188
rect 17604 26042 17632 26182
rect 17592 26036 17644 26042
rect 17592 25978 17644 25984
rect 17604 25498 17632 25978
rect 17592 25492 17644 25498
rect 17592 25434 17644 25440
rect 17328 24806 17632 24834
rect 17696 24818 17724 26250
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 17776 25492 17828 25498
rect 17776 25434 17828 25440
rect 17604 24750 17632 24806
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17592 24744 17644 24750
rect 17592 24686 17644 24692
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 17040 24268 17092 24274
rect 17040 24210 17092 24216
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 16868 22066 16988 22094
rect 16592 19310 16620 22066
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16868 21146 16896 21286
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16960 21026 16988 22066
rect 17052 22030 17080 23598
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 17052 21078 17080 21286
rect 16868 20998 16988 21026
rect 17040 21072 17092 21078
rect 17040 21014 17092 21020
rect 16868 20806 16896 20998
rect 16948 20868 17000 20874
rect 16948 20810 17000 20816
rect 16856 20800 16908 20806
rect 16856 20742 16908 20748
rect 16868 20534 16896 20742
rect 16856 20528 16908 20534
rect 16856 20470 16908 20476
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16408 18278 16528 18306
rect 16670 18320 16726 18329
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16408 17746 16436 18278
rect 16670 18255 16726 18264
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 16120 13252 16172 13258
rect 16120 13194 16172 13200
rect 16132 12986 16160 13194
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16132 12714 16160 12922
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 15304 800 15332 2450
rect 15672 800 15700 2926
rect 15948 2650 15976 12310
rect 16224 9654 16252 17614
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16408 17066 16436 17478
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16302 16824 16358 16833
rect 16302 16759 16358 16768
rect 16316 16454 16344 16759
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16500 16096 16528 18158
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16592 17338 16620 18022
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16580 16108 16632 16114
rect 16500 16068 16580 16096
rect 16580 16050 16632 16056
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16316 11082 16344 15030
rect 16592 14498 16620 16050
rect 16684 14906 16712 18255
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16776 15026 16804 15302
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16684 14878 16804 14906
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16408 14482 16620 14498
rect 16396 14476 16620 14482
rect 16448 14470 16620 14476
rect 16396 14418 16448 14424
rect 16592 13938 16620 14470
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11694 16528 12106
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16684 4146 16712 14758
rect 16776 11830 16804 14878
rect 16868 12434 16896 16934
rect 16960 15026 16988 20810
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 17052 16182 17080 17682
rect 17144 17202 17172 24006
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 17236 21622 17264 23666
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17236 16998 17264 21354
rect 17328 21010 17356 24550
rect 17604 24410 17632 24686
rect 17592 24404 17644 24410
rect 17592 24346 17644 24352
rect 17696 24342 17724 24754
rect 17684 24336 17736 24342
rect 17684 24278 17736 24284
rect 17696 24070 17724 24278
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17684 24064 17736 24070
rect 17684 24006 17736 24012
rect 17316 21004 17368 21010
rect 17316 20946 17368 20952
rect 17314 20632 17370 20641
rect 17314 20567 17316 20576
rect 17368 20567 17370 20576
rect 17316 20538 17368 20544
rect 17316 20256 17368 20262
rect 17316 20198 17368 20204
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 17052 14618 17080 16118
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17144 14482 17172 16390
rect 17236 16182 17264 16390
rect 17328 16250 17356 20198
rect 17420 19922 17448 24006
rect 17788 23322 17816 25434
rect 17880 25158 17908 25774
rect 18340 25158 18368 26726
rect 18432 25702 18460 29446
rect 18524 29034 18552 29446
rect 18512 29028 18564 29034
rect 18512 28970 18564 28976
rect 18420 25696 18472 25702
rect 18420 25638 18472 25644
rect 17868 25152 17920 25158
rect 17868 25094 17920 25100
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 18340 24886 18368 25094
rect 18524 24886 18552 28970
rect 18616 28014 18644 31962
rect 18708 30938 18736 37606
rect 18800 36378 18828 38150
rect 18892 37942 18920 38354
rect 18880 37936 18932 37942
rect 18880 37878 18932 37884
rect 18984 37806 19012 41618
rect 19156 41472 19208 41478
rect 19156 41414 19208 41420
rect 19168 40934 19196 41414
rect 19260 41274 19288 41618
rect 19248 41268 19300 41274
rect 19248 41210 19300 41216
rect 19156 40928 19208 40934
rect 19156 40870 19208 40876
rect 19168 40458 19196 40870
rect 19352 40526 19380 42502
rect 19524 42220 19576 42226
rect 19524 42162 19576 42168
rect 19432 40928 19484 40934
rect 19432 40870 19484 40876
rect 19340 40520 19392 40526
rect 19340 40462 19392 40468
rect 19156 40452 19208 40458
rect 19156 40394 19208 40400
rect 19064 39840 19116 39846
rect 19064 39782 19116 39788
rect 19076 39642 19104 39782
rect 19064 39636 19116 39642
rect 19064 39578 19116 39584
rect 19076 38350 19104 39578
rect 19168 39114 19196 40394
rect 19444 39506 19472 40870
rect 19536 39914 19564 42162
rect 19524 39908 19576 39914
rect 19524 39850 19576 39856
rect 19628 39642 19656 45526
rect 19800 44804 19852 44810
rect 19800 44746 19852 44752
rect 19812 44538 19840 44746
rect 19800 44532 19852 44538
rect 19800 44474 19852 44480
rect 19800 42356 19852 42362
rect 19800 42298 19852 42304
rect 19708 42152 19760 42158
rect 19708 42094 19760 42100
rect 19720 41546 19748 42094
rect 19708 41540 19760 41546
rect 19708 41482 19760 41488
rect 19616 39636 19668 39642
rect 19616 39578 19668 39584
rect 19614 39536 19670 39545
rect 19432 39500 19484 39506
rect 19614 39471 19670 39480
rect 19432 39442 19484 39448
rect 19168 39086 19288 39114
rect 19156 38888 19208 38894
rect 19156 38830 19208 38836
rect 19064 38344 19116 38350
rect 19064 38286 19116 38292
rect 18972 37800 19024 37806
rect 18972 37742 19024 37748
rect 19076 37738 19104 38286
rect 19064 37732 19116 37738
rect 19064 37674 19116 37680
rect 18972 37664 19024 37670
rect 18972 37606 19024 37612
rect 18788 36372 18840 36378
rect 18788 36314 18840 36320
rect 18788 34196 18840 34202
rect 18788 34138 18840 34144
rect 18800 33590 18828 34138
rect 18788 33584 18840 33590
rect 18788 33526 18840 33532
rect 18788 31952 18840 31958
rect 18788 31894 18840 31900
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18694 30288 18750 30297
rect 18694 30223 18696 30232
rect 18748 30223 18750 30232
rect 18696 30194 18748 30200
rect 18696 30116 18748 30122
rect 18696 30058 18748 30064
rect 18604 28008 18656 28014
rect 18604 27950 18656 27956
rect 18604 27668 18656 27674
rect 18604 27610 18656 27616
rect 18328 24880 18380 24886
rect 18328 24822 18380 24828
rect 18512 24880 18564 24886
rect 18512 24822 18564 24828
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17880 23798 17908 24754
rect 18616 24698 18644 27610
rect 18432 24670 18644 24698
rect 18708 24682 18736 30058
rect 18800 28762 18828 31894
rect 18880 31748 18932 31754
rect 18880 31690 18932 31696
rect 18892 31278 18920 31690
rect 18880 31272 18932 31278
rect 18880 31214 18932 31220
rect 18880 30388 18932 30394
rect 18880 30330 18932 30336
rect 18892 29238 18920 30330
rect 18984 29850 19012 37606
rect 19168 35562 19196 38830
rect 19260 38400 19288 39086
rect 19260 38372 19472 38400
rect 19248 38276 19300 38282
rect 19248 38218 19300 38224
rect 19340 38276 19392 38282
rect 19340 38218 19392 38224
rect 19260 36378 19288 38218
rect 19248 36372 19300 36378
rect 19248 36314 19300 36320
rect 19156 35556 19208 35562
rect 19156 35498 19208 35504
rect 19168 33862 19196 35498
rect 19156 33856 19208 33862
rect 19156 33798 19208 33804
rect 19156 31680 19208 31686
rect 19156 31622 19208 31628
rect 19168 31142 19196 31622
rect 19248 31340 19300 31346
rect 19248 31282 19300 31288
rect 19156 31136 19208 31142
rect 19156 31078 19208 31084
rect 19064 30796 19116 30802
rect 19064 30738 19116 30744
rect 18972 29844 19024 29850
rect 18972 29786 19024 29792
rect 19076 29714 19104 30738
rect 19064 29708 19116 29714
rect 19064 29650 19116 29656
rect 18972 29640 19024 29646
rect 18972 29582 19024 29588
rect 18880 29232 18932 29238
rect 18880 29174 18932 29180
rect 18984 29050 19012 29582
rect 18892 29022 19012 29050
rect 18788 28756 18840 28762
rect 18788 28698 18840 28704
rect 18788 28008 18840 28014
rect 18788 27950 18840 27956
rect 18800 24750 18828 27950
rect 18892 25786 18920 29022
rect 18972 28756 19024 28762
rect 18972 28698 19024 28704
rect 18984 27062 19012 28698
rect 19076 28218 19104 29650
rect 19064 28212 19116 28218
rect 19064 28154 19116 28160
rect 19064 27872 19116 27878
rect 19064 27814 19116 27820
rect 18972 27056 19024 27062
rect 18972 26998 19024 27004
rect 18892 25758 19012 25786
rect 18880 25696 18932 25702
rect 18880 25638 18932 25644
rect 18788 24744 18840 24750
rect 18788 24686 18840 24692
rect 18696 24676 18748 24682
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 17776 23316 17828 23322
rect 17776 23258 17828 23264
rect 17788 23050 17816 23258
rect 17776 23044 17828 23050
rect 17776 22986 17828 22992
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 17512 18290 17540 22714
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17684 21616 17736 21622
rect 17684 21558 17736 21564
rect 17592 21480 17644 21486
rect 17592 21422 17644 21428
rect 17604 20942 17632 21422
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17604 19378 17632 19722
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17512 18086 17540 18226
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17236 14278 17264 16118
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17236 14074 17264 14214
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 16868 12406 16988 12434
rect 16960 12238 16988 12406
rect 17144 12306 17172 13874
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17236 12986 17264 13126
rect 17328 12986 17356 15098
rect 17420 14006 17448 15506
rect 17696 15502 17724 21558
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17960 20528 18012 20534
rect 17960 20470 18012 20476
rect 17868 20324 17920 20330
rect 17868 20266 17920 20272
rect 17774 19952 17830 19961
rect 17774 19887 17830 19896
rect 17788 19854 17816 19887
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17788 18834 17816 19246
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17880 14958 17908 20266
rect 17972 19990 18000 20470
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18340 18970 18368 22578
rect 18432 21434 18460 24670
rect 18696 24618 18748 24624
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18524 22098 18552 24550
rect 18708 24342 18736 24618
rect 18696 24336 18748 24342
rect 18696 24278 18748 24284
rect 18800 24138 18828 24686
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18616 23186 18644 23598
rect 18604 23180 18656 23186
rect 18604 23122 18656 23128
rect 18616 22710 18644 23122
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 18800 22522 18828 24074
rect 18616 22494 18828 22522
rect 18616 22234 18644 22494
rect 18788 22432 18840 22438
rect 18788 22374 18840 22380
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18512 22092 18564 22098
rect 18512 22034 18564 22040
rect 18432 21406 18552 21434
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18524 21298 18552 21406
rect 18432 19938 18460 21286
rect 18524 21270 18644 21298
rect 18510 20632 18566 20641
rect 18510 20567 18566 20576
rect 18524 20466 18552 20567
rect 18616 20534 18644 21270
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18800 20346 18828 22374
rect 18616 20318 18828 20346
rect 18432 19910 18552 19938
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 18432 19417 18460 19722
rect 18418 19408 18474 19417
rect 18418 19343 18474 19352
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18326 18728 18382 18737
rect 18326 18663 18382 18672
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18340 18426 18368 18663
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17972 16454 18000 17206
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17408 14000 17460 14006
rect 17460 13948 17540 13954
rect 17408 13942 17540 13948
rect 17420 13926 17540 13942
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16132 3670 16160 4082
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16040 800 16068 3538
rect 16408 800 16436 4014
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16776 800 16804 2790
rect 16868 2446 16896 9862
rect 16960 7478 16988 12174
rect 17420 12102 17448 13806
rect 17512 12442 17540 13926
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 17052 3058 17080 11494
rect 17604 9602 17632 14826
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17880 13734 17908 13942
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18340 12986 18368 18362
rect 18432 14074 18460 18566
rect 18524 18154 18552 19910
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 18616 17218 18644 20318
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18524 17190 18644 17218
rect 18524 14414 18552 17190
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18616 16250 18644 17070
rect 18708 16726 18736 19450
rect 18696 16720 18748 16726
rect 18696 16662 18748 16668
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18708 16250 18736 16390
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18616 15026 18644 16186
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18708 15162 18736 15302
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18800 15042 18828 20198
rect 18892 19854 18920 25638
rect 18984 23798 19012 25758
rect 19076 25362 19104 27814
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 18972 23792 19024 23798
rect 18972 23734 19024 23740
rect 18984 22438 19012 23734
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 19076 22574 19104 23598
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 19168 22094 19196 31078
rect 19260 24750 19288 31282
rect 19352 29578 19380 38218
rect 19444 37670 19472 38372
rect 19432 37664 19484 37670
rect 19432 37606 19484 37612
rect 19432 37188 19484 37194
rect 19432 37130 19484 37136
rect 19444 36650 19472 37130
rect 19432 36644 19484 36650
rect 19432 36586 19484 36592
rect 19628 36122 19656 39471
rect 19720 36242 19748 41482
rect 19812 36786 19840 42298
rect 19904 41274 19932 45766
rect 20272 45554 20300 47942
rect 20364 47258 20392 52294
rect 20996 49972 21048 49978
rect 20996 49914 21048 49920
rect 20352 47252 20404 47258
rect 20352 47194 20404 47200
rect 20904 46640 20956 46646
rect 20904 46582 20956 46588
rect 20444 46028 20496 46034
rect 20444 45970 20496 45976
rect 20180 45526 20300 45554
rect 20076 45416 20128 45422
rect 20076 45358 20128 45364
rect 19984 44736 20036 44742
rect 19984 44678 20036 44684
rect 19996 43246 20024 44678
rect 20088 43450 20116 45358
rect 20076 43444 20128 43450
rect 20076 43386 20128 43392
rect 19984 43240 20036 43246
rect 19984 43182 20036 43188
rect 19892 41268 19944 41274
rect 19892 41210 19944 41216
rect 19996 41070 20024 43182
rect 19984 41064 20036 41070
rect 19984 41006 20036 41012
rect 19996 40730 20024 41006
rect 19984 40724 20036 40730
rect 19984 40666 20036 40672
rect 19984 40520 20036 40526
rect 19984 40462 20036 40468
rect 19996 40361 20024 40462
rect 19982 40352 20038 40361
rect 19982 40287 20038 40296
rect 19892 39296 19944 39302
rect 19892 39238 19944 39244
rect 19800 36780 19852 36786
rect 19800 36722 19852 36728
rect 19708 36236 19760 36242
rect 19708 36178 19760 36184
rect 19628 36094 19748 36122
rect 19616 36032 19668 36038
rect 19616 35974 19668 35980
rect 19524 34468 19576 34474
rect 19524 34410 19576 34416
rect 19432 31952 19484 31958
rect 19430 31920 19432 31929
rect 19484 31920 19486 31929
rect 19430 31855 19486 31864
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19340 29572 19392 29578
rect 19340 29514 19392 29520
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 19352 27334 19380 28018
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19340 26920 19392 26926
rect 19340 26862 19392 26868
rect 19352 26042 19380 26862
rect 19340 26036 19392 26042
rect 19340 25978 19392 25984
rect 19444 25294 19472 30534
rect 19536 30190 19564 34410
rect 19628 30938 19656 35974
rect 19720 35290 19748 36094
rect 19800 35488 19852 35494
rect 19904 35465 19932 39238
rect 19996 35766 20024 40287
rect 20088 39506 20116 43386
rect 20180 42362 20208 45526
rect 20456 44538 20484 45970
rect 20720 45824 20772 45830
rect 20720 45766 20772 45772
rect 20444 44532 20496 44538
rect 20444 44474 20496 44480
rect 20260 43648 20312 43654
rect 20260 43590 20312 43596
rect 20168 42356 20220 42362
rect 20168 42298 20220 42304
rect 20272 40050 20300 43590
rect 20352 42900 20404 42906
rect 20352 42842 20404 42848
rect 20260 40044 20312 40050
rect 20260 39986 20312 39992
rect 20272 39846 20300 39986
rect 20364 39930 20392 42842
rect 20536 42560 20588 42566
rect 20536 42502 20588 42508
rect 20548 42158 20576 42502
rect 20732 42362 20760 45766
rect 20916 45286 20944 46582
rect 20904 45280 20956 45286
rect 20904 45222 20956 45228
rect 20916 44878 20944 45222
rect 20904 44872 20956 44878
rect 20904 44814 20956 44820
rect 20812 44328 20864 44334
rect 20812 44270 20864 44276
rect 20720 42356 20772 42362
rect 20720 42298 20772 42304
rect 20536 42152 20588 42158
rect 20536 42094 20588 42100
rect 20720 42016 20772 42022
rect 20720 41958 20772 41964
rect 20444 41132 20496 41138
rect 20444 41074 20496 41080
rect 20456 40390 20484 41074
rect 20444 40384 20496 40390
rect 20444 40326 20496 40332
rect 20456 40089 20484 40326
rect 20442 40080 20498 40089
rect 20442 40015 20498 40024
rect 20444 39976 20496 39982
rect 20364 39924 20444 39930
rect 20364 39918 20496 39924
rect 20536 39976 20588 39982
rect 20536 39918 20588 39924
rect 20364 39902 20484 39918
rect 20260 39840 20312 39846
rect 20260 39782 20312 39788
rect 20272 39545 20300 39782
rect 20444 39636 20496 39642
rect 20444 39578 20496 39584
rect 20258 39536 20314 39545
rect 20076 39500 20128 39506
rect 20258 39471 20314 39480
rect 20076 39442 20128 39448
rect 20260 39432 20312 39438
rect 20260 39374 20312 39380
rect 20272 38026 20300 39374
rect 20456 38894 20484 39578
rect 20444 38888 20496 38894
rect 20444 38830 20496 38836
rect 20352 38752 20404 38758
rect 20352 38694 20404 38700
rect 20444 38752 20496 38758
rect 20444 38694 20496 38700
rect 20180 37998 20300 38026
rect 20180 37670 20208 37998
rect 20258 37904 20314 37913
rect 20258 37839 20260 37848
rect 20312 37839 20314 37848
rect 20260 37810 20312 37816
rect 20168 37664 20220 37670
rect 20168 37606 20220 37612
rect 20260 37324 20312 37330
rect 20260 37266 20312 37272
rect 20168 37188 20220 37194
rect 20168 37130 20220 37136
rect 20076 37120 20128 37126
rect 20076 37062 20128 37068
rect 20088 36582 20116 37062
rect 20076 36576 20128 36582
rect 20076 36518 20128 36524
rect 19984 35760 20036 35766
rect 19984 35702 20036 35708
rect 19800 35430 19852 35436
rect 19890 35456 19946 35465
rect 19708 35284 19760 35290
rect 19708 35226 19760 35232
rect 19708 35012 19760 35018
rect 19708 34954 19760 34960
rect 19720 34678 19748 34954
rect 19812 34746 19840 35430
rect 19890 35391 19946 35400
rect 19892 34944 19944 34950
rect 19892 34886 19944 34892
rect 19800 34740 19852 34746
rect 19800 34682 19852 34688
rect 19708 34672 19760 34678
rect 19708 34614 19760 34620
rect 19904 33658 19932 34886
rect 20088 33998 20116 36518
rect 20180 35154 20208 37130
rect 20168 35148 20220 35154
rect 20168 35090 20220 35096
rect 20272 34746 20300 37266
rect 20364 36242 20392 38694
rect 20456 38350 20484 38694
rect 20444 38344 20496 38350
rect 20444 38286 20496 38292
rect 20456 36922 20484 38286
rect 20548 37806 20576 39918
rect 20628 38344 20680 38350
rect 20628 38286 20680 38292
rect 20640 38010 20668 38286
rect 20628 38004 20680 38010
rect 20628 37946 20680 37952
rect 20536 37800 20588 37806
rect 20536 37742 20588 37748
rect 20640 37652 20668 37946
rect 20548 37624 20668 37652
rect 20548 37398 20576 37624
rect 20536 37392 20588 37398
rect 20536 37334 20588 37340
rect 20444 36916 20496 36922
rect 20444 36858 20496 36864
rect 20444 36644 20496 36650
rect 20444 36586 20496 36592
rect 20352 36236 20404 36242
rect 20352 36178 20404 36184
rect 20352 35284 20404 35290
rect 20352 35226 20404 35232
rect 20260 34740 20312 34746
rect 20260 34682 20312 34688
rect 20168 34400 20220 34406
rect 20168 34342 20220 34348
rect 20076 33992 20128 33998
rect 20076 33934 20128 33940
rect 20180 33674 20208 34342
rect 20272 33930 20300 34682
rect 20260 33924 20312 33930
rect 20260 33866 20312 33872
rect 19892 33652 19944 33658
rect 19892 33594 19944 33600
rect 20088 33646 20208 33674
rect 19904 31958 19932 33594
rect 19982 32056 20038 32065
rect 19982 31991 20038 32000
rect 19892 31952 19944 31958
rect 19892 31894 19944 31900
rect 19996 31754 20024 31991
rect 19812 31726 20024 31754
rect 19616 30932 19668 30938
rect 19616 30874 19668 30880
rect 19524 30184 19576 30190
rect 19524 30126 19576 30132
rect 19536 28472 19564 30126
rect 19812 29850 19840 31726
rect 19984 31272 20036 31278
rect 19982 31240 19984 31249
rect 20036 31240 20038 31249
rect 19982 31175 20038 31184
rect 19890 30832 19946 30841
rect 19890 30767 19892 30776
rect 19944 30767 19946 30776
rect 19984 30796 20036 30802
rect 19892 30738 19944 30744
rect 19984 30738 20036 30744
rect 19800 29844 19852 29850
rect 19800 29786 19852 29792
rect 19812 29306 19840 29786
rect 19800 29300 19852 29306
rect 19800 29242 19852 29248
rect 19616 28484 19668 28490
rect 19536 28444 19616 28472
rect 19536 26926 19564 28444
rect 19616 28426 19668 28432
rect 19996 28014 20024 30738
rect 20088 30734 20116 33646
rect 20260 33584 20312 33590
rect 20258 33552 20260 33561
rect 20312 33552 20314 33561
rect 20258 33487 20314 33496
rect 20168 32428 20220 32434
rect 20168 32370 20220 32376
rect 20180 32337 20208 32370
rect 20166 32328 20222 32337
rect 20166 32263 20222 32272
rect 20260 31952 20312 31958
rect 20260 31894 20312 31900
rect 20168 31136 20220 31142
rect 20168 31078 20220 31084
rect 20076 30728 20128 30734
rect 20076 30670 20128 30676
rect 20180 30580 20208 31078
rect 20088 30552 20208 30580
rect 20088 29238 20116 30552
rect 20168 29300 20220 29306
rect 20168 29242 20220 29248
rect 20076 29232 20128 29238
rect 20076 29174 20128 29180
rect 20088 28948 20116 29174
rect 20180 29102 20208 29242
rect 20168 29096 20220 29102
rect 20166 29064 20168 29073
rect 20220 29064 20222 29073
rect 20166 28999 20222 29008
rect 20088 28920 20208 28948
rect 20074 28384 20130 28393
rect 20074 28319 20130 28328
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19524 26920 19576 26926
rect 19524 26862 19576 26868
rect 19524 26784 19576 26790
rect 19524 26726 19576 26732
rect 19536 26042 19564 26726
rect 19708 26512 19760 26518
rect 19708 26454 19760 26460
rect 19524 26036 19576 26042
rect 19524 25978 19576 25984
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19524 25152 19576 25158
rect 19524 25094 19576 25100
rect 19248 24744 19300 24750
rect 19248 24686 19300 24692
rect 19248 24132 19300 24138
rect 19248 24074 19300 24080
rect 19260 23866 19288 24074
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 19352 23322 19380 23734
rect 19444 23662 19472 24006
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 19352 22982 19380 23258
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 18984 22066 19196 22094
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18984 18970 19012 22066
rect 19156 20868 19208 20874
rect 19156 20810 19208 20816
rect 19168 20777 19196 20810
rect 19154 20768 19210 20777
rect 19154 20703 19210 20712
rect 19064 19712 19116 19718
rect 19064 19654 19116 19660
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 18984 18766 19012 18906
rect 19076 18902 19104 19654
rect 19260 19446 19288 22374
rect 19352 22030 19380 22578
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 19352 20602 19380 21014
rect 19444 21010 19472 21966
rect 19432 21004 19484 21010
rect 19432 20946 19484 20952
rect 19536 20602 19564 25094
rect 19720 22710 19748 26454
rect 19892 24812 19944 24818
rect 19892 24754 19944 24760
rect 19904 24614 19932 24754
rect 19892 24608 19944 24614
rect 19892 24550 19944 24556
rect 19708 22704 19760 22710
rect 19708 22646 19760 22652
rect 19904 22094 19932 24550
rect 19996 23050 20024 27950
rect 20088 27878 20116 28319
rect 20076 27872 20128 27878
rect 20074 27840 20076 27849
rect 20128 27840 20130 27849
rect 20074 27775 20130 27784
rect 20180 27130 20208 28920
rect 20168 27124 20220 27130
rect 20168 27066 20220 27072
rect 20168 26444 20220 26450
rect 20168 26386 20220 26392
rect 20076 25356 20128 25362
rect 20076 25298 20128 25304
rect 20088 23322 20116 25298
rect 20180 24052 20208 26386
rect 20272 26382 20300 31894
rect 20364 31142 20392 35226
rect 20456 33454 20484 36586
rect 20444 33448 20496 33454
rect 20444 33390 20496 33396
rect 20548 32065 20576 37334
rect 20732 37262 20760 41958
rect 20824 41818 20852 44270
rect 20812 41812 20864 41818
rect 20812 41754 20864 41760
rect 20904 41132 20956 41138
rect 20904 41074 20956 41080
rect 20916 40934 20944 41074
rect 21008 41070 21036 49914
rect 21100 45966 21128 52294
rect 21376 46034 21404 52634
rect 21468 52154 21496 53518
rect 21640 52964 21692 52970
rect 21640 52906 21692 52912
rect 21548 52624 21600 52630
rect 21548 52566 21600 52572
rect 21456 52148 21508 52154
rect 21456 52090 21508 52096
rect 21364 46028 21416 46034
rect 21364 45970 21416 45976
rect 21088 45960 21140 45966
rect 21088 45902 21140 45908
rect 21364 43444 21416 43450
rect 21364 43386 21416 43392
rect 21376 42702 21404 43386
rect 21560 43330 21588 52566
rect 21652 47258 21680 52906
rect 21744 52562 21772 56200
rect 22112 55214 22140 56200
rect 22112 55186 22232 55214
rect 22100 53984 22152 53990
rect 22100 53926 22152 53932
rect 22008 53440 22060 53446
rect 22008 53382 22060 53388
rect 22020 53106 22048 53382
rect 22008 53100 22060 53106
rect 22008 53042 22060 53048
rect 21732 52556 21784 52562
rect 21732 52498 21784 52504
rect 22112 52494 22140 53926
rect 22204 53514 22232 55186
rect 22480 53650 22508 56200
rect 22652 53712 22704 53718
rect 22652 53654 22704 53660
rect 22468 53644 22520 53650
rect 22468 53586 22520 53592
rect 22192 53508 22244 53514
rect 22192 53450 22244 53456
rect 22560 52896 22612 52902
rect 22560 52838 22612 52844
rect 22468 52624 22520 52630
rect 22468 52566 22520 52572
rect 22100 52488 22152 52494
rect 22100 52430 22152 52436
rect 22376 51808 22428 51814
rect 22376 51750 22428 51756
rect 21640 47252 21692 47258
rect 21640 47194 21692 47200
rect 21652 47054 21680 47194
rect 21824 47184 21876 47190
rect 21824 47126 21876 47132
rect 21640 47048 21692 47054
rect 21638 47016 21640 47025
rect 21692 47016 21694 47025
rect 21638 46951 21694 46960
rect 21732 46028 21784 46034
rect 21732 45970 21784 45976
rect 21744 45558 21772 45970
rect 21732 45552 21784 45558
rect 21732 45494 21784 45500
rect 21640 44940 21692 44946
rect 21640 44882 21692 44888
rect 21652 44538 21680 44882
rect 21640 44532 21692 44538
rect 21640 44474 21692 44480
rect 21652 43450 21680 44474
rect 21640 43444 21692 43450
rect 21640 43386 21692 43392
rect 21560 43314 21680 43330
rect 21560 43308 21692 43314
rect 21560 43302 21640 43308
rect 21640 43250 21692 43256
rect 21652 43110 21680 43250
rect 21640 43104 21692 43110
rect 21638 43072 21640 43081
rect 21692 43072 21694 43081
rect 21638 43007 21694 43016
rect 21744 42906 21772 45494
rect 21732 42900 21784 42906
rect 21732 42842 21784 42848
rect 21364 42696 21416 42702
rect 21364 42638 21416 42644
rect 21180 42628 21232 42634
rect 21180 42570 21232 42576
rect 21088 42288 21140 42294
rect 21088 42230 21140 42236
rect 20996 41064 21048 41070
rect 20996 41006 21048 41012
rect 20812 40928 20864 40934
rect 20812 40870 20864 40876
rect 20904 40928 20956 40934
rect 20904 40870 20956 40876
rect 20824 39030 20852 40870
rect 20812 39024 20864 39030
rect 20812 38966 20864 38972
rect 20812 38480 20864 38486
rect 20812 38422 20864 38428
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 20824 37194 20852 38422
rect 20812 37188 20864 37194
rect 20812 37130 20864 37136
rect 20916 36174 20944 40870
rect 21008 39098 21036 41006
rect 20996 39092 21048 39098
rect 20996 39034 21048 39040
rect 20996 38888 21048 38894
rect 20996 38830 21048 38836
rect 20904 36168 20956 36174
rect 20904 36110 20956 36116
rect 20904 36032 20956 36038
rect 20904 35974 20956 35980
rect 20720 35488 20772 35494
rect 20720 35430 20772 35436
rect 20732 35222 20760 35430
rect 20720 35216 20772 35222
rect 20720 35158 20772 35164
rect 20732 35018 20760 35158
rect 20720 35012 20772 35018
rect 20720 34954 20772 34960
rect 20732 34202 20760 34954
rect 20812 34740 20864 34746
rect 20812 34682 20864 34688
rect 20720 34196 20772 34202
rect 20720 34138 20772 34144
rect 20628 33856 20680 33862
rect 20628 33798 20680 33804
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20640 33522 20668 33798
rect 20628 33516 20680 33522
rect 20628 33458 20680 33464
rect 20640 32842 20668 33458
rect 20628 32836 20680 32842
rect 20628 32778 20680 32784
rect 20628 32224 20680 32230
rect 20628 32166 20680 32172
rect 20534 32056 20590 32065
rect 20534 31991 20590 32000
rect 20640 31414 20668 32166
rect 20732 31754 20760 33798
rect 20720 31748 20772 31754
rect 20720 31690 20772 31696
rect 20628 31408 20680 31414
rect 20628 31350 20680 31356
rect 20444 31204 20496 31210
rect 20444 31146 20496 31152
rect 20352 31136 20404 31142
rect 20352 31078 20404 31084
rect 20352 30932 20404 30938
rect 20352 30874 20404 30880
rect 20364 29594 20392 30874
rect 20456 30734 20484 31146
rect 20628 31136 20680 31142
rect 20628 31078 20680 31084
rect 20536 30796 20588 30802
rect 20536 30738 20588 30744
rect 20444 30728 20496 30734
rect 20444 30670 20496 30676
rect 20364 29566 20484 29594
rect 20352 29504 20404 29510
rect 20352 29446 20404 29452
rect 20260 26376 20312 26382
rect 20260 26318 20312 26324
rect 20364 26042 20392 29446
rect 20456 27538 20484 29566
rect 20548 29238 20576 30738
rect 20536 29232 20588 29238
rect 20536 29174 20588 29180
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 20444 27124 20496 27130
rect 20444 27066 20496 27072
rect 20352 26036 20404 26042
rect 20352 25978 20404 25984
rect 20260 24064 20312 24070
rect 20180 24024 20260 24052
rect 20260 24006 20312 24012
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 20272 22234 20300 24006
rect 20456 23610 20484 27066
rect 20548 24682 20576 29174
rect 20640 27538 20668 31078
rect 20824 29646 20852 34682
rect 20916 31822 20944 35974
rect 21008 34950 21036 38830
rect 21100 38418 21128 42230
rect 21192 40730 21220 42570
rect 21376 42362 21404 42638
rect 21364 42356 21416 42362
rect 21364 42298 21416 42304
rect 21272 41812 21324 41818
rect 21272 41754 21324 41760
rect 21180 40724 21232 40730
rect 21180 40666 21232 40672
rect 21180 40520 21232 40526
rect 21180 40462 21232 40468
rect 21192 40118 21220 40462
rect 21180 40112 21232 40118
rect 21180 40054 21232 40060
rect 21284 38418 21312 41754
rect 21376 41546 21404 42298
rect 21732 41812 21784 41818
rect 21732 41754 21784 41760
rect 21364 41540 21416 41546
rect 21364 41482 21416 41488
rect 21548 41540 21600 41546
rect 21548 41482 21600 41488
rect 21560 41414 21588 41482
rect 21640 41472 21692 41478
rect 21640 41414 21692 41420
rect 21468 41386 21588 41414
rect 21364 40044 21416 40050
rect 21364 39986 21416 39992
rect 21376 39953 21404 39986
rect 21362 39944 21418 39953
rect 21362 39879 21418 39888
rect 21364 38956 21416 38962
rect 21364 38898 21416 38904
rect 21088 38412 21140 38418
rect 21088 38354 21140 38360
rect 21272 38412 21324 38418
rect 21272 38354 21324 38360
rect 21088 38208 21140 38214
rect 21088 38150 21140 38156
rect 20996 34944 21048 34950
rect 20996 34886 21048 34892
rect 21100 32570 21128 38150
rect 21180 37188 21232 37194
rect 21180 37130 21232 37136
rect 21192 34746 21220 37130
rect 21376 36394 21404 38898
rect 21468 37942 21496 41386
rect 21548 40588 21600 40594
rect 21548 40530 21600 40536
rect 21560 40458 21588 40530
rect 21652 40526 21680 41414
rect 21744 40594 21772 41754
rect 21732 40588 21784 40594
rect 21732 40530 21784 40536
rect 21640 40520 21692 40526
rect 21640 40462 21692 40468
rect 21548 40452 21600 40458
rect 21548 40394 21600 40400
rect 21560 39982 21588 40394
rect 21744 40390 21772 40530
rect 21732 40384 21784 40390
rect 21732 40326 21784 40332
rect 21744 40050 21772 40326
rect 21732 40044 21784 40050
rect 21732 39986 21784 39992
rect 21548 39976 21600 39982
rect 21548 39918 21600 39924
rect 21548 39500 21600 39506
rect 21548 39442 21600 39448
rect 21560 38010 21588 39442
rect 21744 39370 21772 39986
rect 21836 39914 21864 47126
rect 22008 46912 22060 46918
rect 22008 46854 22060 46860
rect 21916 45960 21968 45966
rect 21914 45928 21916 45937
rect 21968 45928 21970 45937
rect 21914 45863 21970 45872
rect 21916 43648 21968 43654
rect 21916 43590 21968 43596
rect 21824 39908 21876 39914
rect 21824 39850 21876 39856
rect 21732 39364 21784 39370
rect 21732 39306 21784 39312
rect 21928 38418 21956 43590
rect 22020 42770 22048 46854
rect 22192 46504 22244 46510
rect 22192 46446 22244 46452
rect 22204 44554 22232 46446
rect 22284 45280 22336 45286
rect 22284 45222 22336 45228
rect 22296 44878 22324 45222
rect 22284 44872 22336 44878
rect 22284 44814 22336 44820
rect 22112 44526 22232 44554
rect 22112 43194 22140 44526
rect 22296 44334 22324 44814
rect 22284 44328 22336 44334
rect 22284 44270 22336 44276
rect 22388 43450 22416 51750
rect 22480 43858 22508 52566
rect 22572 46714 22600 52838
rect 22664 47054 22692 53654
rect 22744 52964 22796 52970
rect 22744 52906 22796 52912
rect 22756 52494 22784 52906
rect 22744 52488 22796 52494
rect 22744 52430 22796 52436
rect 22848 52018 22876 56200
rect 23216 55214 23244 56200
rect 23216 55186 23336 55214
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 23308 52494 23336 55186
rect 23480 53440 23532 53446
rect 23480 53382 23532 53388
rect 23492 53106 23520 53382
rect 23480 53100 23532 53106
rect 23480 53042 23532 53048
rect 22928 52488 22980 52494
rect 22928 52430 22980 52436
rect 23296 52488 23348 52494
rect 23296 52430 23348 52436
rect 22836 52012 22888 52018
rect 22836 51954 22888 51960
rect 22940 51898 22968 52430
rect 23584 52034 23612 56200
rect 24582 56199 24638 56208
rect 24032 54188 24084 54194
rect 24032 54130 24084 54136
rect 23756 53984 23808 53990
rect 23756 53926 23808 53932
rect 23848 53984 23900 53990
rect 23848 53926 23900 53932
rect 23768 53174 23796 53926
rect 23756 53168 23808 53174
rect 23756 53110 23808 53116
rect 23664 52896 23716 52902
rect 23664 52838 23716 52844
rect 23676 52601 23704 52838
rect 23662 52592 23718 52601
rect 23662 52527 23718 52536
rect 23584 52018 23704 52034
rect 23584 52012 23716 52018
rect 23584 52006 23664 52012
rect 23664 51954 23716 51960
rect 22744 51876 22796 51882
rect 22744 51818 22796 51824
rect 22848 51870 22968 51898
rect 22652 47048 22704 47054
rect 22652 46990 22704 46996
rect 22652 46912 22704 46918
rect 22652 46854 22704 46860
rect 22560 46708 22612 46714
rect 22560 46650 22612 46656
rect 22572 46617 22600 46650
rect 22558 46608 22614 46617
rect 22558 46543 22614 46552
rect 22560 44804 22612 44810
rect 22560 44746 22612 44752
rect 22572 44538 22600 44746
rect 22560 44532 22612 44538
rect 22560 44474 22612 44480
rect 22468 43852 22520 43858
rect 22468 43794 22520 43800
rect 22468 43648 22520 43654
rect 22468 43590 22520 43596
rect 22376 43444 22428 43450
rect 22376 43386 22428 43392
rect 22374 43344 22430 43353
rect 22374 43279 22430 43288
rect 22112 43166 22232 43194
rect 22008 42764 22060 42770
rect 22008 42706 22060 42712
rect 22100 42560 22152 42566
rect 22100 42502 22152 42508
rect 22008 41472 22060 41478
rect 22008 41414 22060 41420
rect 22020 41274 22048 41414
rect 22008 41268 22060 41274
rect 22008 41210 22060 41216
rect 22112 40594 22140 42502
rect 22204 41002 22232 43166
rect 22284 41540 22336 41546
rect 22284 41482 22336 41488
rect 22192 40996 22244 41002
rect 22192 40938 22244 40944
rect 22100 40588 22152 40594
rect 22100 40530 22152 40536
rect 22100 40180 22152 40186
rect 22100 40122 22152 40128
rect 22112 39250 22140 40122
rect 22204 39506 22232 40938
rect 22296 39642 22324 41482
rect 22388 40458 22416 43279
rect 22480 41414 22508 43590
rect 22572 42770 22600 44474
rect 22664 44334 22692 46854
rect 22756 46714 22784 51818
rect 22744 46708 22796 46714
rect 22744 46650 22796 46656
rect 22744 46368 22796 46374
rect 22744 46310 22796 46316
rect 22652 44328 22704 44334
rect 22652 44270 22704 44276
rect 22664 43353 22692 44270
rect 22650 43344 22706 43353
rect 22650 43279 22706 43288
rect 22652 43240 22704 43246
rect 22652 43182 22704 43188
rect 22560 42764 22612 42770
rect 22560 42706 22612 42712
rect 22572 41682 22600 42706
rect 22560 41676 22612 41682
rect 22560 41618 22612 41624
rect 22480 41386 22600 41414
rect 22468 41064 22520 41070
rect 22468 41006 22520 41012
rect 22376 40452 22428 40458
rect 22376 40394 22428 40400
rect 22480 40202 22508 41006
rect 22388 40174 22508 40202
rect 22284 39636 22336 39642
rect 22284 39578 22336 39584
rect 22192 39500 22244 39506
rect 22192 39442 22244 39448
rect 22112 39222 22232 39250
rect 22100 39092 22152 39098
rect 22100 39034 22152 39040
rect 22112 38758 22140 39034
rect 22100 38752 22152 38758
rect 22100 38694 22152 38700
rect 21916 38412 21968 38418
rect 21916 38354 21968 38360
rect 21916 38208 21968 38214
rect 21916 38150 21968 38156
rect 21548 38004 21600 38010
rect 21548 37946 21600 37952
rect 21456 37936 21508 37942
rect 21456 37878 21508 37884
rect 21560 37806 21588 37946
rect 21548 37800 21600 37806
rect 21548 37742 21600 37748
rect 21560 37398 21588 37742
rect 21640 37732 21692 37738
rect 21640 37674 21692 37680
rect 21548 37392 21600 37398
rect 21548 37334 21600 37340
rect 21376 36366 21496 36394
rect 21364 36236 21416 36242
rect 21364 36178 21416 36184
rect 21272 35012 21324 35018
rect 21272 34954 21324 34960
rect 21180 34740 21232 34746
rect 21180 34682 21232 34688
rect 21180 33448 21232 33454
rect 21180 33390 21232 33396
rect 21192 32910 21220 33390
rect 21284 32978 21312 34954
rect 21376 34950 21404 36178
rect 21364 34944 21416 34950
rect 21364 34886 21416 34892
rect 21376 34066 21404 34886
rect 21364 34060 21416 34066
rect 21364 34002 21416 34008
rect 21376 33658 21404 34002
rect 21468 33998 21496 36366
rect 21548 35692 21600 35698
rect 21548 35634 21600 35640
rect 21456 33992 21508 33998
rect 21456 33934 21508 33940
rect 21456 33856 21508 33862
rect 21456 33798 21508 33804
rect 21468 33658 21496 33798
rect 21364 33652 21416 33658
rect 21364 33594 21416 33600
rect 21456 33652 21508 33658
rect 21456 33594 21508 33600
rect 21362 33552 21418 33561
rect 21362 33487 21418 33496
rect 21456 33516 21508 33522
rect 21376 33318 21404 33487
rect 21456 33458 21508 33464
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21376 33017 21404 33254
rect 21362 33008 21418 33017
rect 21272 32972 21324 32978
rect 21362 32943 21418 32952
rect 21272 32914 21324 32920
rect 21180 32904 21232 32910
rect 21180 32846 21232 32852
rect 21270 32736 21326 32745
rect 21270 32671 21326 32680
rect 21088 32564 21140 32570
rect 21088 32506 21140 32512
rect 21180 32564 21232 32570
rect 21180 32506 21232 32512
rect 21088 32428 21140 32434
rect 21088 32370 21140 32376
rect 20996 32224 21048 32230
rect 20996 32166 21048 32172
rect 21008 31958 21036 32166
rect 20996 31952 21048 31958
rect 20996 31894 21048 31900
rect 20904 31816 20956 31822
rect 20904 31758 20956 31764
rect 21100 30394 21128 32370
rect 21088 30388 21140 30394
rect 21088 30330 21140 30336
rect 21192 29866 21220 32506
rect 21100 29838 21220 29866
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20904 29504 20956 29510
rect 20904 29446 20956 29452
rect 20916 29306 20944 29446
rect 20904 29300 20956 29306
rect 20904 29242 20956 29248
rect 21100 28150 21128 29838
rect 21180 29708 21232 29714
rect 21180 29650 21232 29656
rect 21192 28762 21220 29650
rect 21180 28756 21232 28762
rect 21180 28698 21232 28704
rect 21088 28144 21140 28150
rect 21088 28086 21140 28092
rect 20628 27532 20680 27538
rect 20628 27474 20680 27480
rect 20640 26858 20668 27474
rect 21192 26926 21220 28698
rect 21284 27470 21312 32671
rect 21468 32434 21496 33458
rect 21560 32978 21588 35634
rect 21652 35290 21680 37674
rect 21732 36372 21784 36378
rect 21732 36314 21784 36320
rect 21640 35284 21692 35290
rect 21640 35226 21692 35232
rect 21652 34610 21680 35226
rect 21640 34604 21692 34610
rect 21640 34546 21692 34552
rect 21744 34490 21772 36314
rect 21824 36100 21876 36106
rect 21824 36042 21876 36048
rect 21652 34462 21772 34490
rect 21548 32972 21600 32978
rect 21548 32914 21600 32920
rect 21456 32428 21508 32434
rect 21456 32370 21508 32376
rect 21364 32360 21416 32366
rect 21364 32302 21416 32308
rect 21376 32230 21404 32302
rect 21560 32230 21588 32914
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 21548 32224 21600 32230
rect 21548 32166 21600 32172
rect 21456 31476 21508 31482
rect 21456 31418 21508 31424
rect 21364 31408 21416 31414
rect 21364 31350 21416 31356
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 20628 26852 20680 26858
rect 20628 26794 20680 26800
rect 21192 26314 21220 26862
rect 21180 26308 21232 26314
rect 21180 26250 21232 26256
rect 21376 25974 21404 31350
rect 21468 29510 21496 31418
rect 21560 31346 21588 32166
rect 21652 31822 21680 34462
rect 21640 31816 21692 31822
rect 21640 31758 21692 31764
rect 21652 31482 21680 31758
rect 21836 31754 21864 36042
rect 21928 34066 21956 38150
rect 22008 37664 22060 37670
rect 22008 37606 22060 37612
rect 22020 34524 22048 37606
rect 22204 35834 22232 39222
rect 22284 38480 22336 38486
rect 22284 38422 22336 38428
rect 22296 36689 22324 38422
rect 22388 37788 22416 40174
rect 22466 40080 22522 40089
rect 22466 40015 22522 40024
rect 22480 37942 22508 40015
rect 22468 37936 22520 37942
rect 22468 37878 22520 37884
rect 22468 37800 22520 37806
rect 22388 37760 22468 37788
rect 22468 37742 22520 37748
rect 22282 36680 22338 36689
rect 22480 36650 22508 37742
rect 22282 36615 22338 36624
rect 22468 36644 22520 36650
rect 22468 36586 22520 36592
rect 22284 36032 22336 36038
rect 22284 35974 22336 35980
rect 22192 35828 22244 35834
rect 22192 35770 22244 35776
rect 22100 35692 22152 35698
rect 22100 35634 22152 35640
rect 22192 35692 22244 35698
rect 22192 35634 22244 35640
rect 22112 34678 22140 35634
rect 22204 35086 22232 35634
rect 22192 35080 22244 35086
rect 22192 35022 22244 35028
rect 22100 34672 22152 34678
rect 22100 34614 22152 34620
rect 22020 34496 22140 34524
rect 22008 34400 22060 34406
rect 22008 34342 22060 34348
rect 21916 34060 21968 34066
rect 21916 34002 21968 34008
rect 21916 32768 21968 32774
rect 21914 32736 21916 32745
rect 21968 32736 21970 32745
rect 21914 32671 21970 32680
rect 21914 32600 21970 32609
rect 21914 32535 21916 32544
rect 21968 32535 21970 32544
rect 21916 32506 21968 32512
rect 21824 31748 21876 31754
rect 21824 31690 21876 31696
rect 21640 31476 21692 31482
rect 21640 31418 21692 31424
rect 21548 31340 21600 31346
rect 21548 31282 21600 31288
rect 21824 30592 21876 30598
rect 21824 30534 21876 30540
rect 21640 30116 21692 30122
rect 21640 30058 21692 30064
rect 21652 29782 21680 30058
rect 21732 30048 21784 30054
rect 21732 29990 21784 29996
rect 21640 29776 21692 29782
rect 21640 29718 21692 29724
rect 21456 29504 21508 29510
rect 21456 29446 21508 29452
rect 21548 29232 21600 29238
rect 21546 29200 21548 29209
rect 21600 29200 21602 29209
rect 21546 29135 21602 29144
rect 21640 27668 21692 27674
rect 21640 27610 21692 27616
rect 21548 27600 21600 27606
rect 21548 27542 21600 27548
rect 21364 25968 21416 25974
rect 21364 25910 21416 25916
rect 21272 25832 21324 25838
rect 21272 25774 21324 25780
rect 21284 25294 21312 25774
rect 21364 25696 21416 25702
rect 21364 25638 21416 25644
rect 21272 25288 21324 25294
rect 21272 25230 21324 25236
rect 20536 24676 20588 24682
rect 20536 24618 20588 24624
rect 20548 23798 20576 24618
rect 20536 23792 20588 23798
rect 20536 23734 20588 23740
rect 20456 23582 20576 23610
rect 20444 23316 20496 23322
rect 20444 23258 20496 23264
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 19904 22066 20024 22094
rect 19996 21894 20024 22066
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 20168 21548 20220 21554
rect 20168 21490 20220 21496
rect 20180 20874 20208 21490
rect 20364 21434 20392 22714
rect 20456 21554 20484 23258
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20260 21412 20312 21418
rect 20364 21406 20484 21434
rect 20260 21354 20312 21360
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20272 20777 20300 21354
rect 20456 21350 20484 21406
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 19982 20768 20038 20777
rect 19982 20703 20038 20712
rect 20258 20768 20314 20777
rect 20258 20703 20314 20712
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 19530 19380 19654
rect 19352 19514 19564 19530
rect 19352 19508 19576 19514
rect 19352 19502 19524 19508
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 18880 17604 18932 17610
rect 18880 17546 18932 17552
rect 18892 15162 18920 17546
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18708 15014 18828 15042
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17880 11898 17908 12106
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18340 11898 18368 12718
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18524 11830 18552 13330
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18340 10674 18368 11494
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18248 10130 18276 10406
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17420 9574 17632 9602
rect 17420 3534 17448 9574
rect 17592 9444 17644 9450
rect 17592 9386 17644 9392
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17144 800 17172 2858
rect 17512 800 17540 4014
rect 17604 2774 17632 9386
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 5710 17724 9318
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17788 4826 17816 5170
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 18340 4622 18368 6598
rect 18616 4622 18644 12582
rect 18708 10062 18736 15014
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18708 4049 18736 4082
rect 18694 4040 18750 4049
rect 18694 3975 18750 3984
rect 18708 3738 18736 3975
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17604 2746 17724 2774
rect 17696 2582 17724 2746
rect 17684 2576 17736 2582
rect 17684 2518 17736 2524
rect 17880 800 17908 3538
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17972 2514 18000 2790
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18340 1170 18368 2314
rect 18248 1142 18368 1170
rect 18248 800 18276 1142
rect 18616 800 18644 3334
rect 18800 3058 18828 14894
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18892 12238 18920 14758
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 19076 9586 19104 18838
rect 19168 18358 19196 19246
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 19168 17134 19196 18294
rect 19260 17882 19288 19178
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19260 16946 19288 17818
rect 19168 16918 19288 16946
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 19168 8566 19196 16918
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19260 13530 19288 14010
rect 19352 13870 19380 19502
rect 19524 19450 19576 19456
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19444 18358 19472 18634
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19352 10674 19380 13398
rect 19444 13326 19472 14214
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19156 8560 19208 8566
rect 19156 8502 19208 8508
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18800 2650 18828 2994
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 18984 800 19012 3606
rect 19352 800 19380 5238
rect 19444 2774 19472 9930
rect 19536 5234 19564 18566
rect 19628 14260 19656 20470
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19720 16046 19748 16730
rect 19708 16040 19760 16046
rect 19708 15982 19760 15988
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19720 15094 19748 15302
rect 19708 15088 19760 15094
rect 19708 15030 19760 15036
rect 19812 15026 19840 20198
rect 19892 15632 19944 15638
rect 19892 15574 19944 15580
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19708 14272 19760 14278
rect 19628 14232 19708 14260
rect 19708 14214 19760 14220
rect 19720 14006 19748 14214
rect 19708 14000 19760 14006
rect 19708 13942 19760 13948
rect 19812 12434 19840 14758
rect 19904 13258 19932 15574
rect 19996 14006 20024 20703
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20180 17610 20208 18022
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 20180 16794 20208 17546
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 19892 13252 19944 13258
rect 19892 13194 19944 13200
rect 19812 12406 19932 12434
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11830 19840 12038
rect 19800 11824 19852 11830
rect 19800 11766 19852 11772
rect 19904 11694 19932 12406
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19996 11898 20024 12242
rect 20180 12170 20208 16390
rect 20272 13938 20300 20703
rect 20456 18766 20484 21286
rect 20548 20058 20576 23582
rect 21088 23520 21140 23526
rect 21088 23462 21140 23468
rect 21100 22982 21128 23462
rect 21088 22976 21140 22982
rect 21088 22918 21140 22924
rect 21180 22568 21232 22574
rect 21180 22510 21232 22516
rect 21192 22234 21220 22510
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20548 19514 20576 19994
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20640 17882 20668 19246
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 20732 17610 20760 18566
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20732 17270 20760 17546
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20456 16590 20484 17070
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20824 16182 20852 19314
rect 20996 19236 21048 19242
rect 20996 19178 21048 19184
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20916 17746 20944 18634
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20916 17338 20944 17682
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20916 16658 20944 17274
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20812 16176 20864 16182
rect 20812 16118 20864 16124
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19628 10810 19656 10950
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19904 7886 19932 11630
rect 19996 10606 20024 11834
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 20364 5710 20392 13806
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 10674 20576 12582
rect 20640 11150 20668 15302
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20732 13530 20760 13874
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20824 11830 20852 14418
rect 20916 14414 20944 16594
rect 21008 15638 21036 19178
rect 21100 16250 21128 19314
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 20996 15632 21048 15638
rect 20996 15574 21048 15580
rect 21192 15570 21220 16390
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21192 14482 21220 15506
rect 21284 15502 21312 21286
rect 21376 19514 21404 25638
rect 21560 21894 21588 27542
rect 21652 26314 21680 27610
rect 21640 26308 21692 26314
rect 21640 26250 21692 26256
rect 21652 24138 21680 26250
rect 21744 24206 21772 29990
rect 21836 26568 21864 30534
rect 22020 29646 22048 34342
rect 22112 33522 22140 34496
rect 22204 33522 22232 35022
rect 22296 34746 22324 35974
rect 22468 35624 22520 35630
rect 22468 35566 22520 35572
rect 22376 35556 22428 35562
rect 22376 35498 22428 35504
rect 22388 34950 22416 35498
rect 22376 34944 22428 34950
rect 22376 34886 22428 34892
rect 22284 34740 22336 34746
rect 22284 34682 22336 34688
rect 22480 34678 22508 35566
rect 22572 35562 22600 41386
rect 22664 41070 22692 43182
rect 22756 41682 22784 46310
rect 22848 43654 22876 51870
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 23860 45554 23888 53926
rect 23940 52896 23992 52902
rect 23940 52838 23992 52844
rect 23584 45526 23888 45554
rect 23388 45348 23440 45354
rect 23388 45290 23440 45296
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 23400 44742 23428 45290
rect 23388 44736 23440 44742
rect 23388 44678 23440 44684
rect 23296 44192 23348 44198
rect 23296 44134 23348 44140
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 23308 43994 23336 44134
rect 23296 43988 23348 43994
rect 23296 43930 23348 43936
rect 23296 43852 23348 43858
rect 23296 43794 23348 43800
rect 22836 43648 22888 43654
rect 22836 43590 22888 43596
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22836 42696 22888 42702
rect 22836 42638 22888 42644
rect 22848 42158 22876 42638
rect 23308 42362 23336 43794
rect 23296 42356 23348 42362
rect 23296 42298 23348 42304
rect 22836 42152 22888 42158
rect 22836 42094 22888 42100
rect 22744 41676 22796 41682
rect 22744 41618 22796 41624
rect 22848 41070 22876 42094
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22652 41064 22704 41070
rect 22652 41006 22704 41012
rect 22836 41064 22888 41070
rect 22836 41006 22888 41012
rect 22744 40724 22796 40730
rect 22744 40666 22796 40672
rect 22652 40180 22704 40186
rect 22652 40122 22704 40128
rect 22664 39982 22692 40122
rect 22756 40050 22784 40666
rect 22848 40118 22876 41006
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 23020 40520 23072 40526
rect 23020 40462 23072 40468
rect 22836 40112 22888 40118
rect 22836 40054 22888 40060
rect 22744 40044 22796 40050
rect 22744 39986 22796 39992
rect 22652 39976 22704 39982
rect 22652 39918 22704 39924
rect 22756 39370 22784 39986
rect 23032 39982 23060 40462
rect 23020 39976 23072 39982
rect 23020 39918 23072 39924
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 23308 39386 23336 42298
rect 23400 40594 23428 44678
rect 23480 43988 23532 43994
rect 23480 43930 23532 43936
rect 23492 43246 23520 43930
rect 23480 43240 23532 43246
rect 23480 43182 23532 43188
rect 23492 42158 23520 43182
rect 23480 42152 23532 42158
rect 23480 42094 23532 42100
rect 23480 41676 23532 41682
rect 23480 41618 23532 41624
rect 23492 41274 23520 41618
rect 23480 41268 23532 41274
rect 23480 41210 23532 41216
rect 23388 40588 23440 40594
rect 23388 40530 23440 40536
rect 23388 40384 23440 40390
rect 23388 40326 23440 40332
rect 22744 39364 22796 39370
rect 22744 39306 22796 39312
rect 23124 39358 23336 39386
rect 23124 38894 23152 39358
rect 23294 39264 23350 39273
rect 23294 39199 23350 39208
rect 23112 38888 23164 38894
rect 23112 38830 23164 38836
rect 22836 38752 22888 38758
rect 22836 38694 22888 38700
rect 22652 38412 22704 38418
rect 22652 38354 22704 38360
rect 22560 35556 22612 35562
rect 22560 35498 22612 35504
rect 22558 35456 22614 35465
rect 22558 35391 22614 35400
rect 22468 34672 22520 34678
rect 22468 34614 22520 34620
rect 22468 34536 22520 34542
rect 22468 34478 22520 34484
rect 22480 34202 22508 34478
rect 22468 34196 22520 34202
rect 22468 34138 22520 34144
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22100 33516 22152 33522
rect 22100 33458 22152 33464
rect 22192 33516 22244 33522
rect 22192 33458 22244 33464
rect 22100 33040 22152 33046
rect 22100 32982 22152 32988
rect 22112 32502 22140 32982
rect 22100 32496 22152 32502
rect 22100 32438 22152 32444
rect 22204 31278 22232 33458
rect 22284 33312 22336 33318
rect 22284 33254 22336 33260
rect 22296 33046 22324 33254
rect 22374 33144 22430 33153
rect 22480 33114 22508 33798
rect 22374 33079 22430 33088
rect 22468 33108 22520 33114
rect 22284 33040 22336 33046
rect 22284 32982 22336 32988
rect 22388 32910 22416 33079
rect 22468 33050 22520 33056
rect 22466 33008 22522 33017
rect 22466 32943 22522 32952
rect 22376 32904 22428 32910
rect 22376 32846 22428 32852
rect 22374 32736 22430 32745
rect 22374 32671 22430 32680
rect 22388 32570 22416 32671
rect 22376 32564 22428 32570
rect 22376 32506 22428 32512
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22296 31754 22324 32438
rect 22284 31748 22336 31754
rect 22284 31690 22336 31696
rect 22192 31272 22244 31278
rect 22192 31214 22244 31220
rect 22204 30258 22232 31214
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 22284 29640 22336 29646
rect 22284 29582 22336 29588
rect 22008 28620 22060 28626
rect 22008 28562 22060 28568
rect 22020 28082 22048 28562
rect 22192 28484 22244 28490
rect 22192 28426 22244 28432
rect 22204 28150 22232 28426
rect 22192 28144 22244 28150
rect 22192 28086 22244 28092
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 22020 27554 22048 28018
rect 22204 27674 22232 28086
rect 22192 27668 22244 27674
rect 22192 27610 22244 27616
rect 21928 27538 22048 27554
rect 21916 27532 22048 27538
rect 21968 27526 22048 27532
rect 21916 27474 21968 27480
rect 22020 26926 22048 27526
rect 22100 27396 22152 27402
rect 22100 27338 22152 27344
rect 22192 27396 22244 27402
rect 22192 27338 22244 27344
rect 22008 26920 22060 26926
rect 22008 26862 22060 26868
rect 21916 26580 21968 26586
rect 21836 26540 21916 26568
rect 21916 26522 21968 26528
rect 22020 26518 22048 26862
rect 22008 26512 22060 26518
rect 22008 26454 22060 26460
rect 22020 24818 22048 26454
rect 22112 25226 22140 27338
rect 22204 26518 22232 27338
rect 22192 26512 22244 26518
rect 22192 26454 22244 26460
rect 22204 25906 22232 26454
rect 22296 25906 22324 29582
rect 22388 26042 22416 32506
rect 22480 30734 22508 32943
rect 22572 32434 22600 35391
rect 22664 35018 22692 38354
rect 22744 37868 22796 37874
rect 22744 37810 22796 37816
rect 22652 35012 22704 35018
rect 22652 34954 22704 34960
rect 22652 34536 22704 34542
rect 22652 34478 22704 34484
rect 22560 32428 22612 32434
rect 22560 32370 22612 32376
rect 22560 32224 22612 32230
rect 22560 32166 22612 32172
rect 22572 32026 22600 32166
rect 22560 32020 22612 32026
rect 22560 31962 22612 31968
rect 22664 31142 22692 34478
rect 22756 32774 22784 37810
rect 22848 37806 22876 38694
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 23308 37874 23336 39199
rect 23296 37868 23348 37874
rect 23296 37810 23348 37816
rect 22836 37800 22888 37806
rect 22836 37742 22888 37748
rect 22848 37194 22876 37742
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 22836 37188 22888 37194
rect 22836 37130 22888 37136
rect 22848 36718 22876 37130
rect 22836 36712 22888 36718
rect 22836 36654 22888 36660
rect 22848 35698 22876 36654
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 23204 36372 23256 36378
rect 23204 36314 23256 36320
rect 23216 36038 23244 36314
rect 23204 36032 23256 36038
rect 23204 35974 23256 35980
rect 23400 35714 23428 40326
rect 23492 39506 23520 41210
rect 23480 39500 23532 39506
rect 23480 39442 23532 39448
rect 23584 38978 23612 45526
rect 23848 43240 23900 43246
rect 23848 43182 23900 43188
rect 23664 42696 23716 42702
rect 23664 42638 23716 42644
rect 23756 42696 23808 42702
rect 23756 42638 23808 42644
rect 23676 40186 23704 42638
rect 23768 41614 23796 42638
rect 23860 41682 23888 43182
rect 23848 41676 23900 41682
rect 23848 41618 23900 41624
rect 23756 41608 23808 41614
rect 23756 41550 23808 41556
rect 23768 40712 23796 41550
rect 23848 41472 23900 41478
rect 23848 41414 23900 41420
rect 23860 41313 23888 41414
rect 23846 41304 23902 41313
rect 23846 41239 23902 41248
rect 23768 40684 23888 40712
rect 23756 40452 23808 40458
rect 23756 40394 23808 40400
rect 23768 40186 23796 40394
rect 23664 40180 23716 40186
rect 23664 40122 23716 40128
rect 23756 40180 23808 40186
rect 23756 40122 23808 40128
rect 23756 39840 23808 39846
rect 23676 39800 23756 39828
rect 23676 39030 23704 39800
rect 23756 39782 23808 39788
rect 23860 39273 23888 40684
rect 23952 39953 23980 52838
rect 24044 52698 24072 54130
rect 24596 53582 24624 56199
rect 24674 55448 24730 55457
rect 24674 55383 24730 55392
rect 24688 54194 24716 55383
rect 24766 54632 24822 54641
rect 24766 54567 24822 54576
rect 24676 54188 24728 54194
rect 24676 54130 24728 54136
rect 24674 53816 24730 53825
rect 24674 53751 24730 53760
rect 24584 53576 24636 53582
rect 24584 53518 24636 53524
rect 24596 52698 24624 53518
rect 24032 52692 24084 52698
rect 24032 52634 24084 52640
rect 24584 52692 24636 52698
rect 24584 52634 24636 52640
rect 24688 52018 24716 53751
rect 24780 53106 24808 54567
rect 25044 54052 25096 54058
rect 25044 53994 25096 54000
rect 25056 53106 25084 53994
rect 25964 53576 26016 53582
rect 25964 53518 26016 53524
rect 24768 53100 24820 53106
rect 24768 53042 24820 53048
rect 25044 53100 25096 53106
rect 25044 53042 25096 53048
rect 24780 52698 24808 53042
rect 25056 53009 25084 53042
rect 25042 53000 25098 53009
rect 25042 52935 25098 52944
rect 24952 52896 25004 52902
rect 24952 52838 25004 52844
rect 24768 52692 24820 52698
rect 24768 52634 24820 52640
rect 24768 52488 24820 52494
rect 24768 52430 24820 52436
rect 24780 52193 24808 52430
rect 24766 52184 24822 52193
rect 24766 52119 24822 52128
rect 24676 52012 24728 52018
rect 24676 51954 24728 51960
rect 24400 47660 24452 47666
rect 24400 47602 24452 47608
rect 24216 46572 24268 46578
rect 24216 46514 24268 46520
rect 24032 45960 24084 45966
rect 24032 45902 24084 45908
rect 23938 39944 23994 39953
rect 23938 39879 23994 39888
rect 23846 39264 23902 39273
rect 23846 39199 23902 39208
rect 23492 38950 23612 38978
rect 23664 39024 23716 39030
rect 23664 38966 23716 38972
rect 23492 37670 23520 38950
rect 23676 38876 23704 38966
rect 23584 38848 23704 38876
rect 23756 38888 23808 38894
rect 23584 38298 23612 38848
rect 23756 38830 23808 38836
rect 23664 38752 23716 38758
rect 23664 38694 23716 38700
rect 23676 38418 23704 38694
rect 23768 38418 23796 38830
rect 23664 38412 23716 38418
rect 23664 38354 23716 38360
rect 23756 38412 23808 38418
rect 23756 38354 23808 38360
rect 23848 38344 23900 38350
rect 23584 38270 23704 38298
rect 23848 38286 23900 38292
rect 23676 38214 23704 38270
rect 23572 38208 23624 38214
rect 23572 38150 23624 38156
rect 23664 38208 23716 38214
rect 23664 38150 23716 38156
rect 23756 38208 23808 38214
rect 23756 38150 23808 38156
rect 23480 37664 23532 37670
rect 23480 37606 23532 37612
rect 23584 37466 23612 38150
rect 23664 37664 23716 37670
rect 23664 37606 23716 37612
rect 23480 37460 23532 37466
rect 23480 37402 23532 37408
rect 23572 37460 23624 37466
rect 23572 37402 23624 37408
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 23308 35686 23428 35714
rect 22836 35556 22888 35562
rect 22836 35498 22888 35504
rect 22744 32768 22796 32774
rect 22744 32710 22796 32716
rect 22756 32570 22784 32710
rect 22744 32564 22796 32570
rect 22744 32506 22796 32512
rect 22744 32224 22796 32230
rect 22744 32166 22796 32172
rect 22652 31136 22704 31142
rect 22652 31078 22704 31084
rect 22468 30728 22520 30734
rect 22468 30670 22520 30676
rect 22756 30002 22784 32166
rect 22664 29974 22784 30002
rect 22560 29708 22612 29714
rect 22560 29650 22612 29656
rect 22468 29096 22520 29102
rect 22468 29038 22520 29044
rect 22480 26314 22508 29038
rect 22572 26602 22600 29650
rect 22664 27538 22692 29974
rect 22848 29866 22876 35498
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23204 34944 23256 34950
rect 23204 34886 23256 34892
rect 23216 34490 23244 34886
rect 23308 34610 23336 35686
rect 23388 35624 23440 35630
rect 23388 35566 23440 35572
rect 23400 34950 23428 35566
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 23296 34604 23348 34610
rect 23296 34546 23348 34552
rect 23216 34462 23336 34490
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23308 31482 23336 34462
rect 23400 34066 23428 34886
rect 23492 34626 23520 37402
rect 23572 36712 23624 36718
rect 23572 36654 23624 36660
rect 23584 35834 23612 36654
rect 23676 36122 23704 37606
rect 23768 36242 23796 38150
rect 23860 37806 23888 38286
rect 23952 38282 23980 39879
rect 23940 38276 23992 38282
rect 23940 38218 23992 38224
rect 23848 37800 23900 37806
rect 23848 37742 23900 37748
rect 23860 36718 23888 37742
rect 24044 37330 24072 45902
rect 24228 41414 24256 46514
rect 24308 45280 24360 45286
rect 24308 45222 24360 45228
rect 24320 44742 24348 45222
rect 24308 44736 24360 44742
rect 24308 44678 24360 44684
rect 24320 44470 24348 44678
rect 24308 44464 24360 44470
rect 24308 44406 24360 44412
rect 24320 43654 24348 44406
rect 24308 43648 24360 43654
rect 24308 43590 24360 43596
rect 24320 43382 24348 43590
rect 24308 43376 24360 43382
rect 24308 43318 24360 43324
rect 24320 42770 24348 43318
rect 24308 42764 24360 42770
rect 24308 42706 24360 42712
rect 24320 42294 24348 42706
rect 24308 42288 24360 42294
rect 24308 42230 24360 42236
rect 24320 41478 24348 42230
rect 24308 41472 24360 41478
rect 24308 41414 24360 41420
rect 24136 41386 24256 41414
rect 24032 37324 24084 37330
rect 24032 37266 24084 37272
rect 23940 37120 23992 37126
rect 23940 37062 23992 37068
rect 23952 36922 23980 37062
rect 23940 36916 23992 36922
rect 23940 36858 23992 36864
rect 23848 36712 23900 36718
rect 23848 36654 23900 36660
rect 23756 36236 23808 36242
rect 23756 36178 23808 36184
rect 23676 36094 23796 36122
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23572 35828 23624 35834
rect 23572 35770 23624 35776
rect 23676 34746 23704 35974
rect 23664 34740 23716 34746
rect 23664 34682 23716 34688
rect 23492 34598 23612 34626
rect 23480 34536 23532 34542
rect 23480 34478 23532 34484
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23388 33924 23440 33930
rect 23388 33866 23440 33872
rect 23400 32042 23428 33866
rect 23492 33386 23520 34478
rect 23480 33380 23532 33386
rect 23480 33322 23532 33328
rect 23584 33114 23612 34598
rect 23768 33538 23796 36094
rect 23860 34542 23888 36654
rect 24136 36174 24164 41386
rect 24412 40526 24440 47602
rect 24768 46980 24820 46986
rect 24768 46922 24820 46928
rect 24492 46504 24544 46510
rect 24780 46481 24808 46922
rect 24492 46446 24544 46452
rect 24766 46472 24822 46481
rect 24504 46170 24532 46446
rect 24766 46407 24822 46416
rect 24492 46164 24544 46170
rect 24492 46106 24544 46112
rect 24860 45824 24912 45830
rect 24860 45766 24912 45772
rect 24872 45665 24900 45766
rect 24858 45656 24914 45665
rect 24858 45591 24914 45600
rect 24964 45554 24992 52838
rect 25136 52624 25188 52630
rect 25136 52566 25188 52572
rect 25044 51400 25096 51406
rect 25042 51368 25044 51377
rect 25096 51368 25098 51377
rect 25042 51303 25098 51312
rect 25044 50924 25096 50930
rect 25044 50866 25096 50872
rect 25056 50561 25084 50866
rect 25042 50552 25098 50561
rect 25042 50487 25098 50496
rect 25148 48314 25176 52566
rect 25780 51808 25832 51814
rect 25780 51750 25832 51756
rect 25688 50720 25740 50726
rect 25688 50662 25740 50668
rect 25320 50176 25372 50182
rect 25320 50118 25372 50124
rect 25332 49842 25360 50118
rect 25320 49836 25372 49842
rect 25320 49778 25372 49784
rect 25332 49745 25360 49778
rect 25318 49736 25374 49745
rect 25318 49671 25374 49680
rect 25320 49224 25372 49230
rect 25320 49166 25372 49172
rect 25332 48929 25360 49166
rect 25318 48920 25374 48929
rect 25318 48855 25374 48864
rect 25504 48544 25556 48550
rect 25504 48486 25556 48492
rect 25148 48286 25452 48314
rect 25320 48136 25372 48142
rect 25318 48104 25320 48113
rect 25372 48104 25374 48113
rect 25318 48039 25374 48048
rect 24872 45526 24992 45554
rect 24492 45416 24544 45422
rect 24492 45358 24544 45364
rect 24676 45416 24728 45422
rect 24676 45358 24728 45364
rect 24504 44742 24532 45358
rect 24492 44736 24544 44742
rect 24492 44678 24544 44684
rect 24490 41304 24546 41313
rect 24490 41239 24546 41248
rect 24504 41206 24532 41239
rect 24492 41200 24544 41206
rect 24492 41142 24544 41148
rect 24400 40520 24452 40526
rect 24400 40462 24452 40468
rect 24504 40390 24532 41142
rect 24216 40384 24268 40390
rect 24216 40326 24268 40332
rect 24492 40384 24544 40390
rect 24584 40384 24636 40390
rect 24492 40326 24544 40332
rect 24582 40352 24584 40361
rect 24636 40352 24638 40361
rect 24228 38962 24256 40326
rect 24504 40118 24532 40326
rect 24582 40287 24638 40296
rect 24492 40112 24544 40118
rect 24544 40060 24624 40066
rect 24492 40054 24624 40060
rect 24504 40038 24624 40054
rect 24492 39976 24544 39982
rect 24492 39918 24544 39924
rect 24216 38956 24268 38962
rect 24216 38898 24268 38904
rect 24504 37806 24532 39918
rect 24596 38894 24624 40038
rect 24584 38888 24636 38894
rect 24584 38830 24636 38836
rect 24596 37942 24624 38830
rect 24688 38486 24716 45358
rect 24768 44328 24820 44334
rect 24768 44270 24820 44276
rect 24780 43217 24808 44270
rect 24766 43208 24822 43217
rect 24766 43143 24822 43152
rect 24872 42702 24900 45526
rect 25320 44396 25372 44402
rect 25320 44338 25372 44344
rect 25332 43654 25360 44338
rect 25320 43648 25372 43654
rect 25320 43590 25372 43596
rect 25332 43217 25360 43590
rect 25318 43208 25374 43217
rect 25318 43143 25374 43152
rect 24952 43104 25004 43110
rect 24952 43046 25004 43052
rect 25228 43104 25280 43110
rect 25228 43046 25280 43052
rect 24860 42696 24912 42702
rect 24860 42638 24912 42644
rect 24860 42560 24912 42566
rect 24860 42502 24912 42508
rect 24872 42401 24900 42502
rect 24858 42392 24914 42401
rect 24858 42327 24914 42336
rect 24860 41472 24912 41478
rect 24860 41414 24912 41420
rect 24872 41070 24900 41414
rect 24860 41064 24912 41070
rect 24860 41006 24912 41012
rect 24768 40520 24820 40526
rect 24768 40462 24820 40468
rect 24780 39953 24808 40462
rect 24766 39944 24822 39953
rect 24766 39879 24822 39888
rect 24768 39296 24820 39302
rect 24768 39238 24820 39244
rect 24676 38480 24728 38486
rect 24676 38422 24728 38428
rect 24676 38208 24728 38214
rect 24676 38150 24728 38156
rect 24688 38010 24716 38150
rect 24676 38004 24728 38010
rect 24676 37946 24728 37952
rect 24584 37936 24636 37942
rect 24636 37884 24716 37890
rect 24584 37878 24716 37884
rect 24596 37862 24716 37878
rect 24492 37800 24544 37806
rect 24492 37742 24544 37748
rect 24400 36304 24452 36310
rect 24400 36246 24452 36252
rect 24124 36168 24176 36174
rect 24124 36110 24176 36116
rect 24308 34944 24360 34950
rect 24308 34886 24360 34892
rect 23848 34536 23900 34542
rect 23848 34478 23900 34484
rect 23848 34128 23900 34134
rect 23848 34070 23900 34076
rect 23676 33510 23796 33538
rect 23572 33108 23624 33114
rect 23572 33050 23624 33056
rect 23676 33046 23704 33510
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 23664 33040 23716 33046
rect 23664 32982 23716 32988
rect 23400 32014 23612 32042
rect 23584 31958 23612 32014
rect 23388 31952 23440 31958
rect 23388 31894 23440 31900
rect 23572 31952 23624 31958
rect 23572 31894 23624 31900
rect 23296 31476 23348 31482
rect 23296 31418 23348 31424
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 22756 29838 22876 29866
rect 22756 29170 22784 29838
rect 22836 29776 22888 29782
rect 22836 29718 22888 29724
rect 22848 29306 22876 29718
rect 23400 29714 23428 31894
rect 23480 31884 23532 31890
rect 23480 31826 23532 31832
rect 23492 31226 23520 31826
rect 23492 31198 23612 31226
rect 23584 31142 23612 31198
rect 23572 31136 23624 31142
rect 23572 31078 23624 31084
rect 23584 30326 23612 31078
rect 23572 30320 23624 30326
rect 23572 30262 23624 30268
rect 23388 29708 23440 29714
rect 23388 29650 23440 29656
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 23308 29034 23336 29446
rect 23584 29102 23612 30262
rect 23768 30190 23796 33390
rect 23860 30734 23888 34070
rect 24320 33930 24348 34886
rect 24032 33924 24084 33930
rect 24032 33866 24084 33872
rect 24308 33924 24360 33930
rect 24308 33866 24360 33872
rect 24044 33590 24072 33866
rect 24032 33584 24084 33590
rect 23952 33532 24032 33538
rect 23952 33526 24084 33532
rect 23952 33510 24072 33526
rect 23952 31822 23980 33510
rect 24032 32972 24084 32978
rect 24032 32914 24084 32920
rect 23940 31816 23992 31822
rect 23940 31758 23992 31764
rect 23952 31414 23980 31758
rect 23940 31408 23992 31414
rect 23940 31350 23992 31356
rect 23848 30728 23900 30734
rect 23848 30670 23900 30676
rect 23952 30394 23980 31350
rect 23940 30388 23992 30394
rect 23940 30330 23992 30336
rect 23756 30184 23808 30190
rect 23756 30126 23808 30132
rect 23768 29714 23796 30126
rect 23756 29708 23808 29714
rect 23756 29650 23808 29656
rect 23572 29096 23624 29102
rect 23572 29038 23624 29044
rect 23296 29028 23348 29034
rect 23296 28970 23348 28976
rect 23388 29028 23440 29034
rect 23388 28970 23440 28976
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 23400 28234 23428 28970
rect 23308 28206 23428 28234
rect 22744 27872 22796 27878
rect 22744 27814 22796 27820
rect 22652 27532 22704 27538
rect 22652 27474 22704 27480
rect 22572 26574 22692 26602
rect 22560 26512 22612 26518
rect 22560 26454 22612 26460
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 22376 26036 22428 26042
rect 22376 25978 22428 25984
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22284 25764 22336 25770
rect 22284 25706 22336 25712
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 22112 24682 22140 24754
rect 22100 24676 22152 24682
rect 22100 24618 22152 24624
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 21836 24138 21864 24346
rect 22112 24274 22140 24618
rect 22100 24268 22152 24274
rect 22100 24210 22152 24216
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 21652 23866 21680 24074
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 22112 23730 22140 24210
rect 22192 24132 22244 24138
rect 22192 24074 22244 24080
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22020 22642 22048 23666
rect 22204 23066 22232 24074
rect 22112 23038 22232 23066
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21652 20806 21680 22510
rect 22020 22098 22048 22578
rect 22008 22092 22060 22098
rect 22008 22034 22060 22040
rect 22020 21622 22048 22034
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21652 20398 21680 20742
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 21928 19310 21956 19450
rect 21916 19304 21968 19310
rect 21916 19246 21968 19252
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 21928 18612 21956 19246
rect 22020 18766 22048 19246
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 21928 18584 22048 18612
rect 21456 18148 21508 18154
rect 21456 18090 21508 18096
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20916 12986 20944 14350
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 21008 12986 21036 13262
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21192 12782 21220 13126
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20640 10554 20668 11086
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20548 10526 20668 10554
rect 20824 10538 20852 11018
rect 20812 10532 20864 10538
rect 20548 7886 20576 10526
rect 20812 10474 20864 10480
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20640 8974 20668 10406
rect 21008 10198 21036 12038
rect 20996 10192 21048 10198
rect 20996 10134 21048 10140
rect 21100 9586 21128 12038
rect 21192 11898 21220 12718
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 21284 8566 21312 14758
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 21376 10062 21404 13194
rect 21468 12918 21496 18090
rect 21732 17060 21784 17066
rect 21732 17002 21784 17008
rect 21548 15428 21600 15434
rect 21548 15370 21600 15376
rect 21456 12912 21508 12918
rect 21456 12854 21508 12860
rect 21560 12306 21588 15370
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 21272 8560 21324 8566
rect 21272 8502 21324 8508
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20732 7410 20760 8298
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19708 3460 19760 3466
rect 19708 3402 19760 3408
rect 19444 2746 19564 2774
rect 19536 2446 19564 2746
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19720 800 19748 3402
rect 19904 3398 19932 4626
rect 20168 4548 20220 4554
rect 20168 4490 20220 4496
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 20088 800 20116 4014
rect 20180 2990 20208 4490
rect 20272 4146 20300 5102
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 20456 800 20484 5714
rect 20640 5710 20668 7210
rect 20824 6798 20852 7686
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20732 4010 20760 6190
rect 20916 5914 20944 7278
rect 21100 6322 21128 7686
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 21180 5636 21232 5642
rect 21180 5578 21232 5584
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 20824 800 20852 2790
rect 21192 800 21220 5578
rect 21284 4622 21312 8298
rect 21364 7336 21416 7342
rect 21364 7278 21416 7284
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21376 2417 21404 7278
rect 21456 6248 21508 6254
rect 21456 6190 21508 6196
rect 21468 3194 21496 6190
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21362 2408 21418 2417
rect 21362 2343 21418 2352
rect 21560 800 21588 5714
rect 21652 3534 21680 14554
rect 21744 13326 21772 17002
rect 22020 16658 22048 18584
rect 22112 17202 22140 23038
rect 22296 22930 22324 25706
rect 22388 25498 22416 25978
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 22204 22902 22324 22930
rect 22204 19292 22232 22902
rect 22284 22092 22336 22098
rect 22284 22034 22336 22040
rect 22376 22092 22428 22098
rect 22376 22034 22428 22040
rect 22296 21486 22324 22034
rect 22388 21962 22416 22034
rect 22376 21956 22428 21962
rect 22376 21898 22428 21904
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22388 21146 22416 21898
rect 22572 21690 22600 26454
rect 22664 26246 22692 26574
rect 22652 26240 22704 26246
rect 22652 26182 22704 26188
rect 22664 25362 22692 26182
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 22664 24886 22692 25298
rect 22652 24880 22704 24886
rect 22652 24822 22704 24828
rect 22756 22094 22784 27814
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 22836 27668 22888 27674
rect 22836 27610 22888 27616
rect 22848 27402 22876 27610
rect 22836 27396 22888 27402
rect 22836 27338 22888 27344
rect 23112 27328 23164 27334
rect 23112 27270 23164 27276
rect 23124 27062 23152 27270
rect 23112 27056 23164 27062
rect 23112 26998 23164 27004
rect 23124 26926 23152 26998
rect 23112 26920 23164 26926
rect 23112 26862 23164 26868
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 22836 24744 22888 24750
rect 22836 24686 22888 24692
rect 22848 23866 22876 24686
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23308 24206 23336 28206
rect 23388 27872 23440 27878
rect 23388 27814 23440 27820
rect 23400 27674 23428 27814
rect 23388 27668 23440 27674
rect 23388 27610 23440 27616
rect 23400 27062 23428 27610
rect 23388 27056 23440 27062
rect 23440 27004 23612 27010
rect 23388 26998 23612 27004
rect 23400 26982 23612 26998
rect 23480 26920 23532 26926
rect 23400 26880 23480 26908
rect 23400 26246 23428 26880
rect 23480 26862 23532 26868
rect 23584 26586 23612 26982
rect 23848 26784 23900 26790
rect 23848 26726 23900 26732
rect 23572 26580 23624 26586
rect 23572 26522 23624 26528
rect 23388 26240 23440 26246
rect 23388 26182 23440 26188
rect 23860 25906 23888 26726
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 23400 25498 23428 25842
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 24044 25294 24072 32914
rect 24308 32020 24360 32026
rect 24308 31962 24360 31968
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 24136 27713 24164 29106
rect 24216 28484 24268 28490
rect 24216 28426 24268 28432
rect 24122 27704 24178 27713
rect 24228 27674 24256 28426
rect 24122 27639 24178 27648
rect 24216 27668 24268 27674
rect 24216 27610 24268 27616
rect 24320 25294 24348 31962
rect 24412 31346 24440 36246
rect 24504 36242 24532 37742
rect 24688 37466 24716 37862
rect 24676 37460 24728 37466
rect 24676 37402 24728 37408
rect 24688 36854 24716 37402
rect 24676 36848 24728 36854
rect 24676 36790 24728 36796
rect 24492 36236 24544 36242
rect 24492 36178 24544 36184
rect 24688 35766 24716 36790
rect 24676 35760 24728 35766
rect 24676 35702 24728 35708
rect 24492 34944 24544 34950
rect 24492 34886 24544 34892
rect 24400 31340 24452 31346
rect 24400 31282 24452 31288
rect 24400 31136 24452 31142
rect 24400 31078 24452 31084
rect 24412 26382 24440 31078
rect 24504 30666 24532 34886
rect 24676 34740 24728 34746
rect 24676 34682 24728 34688
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24492 30660 24544 30666
rect 24492 30602 24544 30608
rect 24596 29238 24624 33798
rect 24584 29232 24636 29238
rect 24584 29174 24636 29180
rect 24584 28416 24636 28422
rect 24584 28358 24636 28364
rect 24596 27130 24624 28358
rect 24688 28150 24716 34682
rect 24780 33998 24808 39238
rect 24858 39128 24914 39137
rect 24858 39063 24914 39072
rect 24872 38962 24900 39063
rect 24860 38956 24912 38962
rect 24860 38898 24912 38904
rect 24964 38418 24992 43046
rect 25240 42158 25268 43046
rect 25228 42152 25280 42158
rect 25228 42094 25280 42100
rect 25044 41744 25096 41750
rect 25044 41686 25096 41692
rect 25056 39506 25084 41686
rect 25136 41472 25188 41478
rect 25136 41414 25188 41420
rect 25148 39574 25176 41414
rect 25136 39568 25188 39574
rect 25136 39510 25188 39516
rect 25240 39506 25268 42094
rect 25320 41608 25372 41614
rect 25318 41576 25320 41585
rect 25372 41576 25374 41585
rect 25318 41511 25374 41520
rect 25320 41472 25372 41478
rect 25320 41414 25372 41420
rect 25332 41138 25360 41414
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 25332 40769 25360 41074
rect 25318 40760 25374 40769
rect 25318 40695 25374 40704
rect 25320 40384 25372 40390
rect 25320 40326 25372 40332
rect 25044 39500 25096 39506
rect 25044 39442 25096 39448
rect 25228 39500 25280 39506
rect 25228 39442 25280 39448
rect 25332 38962 25360 40326
rect 25424 39030 25452 48286
rect 25516 47598 25544 48486
rect 25504 47592 25556 47598
rect 25504 47534 25556 47540
rect 25516 47297 25544 47534
rect 25502 47288 25558 47297
rect 25502 47223 25558 47232
rect 25504 46164 25556 46170
rect 25504 46106 25556 46112
rect 25516 44849 25544 46106
rect 25502 44840 25558 44849
rect 25502 44775 25558 44784
rect 25504 44736 25556 44742
rect 25504 44678 25556 44684
rect 25516 44033 25544 44678
rect 25502 44024 25558 44033
rect 25502 43959 25558 43968
rect 25700 40089 25728 50662
rect 25792 40730 25820 51750
rect 25872 51264 25924 51270
rect 25872 51206 25924 51212
rect 25884 41818 25912 51206
rect 25872 41812 25924 41818
rect 25872 41754 25924 41760
rect 25780 40724 25832 40730
rect 25780 40666 25832 40672
rect 25686 40080 25742 40089
rect 25686 40015 25742 40024
rect 25412 39024 25464 39030
rect 25412 38966 25464 38972
rect 25320 38956 25372 38962
rect 25320 38898 25372 38904
rect 25136 38752 25188 38758
rect 25136 38694 25188 38700
rect 24952 38412 25004 38418
rect 24952 38354 25004 38360
rect 25044 37392 25096 37398
rect 25044 37334 25096 37340
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 25056 33658 25084 37334
rect 25148 36378 25176 38694
rect 25332 38321 25360 38898
rect 25976 38554 26004 53518
rect 25964 38548 26016 38554
rect 25964 38490 26016 38496
rect 25318 38312 25374 38321
rect 25318 38247 25374 38256
rect 25318 37496 25374 37505
rect 25318 37431 25374 37440
rect 25332 37262 25360 37431
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 25320 37120 25372 37126
rect 25320 37062 25372 37068
rect 25332 36786 25360 37062
rect 25320 36780 25372 36786
rect 25320 36722 25372 36728
rect 25332 36689 25360 36722
rect 25318 36680 25374 36689
rect 25318 36615 25374 36624
rect 25136 36372 25188 36378
rect 25136 36314 25188 36320
rect 25320 36168 25372 36174
rect 25320 36110 25372 36116
rect 25332 35873 25360 36110
rect 25318 35864 25374 35873
rect 25318 35799 25374 35808
rect 25228 35760 25280 35766
rect 25228 35702 25280 35708
rect 25240 35494 25268 35702
rect 25228 35488 25280 35494
rect 25228 35430 25280 35436
rect 25320 35488 25372 35494
rect 25320 35430 25372 35436
rect 25240 35018 25268 35430
rect 25332 35086 25360 35430
rect 25320 35080 25372 35086
rect 25318 35048 25320 35057
rect 25372 35048 25374 35057
rect 25228 35012 25280 35018
rect 25318 34983 25374 34992
rect 25228 34954 25280 34960
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25332 34241 25360 34546
rect 25318 34232 25374 34241
rect 25318 34167 25320 34176
rect 25372 34167 25374 34176
rect 25320 34138 25372 34144
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 25410 33416 25466 33425
rect 25410 33351 25466 33360
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 25332 32609 25360 32846
rect 25318 32600 25374 32609
rect 25318 32535 25374 32544
rect 25424 32434 25452 33351
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25134 32328 25190 32337
rect 25134 32263 25136 32272
rect 25188 32263 25190 32272
rect 25136 32234 25188 32240
rect 25320 31816 25372 31822
rect 25318 31784 25320 31793
rect 25372 31784 25374 31793
rect 25318 31719 25374 31728
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 25332 30977 25360 31282
rect 25318 30968 25374 30977
rect 25318 30903 25320 30912
rect 25372 30903 25374 30912
rect 25320 30874 25372 30880
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 25136 30592 25188 30598
rect 25136 30534 25188 30540
rect 24768 29776 24820 29782
rect 24768 29718 24820 29724
rect 24780 28558 24808 29718
rect 24768 28552 24820 28558
rect 24768 28494 24820 28500
rect 24858 28520 24914 28529
rect 24858 28455 24860 28464
rect 24912 28455 24914 28464
rect 24860 28426 24912 28432
rect 24676 28144 24728 28150
rect 24676 28086 24728 28092
rect 24676 28008 24728 28014
rect 24676 27950 24728 27956
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24492 26444 24544 26450
rect 24492 26386 24544 26392
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 24400 25764 24452 25770
rect 24400 25706 24452 25712
rect 24032 25288 24084 25294
rect 23754 25256 23810 25265
rect 24032 25230 24084 25236
rect 24308 25288 24360 25294
rect 24308 25230 24360 25236
rect 23754 25191 23810 25200
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 23204 23792 23256 23798
rect 23204 23734 23256 23740
rect 23216 23662 23244 23734
rect 23204 23656 23256 23662
rect 23204 23598 23256 23604
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22836 22976 22888 22982
rect 22836 22918 22888 22924
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 22664 22066 22784 22094
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22388 20942 22416 21082
rect 22664 20942 22692 22066
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22388 20806 22416 20878
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22284 19304 22336 19310
rect 22204 19264 22284 19292
rect 22284 19246 22336 19252
rect 22296 18970 22324 19246
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 22296 16046 22324 18906
rect 22388 18630 22416 20742
rect 22560 19440 22612 19446
rect 22560 19382 22612 19388
rect 22572 18850 22600 19382
rect 22848 19310 22876 22918
rect 23296 22772 23348 22778
rect 23296 22714 23348 22720
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 22098 23336 22714
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 23492 21570 23520 22918
rect 23308 21554 23520 21570
rect 23296 21548 23520 21554
rect 23348 21542 23520 21548
rect 23296 21490 23348 21496
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23386 21176 23442 21185
rect 23386 21111 23442 21120
rect 23400 20534 23428 21111
rect 23480 21072 23532 21078
rect 23480 21014 23532 21020
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23294 19544 23350 19553
rect 23294 19479 23350 19488
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22572 18822 22784 18850
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22572 17882 22600 18634
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21836 12714 21864 14214
rect 21824 12708 21876 12714
rect 21824 12650 21876 12656
rect 21836 12306 21864 12650
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 21732 9920 21784 9926
rect 21732 9862 21784 9868
rect 21744 5574 21772 9862
rect 21928 9654 21956 15302
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 22020 12238 22048 13126
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 22008 11620 22060 11626
rect 22008 11562 22060 11568
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 21732 5568 21784 5574
rect 21732 5510 21784 5516
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21744 3466 21772 4626
rect 21732 3460 21784 3466
rect 21732 3402 21784 3408
rect 21836 3398 21864 6666
rect 22020 6322 22048 11562
rect 22112 6914 22140 13806
rect 22204 12306 22232 15846
rect 22388 15162 22416 16050
rect 22572 16046 22600 17818
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22664 16522 22692 16594
rect 22652 16516 22704 16522
rect 22652 16458 22704 16464
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22296 13530 22324 14350
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22112 6886 22232 6914
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21824 3392 21876 3398
rect 21824 3334 21876 3340
rect 21928 800 21956 6190
rect 22204 5234 22232 6886
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22112 4049 22140 4082
rect 22098 4040 22154 4049
rect 22098 3975 22154 3984
rect 22296 800 22324 7278
rect 22388 4146 22416 14010
rect 22480 12850 22508 15846
rect 22664 14414 22692 16458
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22468 9104 22520 9110
rect 22468 9046 22520 9052
rect 22480 7750 22508 9046
rect 22664 8974 22692 14010
rect 22756 13938 22784 18822
rect 22928 18624 22980 18630
rect 22928 18566 22980 18572
rect 22940 18222 22968 18566
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23308 17134 23336 19479
rect 23386 18728 23442 18737
rect 23386 18663 23442 18672
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23400 16046 23428 18663
rect 23492 16114 23520 21014
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23388 16040 23440 16046
rect 23388 15982 23440 15988
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23584 15026 23612 24006
rect 23664 23656 23716 23662
rect 23664 23598 23716 23604
rect 23676 22778 23704 23598
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23664 22636 23716 22642
rect 23664 22578 23716 22584
rect 23676 21622 23704 22578
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23676 17610 23704 18158
rect 23664 17604 23716 17610
rect 23664 17546 23716 17552
rect 23676 16658 23704 17546
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 23664 15972 23716 15978
rect 23664 15914 23716 15920
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 23294 13832 23350 13841
rect 23294 13767 23350 13776
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23308 12850 23336 13767
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22572 7206 22600 8774
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22480 2854 22508 5102
rect 22572 3942 22600 6258
rect 22664 4758 22692 8434
rect 22652 4752 22704 4758
rect 22652 4694 22704 4700
rect 22756 4622 22784 9318
rect 22848 8090 22876 11698
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23386 11384 23442 11393
rect 23386 11319 23442 11328
rect 23296 10464 23348 10470
rect 23296 10406 23348 10412
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23308 8514 23336 10406
rect 23400 9518 23428 11319
rect 23676 10674 23704 15914
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23308 8486 23428 8514
rect 23296 8424 23348 8430
rect 23296 8366 23348 8372
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 22848 6798 22876 7686
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22468 2848 22520 2854
rect 22468 2790 22520 2796
rect 22664 800 22692 3130
rect 22848 2530 22876 3334
rect 23124 3194 23152 3470
rect 23308 3233 23336 8366
rect 23400 7410 23428 8486
rect 23492 7886 23520 8774
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23400 4554 23428 7142
rect 23388 4548 23440 4554
rect 23388 4490 23440 4496
rect 23294 3224 23350 3233
rect 23112 3188 23164 3194
rect 23294 3159 23350 3168
rect 23112 3130 23164 3136
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22848 2502 23060 2530
rect 23032 800 23060 2502
rect 23400 800 23428 2926
rect 23768 800 23796 25191
rect 23940 25152 23992 25158
rect 23940 25094 23992 25100
rect 23846 23624 23902 23633
rect 23846 23559 23902 23568
rect 23860 23186 23888 23559
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 23860 13938 23888 19722
rect 23952 17202 23980 25094
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 24320 23730 24348 24754
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24216 23520 24268 23526
rect 24216 23462 24268 23468
rect 24228 22098 24256 23462
rect 24320 22778 24348 23666
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 24216 22092 24268 22098
rect 24216 22034 24268 22040
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24032 19168 24084 19174
rect 24032 19110 24084 19116
rect 24044 18290 24072 19110
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24044 18086 24072 18226
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 24044 11694 24072 18022
rect 24136 15026 24164 21966
rect 24216 21616 24268 21622
rect 24216 21558 24268 21564
rect 24228 21146 24256 21558
rect 24216 21140 24268 21146
rect 24216 21082 24268 21088
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24228 15502 24256 17478
rect 24412 16182 24440 25706
rect 24504 23662 24532 26386
rect 24688 24750 24716 27950
rect 25148 27062 25176 30534
rect 25318 30152 25374 30161
rect 25318 30087 25374 30096
rect 25332 29646 25360 30087
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25332 29306 25360 29582
rect 25516 29345 25544 30670
rect 25688 29844 25740 29850
rect 25688 29786 25740 29792
rect 25502 29336 25558 29345
rect 25320 29300 25372 29306
rect 25502 29271 25504 29280
rect 25320 29242 25372 29248
rect 25556 29271 25558 29280
rect 25504 29242 25556 29248
rect 25596 27396 25648 27402
rect 25596 27338 25648 27344
rect 25228 27328 25280 27334
rect 25228 27270 25280 27276
rect 25136 27056 25188 27062
rect 25136 26998 25188 27004
rect 25240 26586 25268 27270
rect 25502 26888 25558 26897
rect 25412 26852 25464 26858
rect 25502 26823 25558 26832
rect 25412 26794 25464 26800
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 25228 26580 25280 26586
rect 25228 26522 25280 26528
rect 25056 25498 25084 26522
rect 25228 26308 25280 26314
rect 25228 26250 25280 26256
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 25044 25492 25096 25498
rect 25044 25434 25096 25440
rect 24872 24818 24900 25434
rect 24952 25424 25004 25430
rect 24952 25366 25004 25372
rect 24860 24812 24912 24818
rect 24860 24754 24912 24760
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 24584 24608 24636 24614
rect 24584 24550 24636 24556
rect 24492 23656 24544 23662
rect 24492 23598 24544 23604
rect 24504 23254 24532 23598
rect 24492 23248 24544 23254
rect 24492 23190 24544 23196
rect 24504 22642 24532 23190
rect 24596 23186 24624 24550
rect 24688 24410 24716 24686
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24676 24404 24728 24410
rect 24676 24346 24728 24352
rect 24780 24342 24808 24550
rect 24858 24440 24914 24449
rect 24858 24375 24914 24384
rect 24768 24336 24820 24342
rect 24768 24278 24820 24284
rect 24872 24274 24900 24375
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24964 24206 24992 25366
rect 25148 25265 25176 25774
rect 25134 25256 25190 25265
rect 25044 25220 25096 25226
rect 25134 25191 25190 25200
rect 25044 25162 25096 25168
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24584 23180 24636 23186
rect 24584 23122 24636 23128
rect 24674 22808 24730 22817
rect 24674 22743 24730 22752
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 24688 20398 24716 22743
rect 25056 22094 25084 25162
rect 25056 22066 25176 22094
rect 24858 21992 24914 22001
rect 24858 21927 24914 21936
rect 24872 21010 24900 21927
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 25044 20868 25096 20874
rect 25044 20810 25096 20816
rect 24676 20392 24728 20398
rect 24676 20334 24728 20340
rect 24950 20360 25006 20369
rect 24950 20295 25006 20304
rect 24964 19922 24992 20295
rect 24952 19916 25004 19922
rect 24952 19858 25004 19864
rect 24858 17912 24914 17921
rect 24858 17847 24914 17856
rect 24872 17270 24900 17847
rect 25056 17678 25084 20810
rect 25148 20534 25176 22066
rect 25136 20528 25188 20534
rect 25136 20470 25188 20476
rect 25240 20466 25268 26250
rect 25318 26072 25374 26081
rect 25318 26007 25374 26016
rect 25332 23730 25360 26007
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 25332 22778 25360 23666
rect 25424 23050 25452 26794
rect 25516 25498 25544 26823
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 25516 24818 25544 25434
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25412 23044 25464 23050
rect 25412 22986 25464 22992
rect 25320 22772 25372 22778
rect 25320 22714 25372 22720
rect 25228 20460 25280 20466
rect 25228 20402 25280 20408
rect 25608 19854 25636 27338
rect 25700 24206 25728 29786
rect 25688 24200 25740 24206
rect 25688 24142 25740 24148
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 24860 17264 24912 17270
rect 24860 17206 24912 17212
rect 24766 17096 24822 17105
rect 24766 17031 24822 17040
rect 24674 16280 24730 16289
rect 24674 16215 24730 16224
rect 24400 16176 24452 16182
rect 24400 16118 24452 16124
rect 24216 15496 24268 15502
rect 24216 15438 24268 15444
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24688 13870 24716 16215
rect 24780 14958 24808 17031
rect 24950 15464 25006 15473
rect 24950 15399 24952 15408
rect 25004 15399 25006 15408
rect 24952 15370 25004 15376
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24766 14648 24822 14657
rect 24766 14583 24822 14592
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24780 12782 24808 14583
rect 25504 13252 25556 13258
rect 25504 13194 25556 13200
rect 25516 13025 25544 13194
rect 25502 13016 25558 13025
rect 25502 12951 25558 12960
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24860 12368 24912 12374
rect 24860 12310 24912 12316
rect 24766 12200 24822 12209
rect 24766 12135 24822 12144
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 23952 8498 23980 11018
rect 24780 10606 24808 12135
rect 24768 10600 24820 10606
rect 24674 10568 24730 10577
rect 24768 10542 24820 10548
rect 24674 10503 24730 10512
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 24044 5234 24072 9862
rect 24688 8430 24716 10503
rect 24872 8974 24900 12310
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24964 9761 24992 9998
rect 24950 9752 25006 9761
rect 24950 9687 25006 9696
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 24766 8120 24822 8129
rect 24766 8055 24822 8064
rect 24492 7812 24544 7818
rect 24492 7754 24544 7760
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 24504 4865 24532 7754
rect 24674 7304 24730 7313
rect 24674 7239 24730 7248
rect 24688 6746 24716 7239
rect 24596 6718 24716 6746
rect 24596 5166 24624 6718
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24584 5160 24636 5166
rect 24584 5102 24636 5108
rect 24490 4856 24546 4865
rect 24490 4791 24546 4800
rect 24688 4146 24716 6598
rect 24780 6254 24808 8055
rect 24860 7880 24912 7886
rect 24860 7822 24912 7828
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24766 5672 24822 5681
rect 24766 5607 24822 5616
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24780 4078 24808 5607
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24124 2848 24176 2854
rect 24124 2790 24176 2796
rect 24136 800 24164 2790
rect 24596 2446 24624 3334
rect 24872 3194 24900 7822
rect 25056 6914 25084 12038
rect 25134 8936 25190 8945
rect 25134 8871 25190 8880
rect 25148 7478 25176 8871
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 24964 6886 25084 6914
rect 24964 6798 24992 6886
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 25056 6497 25084 6666
rect 25042 6488 25098 6497
rect 25042 6423 25098 6432
rect 24952 4004 25004 4010
rect 24952 3946 25004 3952
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24872 1601 24900 2450
rect 24858 1592 24914 1601
rect 24858 1527 24914 1536
rect 13188 734 13400 762
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 24964 785 24992 3946
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 25332 2650 25360 2994
rect 25320 2644 25372 2650
rect 25320 2586 25372 2592
rect 24950 776 25006 785
rect 24950 711 25006 720
<< via2 >>
rect 1306 52944 1362 53000
rect 1306 50496 1362 50552
rect 2226 53524 2228 53544
rect 2228 53524 2280 53544
rect 2280 53524 2282 53544
rect 2226 53488 2282 53524
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 3974 55392 4030 55448
rect 1306 48068 1362 48104
rect 1306 48048 1308 48068
rect 1308 48048 1360 48068
rect 1360 48048 1362 48068
rect 1306 45620 1362 45656
rect 1306 45600 1308 45620
rect 1308 45600 1360 45620
rect 1360 45600 1362 45620
rect 1214 43152 1270 43208
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 1306 40704 1362 40760
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 1306 38292 1308 38312
rect 1308 38292 1360 38312
rect 1360 38292 1362 38312
rect 1306 38256 1362 38292
rect 1582 35808 1638 35864
rect 1214 33360 1270 33416
rect 1306 30912 1362 30968
rect 1306 28464 1362 28520
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 1306 23604 1308 23624
rect 1308 23604 1360 23624
rect 1360 23604 1362 23624
rect 1306 23568 1362 23604
rect 2778 26016 2834 26072
rect 4434 40704 4490 40760
rect 7378 53488 7434 53544
rect 5446 32444 5448 32464
rect 5448 32444 5500 32464
rect 5500 32444 5502 32464
rect 5446 32408 5502 32444
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7378 39888 7434 39944
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 8206 38256 8262 38312
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 1306 21120 1362 21176
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 1306 18672 1362 18728
rect 1306 16224 1362 16280
rect 1306 13812 1308 13832
rect 1308 13812 1360 13832
rect 1360 13812 1362 13832
rect 1306 13776 1362 13812
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2502 16496 2558 16552
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3606 8880 3662 8936
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3422 1536 3478 1592
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 8482 40724 8538 40760
rect 8482 40704 8484 40724
rect 8484 40704 8536 40724
rect 8536 40704 8538 40724
rect 8574 36080 8630 36136
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 8666 35808 8722 35864
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 8850 38528 8906 38584
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 4066 16496 4122 16552
rect 3882 11600 3938 11656
rect 4066 6432 4122 6488
rect 3790 5752 3846 5808
rect 4986 18128 5042 18184
rect 3698 3984 3754 4040
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 9586 40432 9642 40488
rect 10322 42508 10324 42528
rect 10324 42508 10376 42528
rect 10376 42508 10378 42528
rect 10322 42472 10378 42508
rect 9770 36760 9826 36816
rect 10230 37712 10286 37768
rect 9954 36760 10010 36816
rect 9770 31884 9826 31920
rect 9770 31864 9772 31884
rect 9772 31864 9824 31884
rect 9824 31864 9826 31884
rect 11610 44260 11666 44296
rect 11610 44240 11612 44260
rect 11612 44240 11664 44260
rect 11664 44240 11666 44260
rect 11242 40432 11298 40488
rect 10506 37712 10562 37768
rect 11978 40468 11980 40488
rect 11980 40468 12032 40488
rect 12032 40468 12034 40488
rect 11610 38256 11666 38312
rect 8666 19660 8668 19680
rect 8668 19660 8720 19680
rect 8720 19660 8722 19680
rect 8666 19624 8722 19660
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 9494 16496 9550 16552
rect 8482 5616 8538 5672
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 9586 5072 9642 5128
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 11426 30676 11428 30696
rect 11428 30676 11480 30696
rect 11480 30676 11482 30696
rect 11426 30640 11482 30676
rect 11978 40432 12034 40468
rect 12070 37304 12126 37360
rect 11610 32972 11666 33008
rect 11610 32952 11612 32972
rect 11612 32952 11664 32972
rect 11664 32952 11666 32972
rect 11058 23976 11114 24032
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12530 37848 12586 37904
rect 12438 35808 12494 35864
rect 12254 32308 12256 32328
rect 12256 32308 12308 32328
rect 12308 32308 12310 32328
rect 12254 32272 12310 32308
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 13266 38412 13322 38448
rect 13266 38392 13268 38412
rect 13268 38392 13320 38412
rect 13320 38392 13322 38412
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12530 33260 12532 33280
rect 12532 33260 12584 33280
rect 12584 33260 12586 33280
rect 12530 33224 12586 33260
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 11886 23976 11942 24032
rect 12162 19372 12218 19408
rect 12162 19352 12164 19372
rect 12164 19352 12216 19372
rect 12216 19352 12218 19372
rect 13818 38256 13874 38312
rect 13818 36252 13820 36272
rect 13820 36252 13872 36272
rect 13872 36252 13874 36272
rect 13818 36216 13874 36252
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12530 17876 12586 17912
rect 12530 17856 12532 17876
rect 12532 17856 12584 17876
rect 12584 17856 12586 17876
rect 14002 32408 14058 32464
rect 14278 38528 14334 38584
rect 15198 37324 15254 37360
rect 15198 37304 15200 37324
rect 15200 37304 15252 37324
rect 15252 37304 15254 37324
rect 13542 21956 13598 21992
rect 13542 21936 13544 21956
rect 13544 21936 13596 21956
rect 13596 21936 13598 21956
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12898 18264 12954 18320
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 15474 36896 15530 36952
rect 15658 36100 15714 36136
rect 15658 36080 15660 36100
rect 15660 36080 15712 36100
rect 15712 36080 15714 36100
rect 16394 52536 16450 52592
rect 15842 43052 15844 43072
rect 15844 43052 15896 43072
rect 15896 43052 15898 43072
rect 15842 43016 15898 43052
rect 16026 38700 16028 38720
rect 16028 38700 16080 38720
rect 16080 38700 16082 38720
rect 16026 38664 16082 38700
rect 15842 36660 15844 36680
rect 15844 36660 15896 36680
rect 15896 36660 15898 36680
rect 15842 36624 15898 36660
rect 16118 38004 16174 38040
rect 16118 37984 16120 38004
rect 16120 37984 16172 38004
rect 16172 37984 16174 38004
rect 14738 28328 14794 28384
rect 13542 14048 13598 14104
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 14646 21664 14702 21720
rect 15290 28192 15346 28248
rect 15382 27240 15438 27296
rect 14738 19660 14740 19680
rect 14740 19660 14792 19680
rect 14792 19660 14794 19680
rect 14738 19624 14794 19660
rect 16670 36780 16726 36816
rect 16670 36760 16672 36780
rect 16672 36760 16724 36780
rect 16724 36760 16726 36780
rect 17130 52536 17186 52592
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 24582 56208 24638 56264
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 16854 40024 16910 40080
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 18510 47640 18566 47696
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17130 39888 17186 39944
rect 17314 38528 17370 38584
rect 16578 32408 16634 32464
rect 16118 29144 16174 29200
rect 14738 16244 14794 16280
rect 14738 16224 14740 16244
rect 14740 16224 14792 16244
rect 14792 16224 14794 16244
rect 15934 28212 15990 28248
rect 15934 28192 15936 28212
rect 15936 28192 15988 28212
rect 15988 28192 15990 28212
rect 16394 29028 16450 29064
rect 16394 29008 16396 29028
rect 16396 29008 16448 29028
rect 16448 29008 16450 29028
rect 16026 27956 16028 27976
rect 16028 27956 16080 27976
rect 16080 27956 16082 27976
rect 16026 27920 16082 27956
rect 16762 28364 16764 28384
rect 16764 28364 16816 28384
rect 16816 28364 16818 28384
rect 16762 28328 16818 28364
rect 16118 20712 16174 20768
rect 15934 16224 15990 16280
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 18234 40024 18290 40080
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 18418 38836 18420 38856
rect 18420 38836 18472 38856
rect 18472 38836 18474 38856
rect 18418 38800 18474 38836
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 20074 45908 20076 45928
rect 20076 45908 20128 45928
rect 20128 45908 20130 45928
rect 20074 45872 20130 45908
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17406 31864 17462 31920
rect 17130 27376 17186 27432
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 18234 31728 18290 31784
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 18050 30232 18106 30288
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 18326 28464 18382 28520
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 16670 18264 16726 18320
rect 16302 16768 16358 16824
rect 17314 20596 17370 20632
rect 17314 20576 17316 20596
rect 17316 20576 17368 20596
rect 17368 20576 17370 20596
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 19614 39480 19670 39536
rect 18694 30252 18750 30288
rect 18694 30232 18696 30252
rect 18696 30232 18748 30252
rect 18748 30232 18750 30252
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17774 19896 17830 19952
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18510 20576 18566 20632
rect 18418 19352 18474 19408
rect 18326 18672 18382 18728
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 19982 40296 20038 40352
rect 19430 31900 19432 31920
rect 19432 31900 19484 31920
rect 19484 31900 19486 31920
rect 19430 31864 19486 31900
rect 20442 40024 20498 40080
rect 20258 39480 20314 39536
rect 20258 37868 20314 37904
rect 20258 37848 20260 37868
rect 20260 37848 20312 37868
rect 20312 37848 20314 37868
rect 19890 35400 19946 35456
rect 19982 32000 20038 32056
rect 19982 31220 19984 31240
rect 19984 31220 20036 31240
rect 20036 31220 20038 31240
rect 19982 31184 20038 31220
rect 19890 30796 19946 30832
rect 19890 30776 19892 30796
rect 19892 30776 19944 30796
rect 19944 30776 19946 30796
rect 20258 33532 20260 33552
rect 20260 33532 20312 33552
rect 20312 33532 20314 33552
rect 20258 33496 20314 33532
rect 20166 32272 20222 32328
rect 20166 29044 20168 29064
rect 20168 29044 20220 29064
rect 20220 29044 20222 29064
rect 20166 29008 20222 29044
rect 20074 28328 20130 28384
rect 19154 20712 19210 20768
rect 20074 27820 20076 27840
rect 20076 27820 20128 27840
rect 20128 27820 20130 27840
rect 20074 27784 20130 27820
rect 21638 46996 21640 47016
rect 21640 46996 21692 47016
rect 21692 46996 21694 47016
rect 21638 46960 21694 46996
rect 21638 43052 21640 43072
rect 21640 43052 21692 43072
rect 21692 43052 21694 43072
rect 21638 43016 21694 43052
rect 20534 32000 20590 32056
rect 21362 39888 21418 39944
rect 21914 45908 21916 45928
rect 21916 45908 21968 45928
rect 21968 45908 21970 45928
rect 21914 45872 21970 45908
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 23662 52536 23718 52592
rect 22558 46552 22614 46608
rect 22374 43288 22430 43344
rect 22650 43288 22706 43344
rect 21362 33496 21418 33552
rect 21362 32952 21418 33008
rect 21270 32680 21326 32736
rect 22466 40024 22522 40080
rect 22282 36624 22338 36680
rect 21914 32716 21916 32736
rect 21916 32716 21968 32736
rect 21968 32716 21970 32736
rect 21914 32680 21970 32716
rect 21914 32564 21970 32600
rect 21914 32544 21916 32564
rect 21916 32544 21968 32564
rect 21968 32544 21970 32564
rect 21546 29180 21548 29200
rect 21548 29180 21600 29200
rect 21600 29180 21602 29200
rect 21546 29144 21602 29180
rect 19982 20712 20038 20768
rect 20258 20712 20314 20768
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18694 3984 18750 4040
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 23294 39208 23350 39264
rect 22558 35400 22614 35456
rect 22374 33088 22430 33144
rect 22466 32952 22522 33008
rect 22374 32680 22430 32736
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 23846 41248 23902 41304
rect 24674 55392 24730 55448
rect 24766 54576 24822 54632
rect 24674 53760 24730 53816
rect 25042 52944 25098 53000
rect 24766 52128 24822 52184
rect 23938 39888 23994 39944
rect 23846 39208 23902 39264
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 24766 46416 24822 46472
rect 24858 45600 24914 45656
rect 25042 51348 25044 51368
rect 25044 51348 25096 51368
rect 25096 51348 25098 51368
rect 25042 51312 25098 51348
rect 25042 50496 25098 50552
rect 25318 49680 25374 49736
rect 25318 48864 25374 48920
rect 25318 48084 25320 48104
rect 25320 48084 25372 48104
rect 25372 48084 25374 48104
rect 25318 48048 25374 48084
rect 24490 41248 24546 41304
rect 24582 40332 24584 40352
rect 24584 40332 24636 40352
rect 24636 40332 24638 40352
rect 24582 40296 24638 40332
rect 24766 43152 24822 43208
rect 25318 43152 25374 43208
rect 24858 42336 24914 42392
rect 24766 39888 24822 39944
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 21362 2352 21418 2408
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 24122 27648 24178 27704
rect 24858 39072 24914 39128
rect 25318 41556 25320 41576
rect 25320 41556 25372 41576
rect 25372 41556 25374 41576
rect 25318 41520 25374 41556
rect 25318 40704 25374 40760
rect 25502 47232 25558 47288
rect 25502 44784 25558 44840
rect 25502 43968 25558 44024
rect 25686 40024 25742 40080
rect 25318 38256 25374 38312
rect 25318 37440 25374 37496
rect 25318 36624 25374 36680
rect 25318 35808 25374 35864
rect 25318 35028 25320 35048
rect 25320 35028 25372 35048
rect 25372 35028 25374 35048
rect 25318 34992 25374 35028
rect 25318 34196 25374 34232
rect 25318 34176 25320 34196
rect 25320 34176 25372 34196
rect 25372 34176 25374 34196
rect 25410 33360 25466 33416
rect 25318 32544 25374 32600
rect 25134 32292 25190 32328
rect 25134 32272 25136 32292
rect 25136 32272 25188 32292
rect 25188 32272 25190 32292
rect 25318 31764 25320 31784
rect 25320 31764 25372 31784
rect 25372 31764 25374 31784
rect 25318 31728 25374 31764
rect 25318 30932 25374 30968
rect 25318 30912 25320 30932
rect 25320 30912 25372 30932
rect 25372 30912 25374 30932
rect 24858 28484 24914 28520
rect 24858 28464 24860 28484
rect 24860 28464 24912 28484
rect 24912 28464 24914 28484
rect 23754 25200 23810 25256
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23386 21120 23442 21176
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 23294 19488 23350 19544
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22098 3984 22154 4040
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23386 18672 23442 18728
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 23294 13776 23350 13832
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 23386 11328 23442 11384
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 23294 3168 23350 3224
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 23846 23568 23902 23624
rect 25318 30096 25374 30152
rect 25502 29300 25558 29336
rect 25502 29280 25504 29300
rect 25504 29280 25556 29300
rect 25556 29280 25558 29300
rect 25502 26832 25558 26888
rect 24858 24384 24914 24440
rect 25134 25200 25190 25256
rect 24674 22752 24730 22808
rect 24858 21936 24914 21992
rect 24950 20304 25006 20360
rect 24858 17856 24914 17912
rect 25318 26016 25374 26072
rect 24766 17040 24822 17096
rect 24674 16224 24730 16280
rect 24950 15428 25006 15464
rect 24950 15408 24952 15428
rect 24952 15408 25004 15428
rect 25004 15408 25006 15428
rect 24766 14592 24822 14648
rect 25502 12960 25558 13016
rect 24766 12144 24822 12200
rect 24674 10512 24730 10568
rect 24950 9696 25006 9752
rect 24766 8064 24822 8120
rect 24674 7248 24730 7304
rect 24490 4800 24546 4856
rect 24766 5616 24822 5672
rect 25134 8880 25190 8936
rect 25042 6432 25098 6488
rect 24858 1536 24914 1592
rect 24950 720 25006 776
<< metal3 >>
rect 24577 56266 24643 56269
rect 26200 56266 27000 56296
rect 24577 56264 27000 56266
rect 24577 56208 24582 56264
rect 24638 56208 27000 56264
rect 24577 56206 27000 56208
rect 24577 56203 24643 56206
rect 26200 56176 27000 56206
rect 0 55450 800 55480
rect 3969 55450 4035 55453
rect 0 55448 4035 55450
rect 0 55392 3974 55448
rect 4030 55392 4035 55448
rect 0 55390 4035 55392
rect 0 55360 800 55390
rect 3969 55387 4035 55390
rect 24669 55450 24735 55453
rect 26200 55450 27000 55480
rect 24669 55448 27000 55450
rect 24669 55392 24674 55448
rect 24730 55392 27000 55448
rect 24669 55390 27000 55392
rect 24669 55387 24735 55390
rect 26200 55360 27000 55390
rect 24761 54634 24827 54637
rect 26200 54634 27000 54664
rect 24761 54632 27000 54634
rect 24761 54576 24766 54632
rect 24822 54576 27000 54632
rect 24761 54574 27000 54576
rect 24761 54571 24827 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 24669 53818 24735 53821
rect 26200 53818 27000 53848
rect 24669 53816 27000 53818
rect 24669 53760 24674 53816
rect 24730 53760 27000 53816
rect 24669 53758 27000 53760
rect 24669 53755 24735 53758
rect 26200 53728 27000 53758
rect 2221 53546 2287 53549
rect 7373 53546 7439 53549
rect 2221 53544 7439 53546
rect 2221 53488 2226 53544
rect 2282 53488 7378 53544
rect 7434 53488 7439 53544
rect 2221 53486 7439 53488
rect 2221 53483 2287 53486
rect 7373 53483 7439 53486
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 0 53002 800 53032
rect 1301 53002 1367 53005
rect 0 53000 1367 53002
rect 0 52944 1306 53000
rect 1362 52944 1367 53000
rect 0 52942 1367 52944
rect 0 52912 800 52942
rect 1301 52939 1367 52942
rect 25037 53002 25103 53005
rect 26200 53002 27000 53032
rect 25037 53000 27000 53002
rect 25037 52944 25042 53000
rect 25098 52944 27000 53000
rect 25037 52942 27000 52944
rect 25037 52939 25103 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 16389 52596 16455 52597
rect 17125 52596 17191 52597
rect 16389 52592 16436 52596
rect 16500 52594 16506 52596
rect 16389 52536 16394 52592
rect 16389 52532 16436 52536
rect 16500 52534 16546 52594
rect 17125 52592 17172 52596
rect 17236 52594 17242 52596
rect 23657 52594 23723 52597
rect 23790 52594 23796 52596
rect 17125 52536 17130 52592
rect 16500 52532 16506 52534
rect 17125 52532 17172 52536
rect 17236 52534 17282 52594
rect 23657 52592 23796 52594
rect 23657 52536 23662 52592
rect 23718 52536 23796 52592
rect 23657 52534 23796 52536
rect 17236 52532 17242 52534
rect 16389 52531 16455 52532
rect 17125 52531 17191 52532
rect 23657 52531 23723 52534
rect 23790 52532 23796 52534
rect 23860 52532 23866 52596
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 24761 52186 24827 52189
rect 26200 52186 27000 52216
rect 24761 52184 27000 52186
rect 24761 52128 24766 52184
rect 24822 52128 27000 52184
rect 24761 52126 27000 52128
rect 24761 52123 24827 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 25037 51370 25103 51373
rect 26200 51370 27000 51400
rect 25037 51368 27000 51370
rect 25037 51312 25042 51368
rect 25098 51312 27000 51368
rect 25037 51310 27000 51312
rect 25037 51307 25103 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 0 50554 800 50584
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 1301 50554 1367 50557
rect 0 50552 1367 50554
rect 0 50496 1306 50552
rect 1362 50496 1367 50552
rect 0 50494 1367 50496
rect 0 50464 800 50494
rect 1301 50491 1367 50494
rect 25037 50554 25103 50557
rect 26200 50554 27000 50584
rect 25037 50552 27000 50554
rect 25037 50496 25042 50552
rect 25098 50496 27000 50552
rect 25037 50494 27000 50496
rect 25037 50491 25103 50494
rect 26200 50464 27000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25313 49738 25379 49741
rect 26200 49738 27000 49768
rect 25313 49736 27000 49738
rect 25313 49680 25318 49736
rect 25374 49680 27000 49736
rect 25313 49678 27000 49680
rect 25313 49675 25379 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25313 48922 25379 48925
rect 26200 48922 27000 48952
rect 25313 48920 27000 48922
rect 25313 48864 25318 48920
rect 25374 48864 27000 48920
rect 25313 48862 27000 48864
rect 25313 48859 25379 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 0 48106 800 48136
rect 1301 48106 1367 48109
rect 0 48104 1367 48106
rect 0 48048 1306 48104
rect 1362 48048 1367 48104
rect 0 48046 1367 48048
rect 0 48016 800 48046
rect 1301 48043 1367 48046
rect 25313 48106 25379 48109
rect 26200 48106 27000 48136
rect 25313 48104 27000 48106
rect 25313 48048 25318 48104
rect 25374 48048 27000 48104
rect 25313 48046 27000 48048
rect 25313 48043 25379 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 18505 47698 18571 47701
rect 18638 47698 18644 47700
rect 18505 47696 18644 47698
rect 18505 47640 18510 47696
rect 18566 47640 18644 47696
rect 18505 47638 18644 47640
rect 18505 47635 18571 47638
rect 18638 47636 18644 47638
rect 18708 47636 18714 47700
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25497 47290 25563 47293
rect 26200 47290 27000 47320
rect 25497 47288 27000 47290
rect 25497 47232 25502 47288
rect 25558 47232 27000 47288
rect 25497 47230 27000 47232
rect 25497 47227 25563 47230
rect 26200 47200 27000 47230
rect 21633 47018 21699 47021
rect 21766 47018 21772 47020
rect 21633 47016 21772 47018
rect 21633 46960 21638 47016
rect 21694 46960 21772 47016
rect 21633 46958 21772 46960
rect 21633 46955 21699 46958
rect 21766 46956 21772 46958
rect 21836 46956 21842 47020
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 22553 46610 22619 46613
rect 22686 46610 22692 46612
rect 22553 46608 22692 46610
rect 22553 46552 22558 46608
rect 22614 46552 22692 46608
rect 22553 46550 22692 46552
rect 22553 46547 22619 46550
rect 22686 46548 22692 46550
rect 22756 46548 22762 46612
rect 24761 46474 24827 46477
rect 26200 46474 27000 46504
rect 24761 46472 27000 46474
rect 24761 46416 24766 46472
rect 24822 46416 27000 46472
rect 24761 46414 27000 46416
rect 24761 46411 24827 46414
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 20069 45932 20135 45933
rect 21909 45932 21975 45933
rect 20069 45928 20116 45932
rect 20180 45930 20186 45932
rect 20069 45872 20074 45928
rect 20069 45868 20116 45872
rect 20180 45870 20226 45930
rect 21909 45928 21956 45932
rect 22020 45930 22026 45932
rect 21909 45872 21914 45928
rect 20180 45868 20186 45870
rect 21909 45868 21956 45872
rect 22020 45870 22066 45930
rect 22020 45868 22026 45870
rect 20069 45867 20135 45868
rect 21909 45867 21975 45868
rect 7946 45728 8262 45729
rect 0 45658 800 45688
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 1301 45658 1367 45661
rect 0 45656 1367 45658
rect 0 45600 1306 45656
rect 1362 45600 1367 45656
rect 0 45598 1367 45600
rect 0 45568 800 45598
rect 1301 45595 1367 45598
rect 24853 45658 24919 45661
rect 26200 45658 27000 45688
rect 24853 45656 27000 45658
rect 24853 45600 24858 45656
rect 24914 45600 27000 45656
rect 24853 45598 27000 45600
rect 24853 45595 24919 45598
rect 26200 45568 27000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 25497 44842 25563 44845
rect 26200 44842 27000 44872
rect 25497 44840 27000 44842
rect 25497 44784 25502 44840
rect 25558 44784 27000 44840
rect 25497 44782 27000 44784
rect 25497 44779 25563 44782
rect 26200 44752 27000 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 11605 44300 11671 44301
rect 11605 44298 11652 44300
rect 11560 44296 11652 44298
rect 11560 44240 11610 44296
rect 11560 44238 11652 44240
rect 11605 44236 11652 44238
rect 11716 44236 11722 44300
rect 11605 44235 11671 44236
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 25497 44026 25563 44029
rect 26200 44026 27000 44056
rect 25497 44024 27000 44026
rect 25497 43968 25502 44024
rect 25558 43968 27000 44024
rect 25497 43966 27000 43968
rect 25497 43963 25563 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 22369 43346 22435 43349
rect 22645 43346 22711 43349
rect 22369 43344 22711 43346
rect 22369 43288 22374 43344
rect 22430 43288 22650 43344
rect 22706 43288 22711 43344
rect 22369 43286 22711 43288
rect 22369 43283 22435 43286
rect 22645 43283 22711 43286
rect 0 43210 800 43240
rect 1209 43210 1275 43213
rect 0 43208 1275 43210
rect 0 43152 1214 43208
rect 1270 43152 1275 43208
rect 0 43150 1275 43152
rect 0 43120 800 43150
rect 1209 43147 1275 43150
rect 19742 43148 19748 43212
rect 19812 43210 19818 43212
rect 24761 43210 24827 43213
rect 19812 43208 24827 43210
rect 19812 43152 24766 43208
rect 24822 43152 24827 43208
rect 19812 43150 24827 43152
rect 19812 43148 19818 43150
rect 24761 43147 24827 43150
rect 25313 43210 25379 43213
rect 26200 43210 27000 43240
rect 25313 43208 27000 43210
rect 25313 43152 25318 43208
rect 25374 43152 27000 43208
rect 25313 43150 27000 43152
rect 25313 43147 25379 43150
rect 26200 43120 27000 43150
rect 15837 43074 15903 43077
rect 21633 43076 21699 43077
rect 16062 43074 16068 43076
rect 15837 43072 16068 43074
rect 15837 43016 15842 43072
rect 15898 43016 16068 43072
rect 15837 43014 16068 43016
rect 15837 43011 15903 43014
rect 16062 43012 16068 43014
rect 16132 43012 16138 43076
rect 21582 43012 21588 43076
rect 21652 43074 21699 43076
rect 21652 43072 21744 43074
rect 21694 43016 21744 43072
rect 21652 43014 21744 43016
rect 21652 43012 21699 43014
rect 21633 43011 21699 43012
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 10317 42530 10383 42533
rect 10910 42530 10916 42532
rect 10317 42528 10916 42530
rect 10317 42472 10322 42528
rect 10378 42472 10916 42528
rect 10317 42470 10916 42472
rect 10317 42467 10383 42470
rect 10910 42468 10916 42470
rect 10980 42468 10986 42532
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 24853 42394 24919 42397
rect 26200 42394 27000 42424
rect 24853 42392 27000 42394
rect 24853 42336 24858 42392
rect 24914 42336 27000 42392
rect 24853 42334 27000 42336
rect 24853 42331 24919 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 25313 41578 25379 41581
rect 26200 41578 27000 41608
rect 25313 41576 27000 41578
rect 25313 41520 25318 41576
rect 25374 41520 27000 41576
rect 25313 41518 27000 41520
rect 25313 41515 25379 41518
rect 26200 41488 27000 41518
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 23841 41306 23907 41309
rect 24485 41306 24551 41309
rect 23841 41304 24551 41306
rect 23841 41248 23846 41304
rect 23902 41248 24490 41304
rect 24546 41248 24551 41304
rect 23841 41246 24551 41248
rect 23841 41243 23907 41246
rect 24485 41243 24551 41246
rect 2946 40832 3262 40833
rect 0 40762 800 40792
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 1301 40762 1367 40765
rect 0 40760 1367 40762
rect 0 40704 1306 40760
rect 1362 40704 1367 40760
rect 0 40702 1367 40704
rect 0 40672 800 40702
rect 1301 40699 1367 40702
rect 4429 40762 4495 40765
rect 8477 40762 8543 40765
rect 4429 40760 8543 40762
rect 4429 40704 4434 40760
rect 4490 40704 8482 40760
rect 8538 40704 8543 40760
rect 4429 40702 8543 40704
rect 4429 40699 4495 40702
rect 8477 40699 8543 40702
rect 25313 40762 25379 40765
rect 26200 40762 27000 40792
rect 25313 40760 27000 40762
rect 25313 40704 25318 40760
rect 25374 40704 27000 40760
rect 25313 40702 27000 40704
rect 25313 40699 25379 40702
rect 26200 40672 27000 40702
rect 9581 40490 9647 40493
rect 11237 40490 11303 40493
rect 11973 40490 12039 40493
rect 9581 40488 12039 40490
rect 9581 40432 9586 40488
rect 9642 40432 11242 40488
rect 11298 40432 11978 40488
rect 12034 40432 12039 40488
rect 9581 40430 12039 40432
rect 9581 40427 9647 40430
rect 11237 40427 11303 40430
rect 11973 40427 12039 40430
rect 19977 40354 20043 40357
rect 24577 40354 24643 40357
rect 19977 40352 24643 40354
rect 19977 40296 19982 40352
rect 20038 40296 24582 40352
rect 24638 40296 24643 40352
rect 19977 40294 24643 40296
rect 19977 40291 20043 40294
rect 24577 40291 24643 40294
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 15878 40020 15884 40084
rect 15948 40082 15954 40084
rect 16849 40082 16915 40085
rect 15948 40080 16915 40082
rect 15948 40024 16854 40080
rect 16910 40024 16915 40080
rect 15948 40022 16915 40024
rect 15948 40020 15954 40022
rect 16849 40019 16915 40022
rect 18229 40082 18295 40085
rect 19190 40082 19196 40084
rect 18229 40080 19196 40082
rect 18229 40024 18234 40080
rect 18290 40024 19196 40080
rect 18229 40022 19196 40024
rect 18229 40019 18295 40022
rect 19190 40020 19196 40022
rect 19260 40020 19266 40084
rect 20437 40082 20503 40085
rect 22461 40082 22527 40085
rect 25681 40082 25747 40085
rect 20437 40080 25747 40082
rect 20437 40024 20442 40080
rect 20498 40024 22466 40080
rect 22522 40024 25686 40080
rect 25742 40024 25747 40080
rect 20437 40022 25747 40024
rect 20437 40019 20503 40022
rect 22461 40019 22527 40022
rect 25681 40019 25747 40022
rect 7373 39946 7439 39949
rect 12198 39946 12204 39948
rect 7373 39944 12204 39946
rect 7373 39888 7378 39944
rect 7434 39888 12204 39944
rect 7373 39886 12204 39888
rect 7373 39883 7439 39886
rect 12198 39884 12204 39886
rect 12268 39884 12274 39948
rect 17125 39946 17191 39949
rect 17350 39946 17356 39948
rect 17125 39944 17356 39946
rect 17125 39888 17130 39944
rect 17186 39888 17356 39944
rect 17125 39886 17356 39888
rect 17125 39883 17191 39886
rect 17350 39884 17356 39886
rect 17420 39884 17426 39948
rect 21357 39946 21423 39949
rect 23933 39946 23999 39949
rect 21357 39944 23999 39946
rect 21357 39888 21362 39944
rect 21418 39888 23938 39944
rect 23994 39888 23999 39944
rect 21357 39886 23999 39888
rect 21357 39883 21423 39886
rect 23933 39883 23999 39886
rect 24761 39946 24827 39949
rect 26200 39946 27000 39976
rect 24761 39944 27000 39946
rect 24761 39888 24766 39944
rect 24822 39888 27000 39944
rect 24761 39886 27000 39888
rect 24761 39883 24827 39886
rect 26200 39856 27000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 19609 39538 19675 39541
rect 20253 39538 20319 39541
rect 19609 39536 20319 39538
rect 19609 39480 19614 39536
rect 19670 39480 20258 39536
rect 20314 39480 20319 39536
rect 19609 39478 20319 39480
rect 19609 39475 19675 39478
rect 20253 39475 20319 39478
rect 23289 39266 23355 39269
rect 23841 39266 23907 39269
rect 23289 39264 23907 39266
rect 23289 39208 23294 39264
rect 23350 39208 23846 39264
rect 23902 39208 23907 39264
rect 23289 39206 23907 39208
rect 23289 39203 23355 39206
rect 23841 39203 23907 39206
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 24853 39130 24919 39133
rect 26200 39130 27000 39160
rect 24853 39128 27000 39130
rect 24853 39072 24858 39128
rect 24914 39072 27000 39128
rect 24853 39070 27000 39072
rect 24853 39067 24919 39070
rect 26200 39040 27000 39070
rect 18413 38858 18479 38861
rect 18638 38858 18644 38860
rect 18413 38856 18644 38858
rect 18413 38800 18418 38856
rect 18474 38800 18644 38856
rect 18413 38798 18644 38800
rect 18413 38795 18479 38798
rect 18638 38796 18644 38798
rect 18708 38796 18714 38860
rect 16021 38724 16087 38725
rect 16021 38722 16068 38724
rect 15976 38720 16068 38722
rect 15976 38664 16026 38720
rect 15976 38662 16068 38664
rect 16021 38660 16068 38662
rect 16132 38660 16138 38724
rect 16021 38659 16087 38660
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 8845 38586 8911 38589
rect 12750 38586 12756 38588
rect 8845 38584 12756 38586
rect 8845 38528 8850 38584
rect 8906 38528 12756 38584
rect 8845 38526 12756 38528
rect 8845 38523 8911 38526
rect 12750 38524 12756 38526
rect 12820 38524 12826 38588
rect 14273 38586 14339 38589
rect 17309 38586 17375 38589
rect 14273 38584 17375 38586
rect 14273 38528 14278 38584
rect 14334 38528 17314 38584
rect 17370 38528 17375 38584
rect 14273 38526 17375 38528
rect 14273 38523 14339 38526
rect 17309 38523 17375 38526
rect 13261 38450 13327 38453
rect 19742 38450 19748 38452
rect 13261 38448 19748 38450
rect 13261 38392 13266 38448
rect 13322 38392 19748 38448
rect 13261 38390 19748 38392
rect 13261 38387 13327 38390
rect 19742 38388 19748 38390
rect 19812 38388 19818 38452
rect 0 38314 800 38344
rect 1301 38314 1367 38317
rect 0 38312 1367 38314
rect 0 38256 1306 38312
rect 1362 38256 1367 38312
rect 0 38254 1367 38256
rect 0 38224 800 38254
rect 1301 38251 1367 38254
rect 8201 38314 8267 38317
rect 11605 38314 11671 38317
rect 13813 38314 13879 38317
rect 8201 38312 13879 38314
rect 8201 38256 8206 38312
rect 8262 38256 11610 38312
rect 11666 38256 13818 38312
rect 13874 38256 13879 38312
rect 8201 38254 13879 38256
rect 8201 38251 8267 38254
rect 11605 38251 11671 38254
rect 13813 38251 13879 38254
rect 25313 38314 25379 38317
rect 26200 38314 27000 38344
rect 25313 38312 27000 38314
rect 25313 38256 25318 38312
rect 25374 38256 27000 38312
rect 25313 38254 27000 38256
rect 25313 38251 25379 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 12750 37980 12756 38044
rect 12820 38042 12826 38044
rect 16113 38042 16179 38045
rect 12820 38040 16179 38042
rect 12820 37984 16118 38040
rect 16174 37984 16179 38040
rect 12820 37982 16179 37984
rect 12820 37980 12826 37982
rect 16113 37979 16179 37982
rect 12525 37906 12591 37909
rect 20253 37906 20319 37909
rect 12525 37904 20319 37906
rect 12525 37848 12530 37904
rect 12586 37848 20258 37904
rect 20314 37848 20319 37904
rect 12525 37846 20319 37848
rect 12525 37843 12591 37846
rect 20253 37843 20319 37846
rect 10225 37770 10291 37773
rect 10501 37770 10567 37773
rect 10225 37768 10567 37770
rect 10225 37712 10230 37768
rect 10286 37712 10506 37768
rect 10562 37712 10567 37768
rect 10225 37710 10567 37712
rect 10225 37707 10291 37710
rect 10501 37707 10567 37710
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 25313 37498 25379 37501
rect 26200 37498 27000 37528
rect 25313 37496 27000 37498
rect 25313 37440 25318 37496
rect 25374 37440 27000 37496
rect 25313 37438 27000 37440
rect 25313 37435 25379 37438
rect 26200 37408 27000 37438
rect 12065 37362 12131 37365
rect 15193 37362 15259 37365
rect 12065 37360 15259 37362
rect 12065 37304 12070 37360
rect 12126 37304 15198 37360
rect 15254 37304 15259 37360
rect 12065 37302 15259 37304
rect 12065 37299 12131 37302
rect 15193 37299 15259 37302
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 15469 36954 15535 36957
rect 16246 36954 16252 36956
rect 15469 36952 16252 36954
rect 15469 36896 15474 36952
rect 15530 36896 16252 36952
rect 15469 36894 16252 36896
rect 15469 36891 15535 36894
rect 16246 36892 16252 36894
rect 16316 36892 16322 36956
rect 9765 36818 9831 36821
rect 9949 36818 10015 36821
rect 16665 36818 16731 36821
rect 9765 36816 16731 36818
rect 9765 36760 9770 36816
rect 9826 36760 9954 36816
rect 10010 36760 16670 36816
rect 16726 36760 16731 36816
rect 9765 36758 16731 36760
rect 9765 36755 9831 36758
rect 9949 36755 10015 36758
rect 16665 36755 16731 36758
rect 15837 36682 15903 36685
rect 22277 36682 22343 36685
rect 22502 36682 22508 36684
rect 15837 36680 22508 36682
rect 15837 36624 15842 36680
rect 15898 36624 22282 36680
rect 22338 36624 22508 36680
rect 15837 36622 22508 36624
rect 15837 36619 15903 36622
rect 22277 36619 22343 36622
rect 22502 36620 22508 36622
rect 22572 36620 22578 36684
rect 25313 36682 25379 36685
rect 26200 36682 27000 36712
rect 25313 36680 27000 36682
rect 25313 36624 25318 36680
rect 25374 36624 27000 36680
rect 25313 36622 27000 36624
rect 25313 36619 25379 36622
rect 26200 36592 27000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 12566 36212 12572 36276
rect 12636 36274 12642 36276
rect 13813 36274 13879 36277
rect 12636 36272 13879 36274
rect 12636 36216 13818 36272
rect 13874 36216 13879 36272
rect 12636 36214 13879 36216
rect 12636 36212 12642 36214
rect 13813 36211 13879 36214
rect 8569 36138 8635 36141
rect 15653 36138 15719 36141
rect 8569 36136 15719 36138
rect 8569 36080 8574 36136
rect 8630 36080 15658 36136
rect 15714 36080 15719 36136
rect 8569 36078 15719 36080
rect 8569 36075 8635 36078
rect 15653 36075 15719 36078
rect 7946 35936 8262 35937
rect 0 35866 800 35896
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 1577 35866 1643 35869
rect 0 35864 1643 35866
rect 0 35808 1582 35864
rect 1638 35808 1643 35864
rect 0 35806 1643 35808
rect 0 35776 800 35806
rect 1577 35803 1643 35806
rect 8661 35866 8727 35869
rect 12433 35866 12499 35869
rect 8661 35864 12499 35866
rect 8661 35808 8666 35864
rect 8722 35808 12438 35864
rect 12494 35808 12499 35864
rect 8661 35806 12499 35808
rect 8661 35803 8727 35806
rect 12433 35803 12499 35806
rect 25313 35866 25379 35869
rect 26200 35866 27000 35896
rect 25313 35864 27000 35866
rect 25313 35808 25318 35864
rect 25374 35808 27000 35864
rect 25313 35806 27000 35808
rect 25313 35803 25379 35806
rect 26200 35776 27000 35806
rect 19885 35458 19951 35461
rect 22553 35458 22619 35461
rect 19885 35456 22619 35458
rect 19885 35400 19890 35456
rect 19946 35400 22558 35456
rect 22614 35400 22619 35456
rect 19885 35398 22619 35400
rect 19885 35395 19951 35398
rect 22553 35395 22619 35398
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 25313 35050 25379 35053
rect 26200 35050 27000 35080
rect 25313 35048 27000 35050
rect 25313 34992 25318 35048
rect 25374 34992 27000 35048
rect 25313 34990 27000 34992
rect 25313 34987 25379 34990
rect 26200 34960 27000 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 25313 34234 25379 34237
rect 26200 34234 27000 34264
rect 25313 34232 27000 34234
rect 25313 34176 25318 34232
rect 25374 34176 27000 34232
rect 25313 34174 27000 34176
rect 25313 34171 25379 34174
rect 26200 34144 27000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 20253 33554 20319 33557
rect 21357 33554 21423 33557
rect 20253 33552 21423 33554
rect 20253 33496 20258 33552
rect 20314 33496 21362 33552
rect 21418 33496 21423 33552
rect 20253 33494 21423 33496
rect 20253 33491 20319 33494
rect 21357 33491 21423 33494
rect 0 33418 800 33448
rect 1209 33418 1275 33421
rect 0 33416 1275 33418
rect 0 33360 1214 33416
rect 1270 33360 1275 33416
rect 0 33358 1275 33360
rect 0 33328 800 33358
rect 1209 33355 1275 33358
rect 25405 33418 25471 33421
rect 26200 33418 27000 33448
rect 25405 33416 27000 33418
rect 25405 33360 25410 33416
rect 25466 33360 27000 33416
rect 25405 33358 27000 33360
rect 25405 33355 25471 33358
rect 26200 33328 27000 33358
rect 12525 33284 12591 33285
rect 12525 33282 12572 33284
rect 12480 33280 12572 33282
rect 12480 33224 12530 33280
rect 12480 33222 12572 33224
rect 12525 33220 12572 33222
rect 12636 33220 12642 33284
rect 12525 33219 12591 33220
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 19190 33084 19196 33148
rect 19260 33146 19266 33148
rect 22369 33146 22435 33149
rect 19260 33144 22435 33146
rect 19260 33088 22374 33144
rect 22430 33088 22435 33144
rect 19260 33086 22435 33088
rect 19260 33084 19266 33086
rect 22369 33083 22435 33086
rect 11605 33012 11671 33013
rect 11605 33010 11652 33012
rect 11560 33008 11652 33010
rect 11560 32952 11610 33008
rect 11560 32950 11652 32952
rect 11605 32948 11652 32950
rect 11716 32948 11722 33012
rect 21357 33010 21423 33013
rect 22461 33012 22527 33013
rect 22461 33010 22508 33012
rect 21222 33008 21423 33010
rect 21222 32952 21362 33008
rect 21418 32952 21423 33008
rect 21222 32950 21423 32952
rect 22416 33008 22508 33010
rect 22416 32952 22466 33008
rect 22416 32950 22508 32952
rect 11605 32947 11671 32948
rect 21222 32741 21282 32950
rect 21357 32947 21423 32950
rect 22461 32948 22508 32950
rect 22572 32948 22578 33012
rect 22461 32947 22527 32948
rect 21222 32736 21331 32741
rect 21909 32738 21975 32741
rect 22369 32738 22435 32741
rect 21222 32680 21270 32736
rect 21326 32680 21331 32736
rect 21222 32678 21331 32680
rect 21265 32675 21331 32678
rect 21774 32736 22435 32738
rect 21774 32680 21914 32736
rect 21970 32680 22374 32736
rect 22430 32680 22435 32736
rect 21774 32678 22435 32680
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 5441 32468 5507 32469
rect 5390 32466 5396 32468
rect 5350 32406 5396 32466
rect 5460 32464 5507 32468
rect 5502 32408 5507 32464
rect 5390 32404 5396 32406
rect 5460 32404 5507 32408
rect 5441 32403 5507 32404
rect 13997 32466 14063 32469
rect 14406 32466 14412 32468
rect 13997 32464 14412 32466
rect 13997 32408 14002 32464
rect 14058 32408 14412 32464
rect 13997 32406 14412 32408
rect 13997 32403 14063 32406
rect 14406 32404 14412 32406
rect 14476 32404 14482 32468
rect 16573 32466 16639 32469
rect 21774 32466 21834 32678
rect 21909 32675 21975 32678
rect 22369 32675 22435 32678
rect 21909 32602 21975 32605
rect 23790 32602 23796 32604
rect 21909 32600 23796 32602
rect 21909 32544 21914 32600
rect 21970 32544 23796 32600
rect 21909 32542 23796 32544
rect 21909 32539 21975 32542
rect 23790 32540 23796 32542
rect 23860 32540 23866 32604
rect 25313 32602 25379 32605
rect 26200 32602 27000 32632
rect 25313 32600 27000 32602
rect 25313 32544 25318 32600
rect 25374 32544 27000 32600
rect 25313 32542 27000 32544
rect 25313 32539 25379 32542
rect 26200 32512 27000 32542
rect 16573 32464 21834 32466
rect 16573 32408 16578 32464
rect 16634 32408 21834 32464
rect 16573 32406 21834 32408
rect 16573 32403 16639 32406
rect 12249 32332 12315 32333
rect 12198 32268 12204 32332
rect 12268 32330 12315 32332
rect 20161 32330 20227 32333
rect 25129 32330 25195 32333
rect 12268 32328 12360 32330
rect 12310 32272 12360 32328
rect 12268 32270 12360 32272
rect 20161 32328 25195 32330
rect 20161 32272 20166 32328
rect 20222 32272 25134 32328
rect 25190 32272 25195 32328
rect 20161 32270 25195 32272
rect 12268 32268 12315 32270
rect 12249 32267 12315 32268
rect 20161 32267 20227 32270
rect 25129 32267 25195 32270
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 19977 32058 20043 32061
rect 20529 32058 20595 32061
rect 19977 32056 20595 32058
rect 19977 32000 19982 32056
rect 20038 32000 20534 32056
rect 20590 32000 20595 32056
rect 19977 31998 20595 32000
rect 19977 31995 20043 31998
rect 20529 31995 20595 31998
rect 9765 31922 9831 31925
rect 17401 31922 17467 31925
rect 9765 31920 17467 31922
rect 9765 31864 9770 31920
rect 9826 31864 17406 31920
rect 17462 31864 17467 31920
rect 9765 31862 17467 31864
rect 9765 31859 9831 31862
rect 17401 31859 17467 31862
rect 19425 31922 19491 31925
rect 19558 31922 19564 31924
rect 19425 31920 19564 31922
rect 19425 31864 19430 31920
rect 19486 31864 19564 31920
rect 19425 31862 19564 31864
rect 19425 31859 19491 31862
rect 19558 31860 19564 31862
rect 19628 31860 19634 31924
rect 18229 31786 18295 31789
rect 21766 31786 21772 31788
rect 18229 31784 21772 31786
rect 18229 31728 18234 31784
rect 18290 31728 21772 31784
rect 18229 31726 21772 31728
rect 18229 31723 18295 31726
rect 21766 31724 21772 31726
rect 21836 31724 21842 31788
rect 25313 31786 25379 31789
rect 26200 31786 27000 31816
rect 25313 31784 27000 31786
rect 25313 31728 25318 31784
rect 25374 31728 27000 31784
rect 25313 31726 27000 31728
rect 25313 31723 25379 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 19977 31242 20043 31245
rect 20110 31242 20116 31244
rect 19977 31240 20116 31242
rect 19977 31184 19982 31240
rect 20038 31184 20116 31240
rect 19977 31182 20116 31184
rect 19977 31179 20043 31182
rect 20110 31180 20116 31182
rect 20180 31180 20186 31244
rect 2946 31040 3262 31041
rect 0 30970 800 31000
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 1301 30970 1367 30973
rect 0 30968 1367 30970
rect 0 30912 1306 30968
rect 1362 30912 1367 30968
rect 0 30910 1367 30912
rect 0 30880 800 30910
rect 1301 30907 1367 30910
rect 25313 30970 25379 30973
rect 26200 30970 27000 31000
rect 25313 30968 27000 30970
rect 25313 30912 25318 30968
rect 25374 30912 27000 30968
rect 25313 30910 27000 30912
rect 25313 30907 25379 30910
rect 26200 30880 27000 30910
rect 19742 30772 19748 30836
rect 19812 30834 19818 30836
rect 19885 30834 19951 30837
rect 19812 30832 19951 30834
rect 19812 30776 19890 30832
rect 19946 30776 19951 30832
rect 19812 30774 19951 30776
rect 19812 30772 19818 30774
rect 19885 30771 19951 30774
rect 10174 30636 10180 30700
rect 10244 30698 10250 30700
rect 11421 30698 11487 30701
rect 10244 30696 11487 30698
rect 10244 30640 11426 30696
rect 11482 30640 11487 30696
rect 10244 30638 11487 30640
rect 10244 30636 10250 30638
rect 11421 30635 11487 30638
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 18045 30290 18111 30293
rect 18689 30290 18755 30293
rect 21950 30290 21956 30292
rect 18045 30288 21956 30290
rect 18045 30232 18050 30288
rect 18106 30232 18694 30288
rect 18750 30232 21956 30288
rect 18045 30230 21956 30232
rect 18045 30227 18111 30230
rect 18689 30227 18755 30230
rect 21950 30228 21956 30230
rect 22020 30228 22026 30292
rect 25313 30154 25379 30157
rect 26200 30154 27000 30184
rect 25313 30152 27000 30154
rect 25313 30096 25318 30152
rect 25374 30096 27000 30152
rect 25313 30094 27000 30096
rect 25313 30091 25379 30094
rect 26200 30064 27000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 25497 29338 25563 29341
rect 26200 29338 27000 29368
rect 25497 29336 27000 29338
rect 25497 29280 25502 29336
rect 25558 29280 27000 29336
rect 25497 29278 27000 29280
rect 25497 29275 25563 29278
rect 26200 29248 27000 29278
rect 16113 29202 16179 29205
rect 16246 29202 16252 29204
rect 16113 29200 16252 29202
rect 16113 29144 16118 29200
rect 16174 29144 16252 29200
rect 16113 29142 16252 29144
rect 16113 29139 16179 29142
rect 16246 29140 16252 29142
rect 16316 29202 16322 29204
rect 21541 29202 21607 29205
rect 16316 29200 21607 29202
rect 16316 29144 21546 29200
rect 21602 29144 21607 29200
rect 16316 29142 21607 29144
rect 16316 29140 16322 29142
rect 21541 29139 21607 29142
rect 16389 29068 16455 29069
rect 15694 29004 15700 29068
rect 15764 29066 15770 29068
rect 16389 29066 16436 29068
rect 15764 29064 16436 29066
rect 16500 29066 16506 29068
rect 20161 29066 20227 29069
rect 20478 29066 20484 29068
rect 15764 29008 16394 29064
rect 15764 29006 16436 29008
rect 15764 29004 15770 29006
rect 16389 29004 16436 29006
rect 16500 29006 16582 29066
rect 20161 29064 20484 29066
rect 20161 29008 20166 29064
rect 20222 29008 20484 29064
rect 20161 29006 20484 29008
rect 16500 29004 16506 29006
rect 16389 29003 16455 29004
rect 20161 29003 20227 29006
rect 20478 29004 20484 29006
rect 20548 29004 20554 29068
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 0 28522 800 28552
rect 1301 28522 1367 28525
rect 0 28520 1367 28522
rect 0 28464 1306 28520
rect 1362 28464 1367 28520
rect 0 28462 1367 28464
rect 0 28432 800 28462
rect 1301 28459 1367 28462
rect 18321 28522 18387 28525
rect 21582 28522 21588 28524
rect 18321 28520 21588 28522
rect 18321 28464 18326 28520
rect 18382 28464 21588 28520
rect 18321 28462 21588 28464
rect 18321 28459 18387 28462
rect 21582 28460 21588 28462
rect 21652 28460 21658 28524
rect 24853 28522 24919 28525
rect 26200 28522 27000 28552
rect 24853 28520 27000 28522
rect 24853 28464 24858 28520
rect 24914 28464 27000 28520
rect 24853 28462 27000 28464
rect 24853 28459 24919 28462
rect 26200 28432 27000 28462
rect 14733 28386 14799 28389
rect 16757 28388 16823 28389
rect 16757 28386 16804 28388
rect 14733 28384 16804 28386
rect 14733 28328 14738 28384
rect 14794 28328 16762 28384
rect 14733 28326 16804 28328
rect 14733 28323 14799 28326
rect 16757 28324 16804 28326
rect 16868 28324 16874 28388
rect 20069 28386 20135 28389
rect 22686 28386 22692 28388
rect 20069 28384 22692 28386
rect 20069 28328 20074 28384
rect 20130 28328 22692 28384
rect 20069 28326 22692 28328
rect 16757 28323 16823 28324
rect 20069 28323 20135 28326
rect 22686 28324 22692 28326
rect 22756 28324 22762 28388
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 14958 28188 14964 28252
rect 15028 28250 15034 28252
rect 15285 28250 15351 28253
rect 15929 28252 15995 28253
rect 15028 28248 15351 28250
rect 15028 28192 15290 28248
rect 15346 28192 15351 28248
rect 15028 28190 15351 28192
rect 15028 28188 15034 28190
rect 15285 28187 15351 28190
rect 15878 28188 15884 28252
rect 15948 28250 15995 28252
rect 15948 28248 16040 28250
rect 15990 28192 16040 28248
rect 15948 28190 16040 28192
rect 15948 28188 15995 28190
rect 15929 28187 15995 28188
rect 16021 27978 16087 27981
rect 16246 27978 16252 27980
rect 16021 27976 16252 27978
rect 16021 27920 16026 27976
rect 16082 27920 16252 27976
rect 16021 27918 16252 27920
rect 16021 27915 16087 27918
rect 16246 27916 16252 27918
rect 16316 27916 16322 27980
rect 19742 27780 19748 27844
rect 19812 27842 19818 27844
rect 20069 27842 20135 27845
rect 19812 27840 20135 27842
rect 19812 27784 20074 27840
rect 20130 27784 20135 27840
rect 19812 27782 20135 27784
rect 19812 27780 19818 27782
rect 20069 27779 20135 27782
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 24117 27706 24183 27709
rect 26200 27706 27000 27736
rect 24117 27704 27000 27706
rect 24117 27648 24122 27704
rect 24178 27648 27000 27704
rect 24117 27646 27000 27648
rect 24117 27643 24183 27646
rect 26200 27616 27000 27646
rect 17125 27436 17191 27437
rect 17125 27432 17172 27436
rect 17236 27434 17242 27436
rect 17125 27376 17130 27432
rect 17125 27372 17172 27376
rect 17236 27374 17282 27434
rect 17236 27372 17242 27374
rect 17125 27371 17191 27372
rect 15142 27236 15148 27300
rect 15212 27298 15218 27300
rect 15377 27298 15443 27301
rect 15212 27296 15443 27298
rect 15212 27240 15382 27296
rect 15438 27240 15443 27296
rect 15212 27238 15443 27240
rect 15212 27236 15218 27238
rect 15377 27235 15443 27238
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 25497 26890 25563 26893
rect 26200 26890 27000 26920
rect 25497 26888 27000 26890
rect 25497 26832 25502 26888
rect 25558 26832 27000 26888
rect 25497 26830 27000 26832
rect 25497 26827 25563 26830
rect 26200 26800 27000 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 7946 26144 8262 26145
rect 0 26074 800 26104
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 2773 26074 2839 26077
rect 0 26072 2839 26074
rect 0 26016 2778 26072
rect 2834 26016 2839 26072
rect 0 26014 2839 26016
rect 0 25984 800 26014
rect 2773 26011 2839 26014
rect 25313 26074 25379 26077
rect 26200 26074 27000 26104
rect 25313 26072 27000 26074
rect 25313 26016 25318 26072
rect 25374 26016 27000 26072
rect 25313 26014 27000 26016
rect 25313 26011 25379 26014
rect 26200 25984 27000 26014
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 16798 25196 16804 25260
rect 16868 25258 16874 25260
rect 23749 25258 23815 25261
rect 16868 25256 23815 25258
rect 16868 25200 23754 25256
rect 23810 25200 23815 25256
rect 16868 25198 23815 25200
rect 16868 25196 16874 25198
rect 23749 25195 23815 25198
rect 25129 25258 25195 25261
rect 26200 25258 27000 25288
rect 25129 25256 27000 25258
rect 25129 25200 25134 25256
rect 25190 25200 27000 25256
rect 25129 25198 27000 25200
rect 25129 25195 25195 25198
rect 26200 25168 27000 25198
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 24853 24442 24919 24445
rect 26200 24442 27000 24472
rect 24853 24440 27000 24442
rect 24853 24384 24858 24440
rect 24914 24384 27000 24440
rect 24853 24382 27000 24384
rect 24853 24379 24919 24382
rect 26200 24352 27000 24382
rect 11053 24034 11119 24037
rect 11881 24034 11947 24037
rect 12014 24034 12020 24036
rect 11053 24032 12020 24034
rect 11053 23976 11058 24032
rect 11114 23976 11886 24032
rect 11942 23976 12020 24032
rect 11053 23974 12020 23976
rect 11053 23971 11119 23974
rect 11881 23971 11947 23974
rect 12014 23972 12020 23974
rect 12084 23972 12090 24036
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 0 23626 800 23656
rect 1301 23626 1367 23629
rect 0 23624 1367 23626
rect 0 23568 1306 23624
rect 1362 23568 1367 23624
rect 0 23566 1367 23568
rect 0 23536 800 23566
rect 1301 23563 1367 23566
rect 23841 23626 23907 23629
rect 26200 23626 27000 23656
rect 23841 23624 27000 23626
rect 23841 23568 23846 23624
rect 23902 23568 27000 23624
rect 23841 23566 27000 23568
rect 23841 23563 23907 23566
rect 26200 23536 27000 23566
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 24669 22810 24735 22813
rect 26200 22810 27000 22840
rect 24669 22808 27000 22810
rect 24669 22752 24674 22808
rect 24730 22752 27000 22808
rect 24669 22750 27000 22752
rect 24669 22747 24735 22750
rect 26200 22720 27000 22750
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 13537 21994 13603 21997
rect 16062 21994 16068 21996
rect 13537 21992 16068 21994
rect 13537 21936 13542 21992
rect 13598 21936 16068 21992
rect 13537 21934 16068 21936
rect 13537 21931 13603 21934
rect 16062 21932 16068 21934
rect 16132 21932 16138 21996
rect 24853 21994 24919 21997
rect 26200 21994 27000 22024
rect 24853 21992 27000 21994
rect 24853 21936 24858 21992
rect 24914 21936 27000 21992
rect 24853 21934 27000 21936
rect 24853 21931 24919 21934
rect 26200 21904 27000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 14406 21660 14412 21724
rect 14476 21722 14482 21724
rect 14641 21722 14707 21725
rect 14476 21720 14707 21722
rect 14476 21664 14646 21720
rect 14702 21664 14707 21720
rect 14476 21662 14707 21664
rect 14476 21660 14482 21662
rect 14641 21659 14707 21662
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 1301 21178 1367 21181
rect 0 21176 1367 21178
rect 0 21120 1306 21176
rect 1362 21120 1367 21176
rect 0 21118 1367 21120
rect 0 21088 800 21118
rect 1301 21115 1367 21118
rect 23381 21178 23447 21181
rect 26200 21178 27000 21208
rect 23381 21176 27000 21178
rect 23381 21120 23386 21176
rect 23442 21120 27000 21176
rect 23381 21118 27000 21120
rect 23381 21115 23447 21118
rect 26200 21088 27000 21118
rect 16113 20772 16179 20773
rect 16062 20770 16068 20772
rect 16022 20710 16068 20770
rect 16132 20768 16179 20772
rect 16174 20712 16179 20768
rect 16062 20708 16068 20710
rect 16132 20708 16179 20712
rect 16113 20707 16179 20708
rect 19149 20770 19215 20773
rect 19742 20770 19748 20772
rect 19149 20768 19748 20770
rect 19149 20712 19154 20768
rect 19210 20712 19748 20768
rect 19149 20710 19748 20712
rect 19149 20707 19215 20710
rect 19742 20708 19748 20710
rect 19812 20770 19818 20772
rect 19977 20770 20043 20773
rect 19812 20768 20043 20770
rect 19812 20712 19982 20768
rect 20038 20712 20043 20768
rect 19812 20710 20043 20712
rect 19812 20708 19818 20710
rect 19977 20707 20043 20710
rect 20253 20770 20319 20773
rect 20478 20770 20484 20772
rect 20253 20768 20484 20770
rect 20253 20712 20258 20768
rect 20314 20712 20484 20768
rect 20253 20710 20484 20712
rect 20253 20707 20319 20710
rect 20478 20708 20484 20710
rect 20548 20708 20554 20772
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 17309 20636 17375 20637
rect 17309 20634 17356 20636
rect 17264 20632 17356 20634
rect 17264 20576 17314 20632
rect 17264 20574 17356 20576
rect 17309 20572 17356 20574
rect 17420 20572 17426 20636
rect 18505 20634 18571 20637
rect 19558 20634 19564 20636
rect 18505 20632 19564 20634
rect 18505 20576 18510 20632
rect 18566 20576 19564 20632
rect 18505 20574 19564 20576
rect 17309 20571 17375 20572
rect 18505 20571 18571 20574
rect 19558 20572 19564 20574
rect 19628 20572 19634 20636
rect 24945 20362 25011 20365
rect 26200 20362 27000 20392
rect 24945 20360 27000 20362
rect 24945 20304 24950 20360
rect 25006 20304 27000 20360
rect 24945 20302 27000 20304
rect 24945 20299 25011 20302
rect 26200 20272 27000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 17769 19954 17835 19957
rect 18638 19954 18644 19956
rect 17769 19952 18644 19954
rect 17769 19896 17774 19952
rect 17830 19896 18644 19952
rect 17769 19894 18644 19896
rect 17769 19891 17835 19894
rect 18638 19892 18644 19894
rect 18708 19892 18714 19956
rect 8661 19684 8727 19685
rect 14733 19684 14799 19685
rect 8661 19682 8708 19684
rect 8616 19680 8708 19682
rect 8616 19624 8666 19680
rect 8616 19622 8708 19624
rect 8661 19620 8708 19622
rect 8772 19620 8778 19684
rect 14733 19682 14780 19684
rect 14688 19680 14780 19682
rect 14688 19624 14738 19680
rect 14688 19622 14780 19624
rect 14733 19620 14780 19622
rect 14844 19620 14850 19684
rect 8661 19619 8727 19620
rect 14733 19619 14799 19620
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 23289 19546 23355 19549
rect 26200 19546 27000 19576
rect 23289 19544 27000 19546
rect 23289 19488 23294 19544
rect 23350 19488 27000 19544
rect 23289 19486 27000 19488
rect 23289 19483 23355 19486
rect 26200 19456 27000 19486
rect 12157 19412 12223 19413
rect 18413 19412 18479 19413
rect 12157 19408 12204 19412
rect 12268 19410 12274 19412
rect 12157 19352 12162 19408
rect 12157 19348 12204 19352
rect 12268 19350 12314 19410
rect 18413 19408 18460 19412
rect 18524 19410 18530 19412
rect 18413 19352 18418 19408
rect 12268 19348 12274 19350
rect 18413 19348 18460 19352
rect 18524 19350 18570 19410
rect 18524 19348 18530 19350
rect 12157 19347 12223 19348
rect 18413 19347 18479 19348
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 0 18730 800 18760
rect 1301 18730 1367 18733
rect 0 18728 1367 18730
rect 0 18672 1306 18728
rect 1362 18672 1367 18728
rect 0 18670 1367 18672
rect 0 18640 800 18670
rect 1301 18667 1367 18670
rect 18321 18730 18387 18733
rect 20110 18730 20116 18732
rect 18321 18728 20116 18730
rect 18321 18672 18326 18728
rect 18382 18672 20116 18728
rect 18321 18670 20116 18672
rect 18321 18667 18387 18670
rect 20110 18668 20116 18670
rect 20180 18668 20186 18732
rect 23381 18730 23447 18733
rect 26200 18730 27000 18760
rect 23381 18728 27000 18730
rect 23381 18672 23386 18728
rect 23442 18672 27000 18728
rect 23381 18670 27000 18672
rect 23381 18667 23447 18670
rect 26200 18640 27000 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 12893 18322 12959 18325
rect 15142 18322 15148 18324
rect 12893 18320 15148 18322
rect 12893 18264 12898 18320
rect 12954 18264 15148 18320
rect 12893 18262 15148 18264
rect 12893 18259 12959 18262
rect 15142 18260 15148 18262
rect 15212 18322 15218 18324
rect 16665 18322 16731 18325
rect 15212 18320 16731 18322
rect 15212 18264 16670 18320
rect 16726 18264 16731 18320
rect 15212 18262 16731 18264
rect 15212 18260 15218 18262
rect 16665 18259 16731 18262
rect 4981 18186 5047 18189
rect 5390 18186 5396 18188
rect 4981 18184 5396 18186
rect 4981 18128 4986 18184
rect 5042 18128 5396 18184
rect 4981 18126 5396 18128
rect 4981 18123 5047 18126
rect 5390 18124 5396 18126
rect 5460 18124 5466 18188
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 12525 17916 12591 17917
rect 12525 17914 12572 17916
rect 12480 17912 12572 17914
rect 12480 17856 12530 17912
rect 12480 17854 12572 17856
rect 12525 17852 12572 17854
rect 12636 17852 12642 17916
rect 24853 17914 24919 17917
rect 26200 17914 27000 17944
rect 24853 17912 27000 17914
rect 24853 17856 24858 17912
rect 24914 17856 27000 17912
rect 24853 17854 27000 17856
rect 12525 17851 12591 17852
rect 24853 17851 24919 17854
rect 26200 17824 27000 17854
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 24761 17098 24827 17101
rect 26200 17098 27000 17128
rect 24761 17096 27000 17098
rect 24761 17040 24766 17096
rect 24822 17040 27000 17096
rect 24761 17038 27000 17040
rect 24761 17035 24827 17038
rect 26200 17008 27000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 16297 16828 16363 16829
rect 16246 16826 16252 16828
rect 16206 16766 16252 16826
rect 16316 16824 16363 16828
rect 16358 16768 16363 16824
rect 16246 16764 16252 16766
rect 16316 16764 16363 16768
rect 16297 16763 16363 16764
rect 2497 16554 2563 16557
rect 4061 16554 4127 16557
rect 9489 16554 9555 16557
rect 2497 16552 9555 16554
rect 2497 16496 2502 16552
rect 2558 16496 4066 16552
rect 4122 16496 9494 16552
rect 9550 16496 9555 16552
rect 2497 16494 9555 16496
rect 2497 16491 2563 16494
rect 4061 16491 4127 16494
rect 9489 16491 9555 16494
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 14733 16282 14799 16285
rect 14958 16282 14964 16284
rect 14733 16280 14964 16282
rect 14733 16224 14738 16280
rect 14794 16224 14964 16280
rect 14733 16222 14964 16224
rect 14733 16219 14799 16222
rect 14958 16220 14964 16222
rect 15028 16220 15034 16284
rect 15694 16220 15700 16284
rect 15764 16282 15770 16284
rect 15929 16282 15995 16285
rect 15764 16280 15995 16282
rect 15764 16224 15934 16280
rect 15990 16224 15995 16280
rect 15764 16222 15995 16224
rect 15764 16220 15770 16222
rect 15929 16219 15995 16222
rect 24669 16282 24735 16285
rect 26200 16282 27000 16312
rect 24669 16280 27000 16282
rect 24669 16224 24674 16280
rect 24730 16224 27000 16280
rect 24669 16222 27000 16224
rect 24669 16219 24735 16222
rect 26200 16192 27000 16222
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 24945 15466 25011 15469
rect 26200 15466 27000 15496
rect 24945 15464 27000 15466
rect 24945 15408 24950 15464
rect 25006 15408 27000 15464
rect 24945 15406 27000 15408
rect 24945 15403 25011 15406
rect 26200 15376 27000 15406
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 24761 14650 24827 14653
rect 26200 14650 27000 14680
rect 24761 14648 27000 14650
rect 24761 14592 24766 14648
rect 24822 14592 27000 14648
rect 24761 14590 27000 14592
rect 24761 14587 24827 14590
rect 26200 14560 27000 14590
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 12014 14044 12020 14108
rect 12084 14106 12090 14108
rect 13537 14106 13603 14109
rect 12084 14104 13603 14106
rect 12084 14048 13542 14104
rect 13598 14048 13603 14104
rect 12084 14046 13603 14048
rect 12084 14044 12090 14046
rect 13537 14043 13603 14046
rect 0 13834 800 13864
rect 1301 13834 1367 13837
rect 0 13832 1367 13834
rect 0 13776 1306 13832
rect 1362 13776 1367 13832
rect 0 13774 1367 13776
rect 0 13744 800 13774
rect 1301 13771 1367 13774
rect 23289 13834 23355 13837
rect 26200 13834 27000 13864
rect 23289 13832 27000 13834
rect 23289 13776 23294 13832
rect 23350 13776 27000 13832
rect 23289 13774 27000 13776
rect 23289 13771 23355 13774
rect 26200 13744 27000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 25497 13018 25563 13021
rect 26200 13018 27000 13048
rect 25497 13016 27000 13018
rect 25497 12960 25502 13016
rect 25558 12960 27000 13016
rect 25497 12958 27000 12960
rect 25497 12955 25563 12958
rect 26200 12928 27000 12958
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 24761 12202 24827 12205
rect 26200 12202 27000 12232
rect 24761 12200 27000 12202
rect 24761 12144 24766 12200
rect 24822 12144 27000 12200
rect 24761 12142 27000 12144
rect 24761 12139 24827 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 3877 11658 3943 11661
rect 1902 11656 3943 11658
rect 1902 11600 3882 11656
rect 3938 11600 3943 11656
rect 1902 11598 3943 11600
rect 0 11386 800 11416
rect 1902 11386 1962 11598
rect 3877 11595 3943 11598
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 0 11326 1962 11386
rect 23381 11386 23447 11389
rect 26200 11386 27000 11416
rect 23381 11384 27000 11386
rect 23381 11328 23386 11384
rect 23442 11328 27000 11384
rect 23381 11326 27000 11328
rect 0 11296 800 11326
rect 23381 11323 23447 11326
rect 26200 11296 27000 11326
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 24669 10570 24735 10573
rect 26200 10570 27000 10600
rect 24669 10568 27000 10570
rect 24669 10512 24674 10568
rect 24730 10512 27000 10568
rect 24669 10510 27000 10512
rect 24669 10507 24735 10510
rect 26200 10480 27000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 24945 9754 25011 9757
rect 26200 9754 27000 9784
rect 24945 9752 27000 9754
rect 24945 9696 24950 9752
rect 25006 9696 27000 9752
rect 24945 9694 27000 9696
rect 24945 9691 25011 9694
rect 26200 9664 27000 9694
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 0 8938 800 8968
rect 3601 8938 3667 8941
rect 0 8936 3667 8938
rect 0 8880 3606 8936
rect 3662 8880 3667 8936
rect 0 8878 3667 8880
rect 0 8848 800 8878
rect 3601 8875 3667 8878
rect 25129 8938 25195 8941
rect 26200 8938 27000 8968
rect 25129 8936 27000 8938
rect 25129 8880 25134 8936
rect 25190 8880 27000 8936
rect 25129 8878 27000 8880
rect 25129 8875 25195 8878
rect 26200 8848 27000 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 24761 8122 24827 8125
rect 26200 8122 27000 8152
rect 24761 8120 27000 8122
rect 24761 8064 24766 8120
rect 24822 8064 27000 8120
rect 24761 8062 27000 8064
rect 24761 8059 24827 8062
rect 26200 8032 27000 8062
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 24669 7306 24735 7309
rect 26200 7306 27000 7336
rect 24669 7304 27000 7306
rect 24669 7248 24674 7304
rect 24730 7248 27000 7304
rect 24669 7246 27000 7248
rect 24669 7243 24735 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 4061 6490 4127 6493
rect 0 6488 4127 6490
rect 0 6432 4066 6488
rect 4122 6432 4127 6488
rect 0 6430 4127 6432
rect 0 6400 800 6430
rect 4061 6427 4127 6430
rect 25037 6490 25103 6493
rect 26200 6490 27000 6520
rect 25037 6488 27000 6490
rect 25037 6432 25042 6488
rect 25098 6432 27000 6488
rect 25037 6430 27000 6432
rect 25037 6427 25103 6430
rect 26200 6400 27000 6430
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 3785 5810 3851 5813
rect 8702 5810 8708 5812
rect 3785 5808 8708 5810
rect 3785 5752 3790 5808
rect 3846 5752 8708 5808
rect 3785 5750 8708 5752
rect 3785 5747 3851 5750
rect 8702 5748 8708 5750
rect 8772 5748 8778 5812
rect 8477 5674 8543 5677
rect 10174 5674 10180 5676
rect 8477 5672 10180 5674
rect 8477 5616 8482 5672
rect 8538 5616 10180 5672
rect 8477 5614 10180 5616
rect 8477 5611 8543 5614
rect 10174 5612 10180 5614
rect 10244 5612 10250 5676
rect 24761 5674 24827 5677
rect 26200 5674 27000 5704
rect 24761 5672 27000 5674
rect 24761 5616 24766 5672
rect 24822 5616 27000 5672
rect 24761 5614 27000 5616
rect 24761 5611 24827 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 9581 5130 9647 5133
rect 14774 5130 14780 5132
rect 9581 5128 14780 5130
rect 9581 5072 9586 5128
rect 9642 5072 14780 5128
rect 9581 5070 14780 5072
rect 9581 5067 9647 5070
rect 14774 5068 14780 5070
rect 14844 5068 14850 5132
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 24485 4858 24551 4861
rect 26200 4858 27000 4888
rect 24485 4856 27000 4858
rect 24485 4800 24490 4856
rect 24546 4800 27000 4856
rect 24485 4798 27000 4800
rect 24485 4795 24551 4798
rect 26200 4768 27000 4798
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 0 4042 800 4072
rect 3693 4042 3759 4045
rect 0 4040 3759 4042
rect 0 3984 3698 4040
rect 3754 3984 3759 4040
rect 0 3982 3759 3984
rect 0 3952 800 3982
rect 3693 3979 3759 3982
rect 18454 3980 18460 4044
rect 18524 4042 18530 4044
rect 18689 4042 18755 4045
rect 18524 4040 18755 4042
rect 18524 3984 18694 4040
rect 18750 3984 18755 4040
rect 18524 3982 18755 3984
rect 18524 3980 18530 3982
rect 18689 3979 18755 3982
rect 22093 4042 22159 4045
rect 26200 4042 27000 4072
rect 22093 4040 27000 4042
rect 22093 3984 22098 4040
rect 22154 3984 27000 4040
rect 22093 3982 27000 3984
rect 22093 3979 22159 3982
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 23289 3226 23355 3229
rect 26200 3226 27000 3256
rect 23289 3224 27000 3226
rect 23289 3168 23294 3224
rect 23350 3168 27000 3224
rect 23289 3166 27000 3168
rect 23289 3163 23355 3166
rect 26200 3136 27000 3166
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 21357 2410 21423 2413
rect 26200 2410 27000 2440
rect 21357 2408 27000 2410
rect 21357 2352 21362 2408
rect 21418 2352 27000 2408
rect 21357 2350 27000 2352
rect 21357 2347 21423 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1594 800 1624
rect 3417 1594 3483 1597
rect 0 1592 3483 1594
rect 0 1536 3422 1592
rect 3478 1536 3483 1592
rect 0 1534 3483 1536
rect 0 1504 800 1534
rect 3417 1531 3483 1534
rect 24853 1594 24919 1597
rect 26200 1594 27000 1624
rect 24853 1592 27000 1594
rect 24853 1536 24858 1592
rect 24914 1536 27000 1592
rect 24853 1534 27000 1536
rect 24853 1531 24919 1534
rect 26200 1504 27000 1534
rect 24945 778 25011 781
rect 26200 778 27000 808
rect 24945 776 27000 778
rect 24945 720 24950 776
rect 25006 720 27000 776
rect 24945 718 27000 720
rect 24945 715 25011 718
rect 26200 688 27000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 16436 52592 16500 52596
rect 16436 52536 16450 52592
rect 16450 52536 16500 52592
rect 16436 52532 16500 52536
rect 17172 52592 17236 52596
rect 17172 52536 17186 52592
rect 17186 52536 17236 52592
rect 17172 52532 17236 52536
rect 23796 52532 23860 52596
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 18644 47636 18708 47700
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 21772 46956 21836 47020
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 22692 46548 22756 46612
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 20116 45928 20180 45932
rect 20116 45872 20130 45928
rect 20130 45872 20180 45928
rect 20116 45868 20180 45872
rect 21956 45928 22020 45932
rect 21956 45872 21970 45928
rect 21970 45872 22020 45928
rect 21956 45868 22020 45872
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 11652 44296 11716 44300
rect 11652 44240 11666 44296
rect 11666 44240 11716 44296
rect 11652 44236 11716 44240
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 19748 43148 19812 43212
rect 16068 43012 16132 43076
rect 21588 43072 21652 43076
rect 21588 43016 21638 43072
rect 21638 43016 21652 43072
rect 21588 43012 21652 43016
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 10916 42468 10980 42532
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 15884 40020 15948 40084
rect 19196 40020 19260 40084
rect 12204 39884 12268 39948
rect 17356 39884 17420 39948
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 18644 38796 18708 38860
rect 16068 38720 16132 38724
rect 16068 38664 16082 38720
rect 16082 38664 16132 38720
rect 16068 38660 16132 38664
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 12756 38524 12820 38588
rect 19748 38388 19812 38452
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 12756 37980 12820 38044
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 16252 36892 16316 36956
rect 22508 36620 22572 36684
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 12572 36212 12636 36276
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 12572 33280 12636 33284
rect 12572 33224 12586 33280
rect 12586 33224 12636 33280
rect 12572 33220 12636 33224
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 19196 33084 19260 33148
rect 11652 33008 11716 33012
rect 11652 32952 11666 33008
rect 11666 32952 11716 33008
rect 11652 32948 11716 32952
rect 22508 33008 22572 33012
rect 22508 32952 22522 33008
rect 22522 32952 22572 33008
rect 22508 32948 22572 32952
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 5396 32464 5460 32468
rect 5396 32408 5446 32464
rect 5446 32408 5460 32464
rect 5396 32404 5460 32408
rect 14412 32404 14476 32468
rect 23796 32540 23860 32604
rect 12204 32328 12268 32332
rect 12204 32272 12254 32328
rect 12254 32272 12268 32328
rect 12204 32268 12268 32272
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 19564 31860 19628 31924
rect 21772 31724 21836 31788
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 20116 31180 20180 31244
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 19748 30772 19812 30836
rect 10180 30636 10244 30700
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 21956 30228 22020 30292
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 16252 29140 16316 29204
rect 15700 29004 15764 29068
rect 16436 29064 16500 29068
rect 16436 29008 16450 29064
rect 16450 29008 16500 29064
rect 16436 29004 16500 29008
rect 20484 29004 20548 29068
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 21588 28460 21652 28524
rect 16804 28384 16868 28388
rect 16804 28328 16818 28384
rect 16818 28328 16868 28384
rect 16804 28324 16868 28328
rect 22692 28324 22756 28388
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 14964 28188 15028 28252
rect 15884 28248 15948 28252
rect 15884 28192 15934 28248
rect 15934 28192 15948 28248
rect 15884 28188 15948 28192
rect 16252 27916 16316 27980
rect 19748 27780 19812 27844
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 17172 27432 17236 27436
rect 17172 27376 17186 27432
rect 17186 27376 17236 27432
rect 17172 27372 17236 27376
rect 15148 27236 15212 27300
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 16804 25196 16868 25260
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 12020 23972 12084 24036
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 16068 21932 16132 21996
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 14412 21660 14476 21724
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 16068 20768 16132 20772
rect 16068 20712 16118 20768
rect 16118 20712 16132 20768
rect 16068 20708 16132 20712
rect 19748 20708 19812 20772
rect 20484 20708 20548 20772
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 17356 20632 17420 20636
rect 17356 20576 17370 20632
rect 17370 20576 17420 20632
rect 17356 20572 17420 20576
rect 19564 20572 19628 20636
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 18644 19892 18708 19956
rect 8708 19680 8772 19684
rect 8708 19624 8722 19680
rect 8722 19624 8772 19680
rect 8708 19620 8772 19624
rect 14780 19680 14844 19684
rect 14780 19624 14794 19680
rect 14794 19624 14844 19680
rect 14780 19620 14844 19624
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 12204 19408 12268 19412
rect 12204 19352 12218 19408
rect 12218 19352 12268 19408
rect 12204 19348 12268 19352
rect 18460 19408 18524 19412
rect 18460 19352 18474 19408
rect 18474 19352 18524 19408
rect 18460 19348 18524 19352
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 20116 18668 20180 18732
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 15148 18260 15212 18324
rect 5396 18124 5460 18188
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 12572 17912 12636 17916
rect 12572 17856 12586 17912
rect 12586 17856 12636 17912
rect 12572 17852 12636 17856
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 16252 16824 16316 16828
rect 16252 16768 16302 16824
rect 16302 16768 16316 16824
rect 16252 16764 16316 16768
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 14964 16220 15028 16284
rect 15700 16220 15764 16284
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 12020 14044 12084 14108
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 8708 5748 8772 5812
rect 10180 5612 10244 5676
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 14780 5068 14844 5132
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18460 3980 18524 4044
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 16435 52596 16501 52597
rect 16435 52532 16436 52596
rect 16500 52532 16501 52596
rect 16435 52531 16501 52532
rect 17171 52596 17237 52597
rect 17171 52532 17172 52596
rect 17236 52532 17237 52596
rect 17171 52531 17237 52532
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 11651 44300 11717 44301
rect 11651 44236 11652 44300
rect 11716 44236 11717 44300
rect 11651 44235 11717 44236
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 10915 42532 10981 42533
rect 10915 42468 10916 42532
rect 10980 42468 10981 42532
rect 10915 42467 10981 42468
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 5395 32468 5461 32469
rect 5395 32404 5396 32468
rect 5460 32404 5461 32468
rect 5395 32403 5461 32404
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 5398 18189 5458 32403
rect 7944 31584 8264 32608
rect 10918 31770 10978 42467
rect 11654 33013 11714 44235
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 16067 43076 16133 43077
rect 16067 43012 16068 43076
rect 16132 43012 16133 43076
rect 16067 43011 16133 43012
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12203 39948 12269 39949
rect 12203 39884 12204 39948
rect 12268 39884 12269 39948
rect 12203 39883 12269 39884
rect 12206 38450 12266 39883
rect 12944 39744 13264 40768
rect 15883 40084 15949 40085
rect 15883 40020 15884 40084
rect 15948 40020 15949 40084
rect 15883 40019 15949 40020
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12755 38588 12821 38589
rect 12755 38524 12756 38588
rect 12820 38524 12821 38588
rect 12755 38523 12821 38524
rect 12206 38390 12634 38450
rect 12574 36277 12634 38390
rect 12758 38045 12818 38523
rect 12755 38044 12821 38045
rect 12755 37980 12756 38044
rect 12820 37980 12821 38044
rect 12755 37979 12821 37980
rect 12571 36276 12637 36277
rect 12571 36212 12572 36276
rect 12636 36212 12637 36276
rect 12571 36211 12637 36212
rect 12574 35910 12634 36211
rect 12206 35850 12634 35910
rect 11651 33012 11717 33013
rect 11651 32948 11652 33012
rect 11716 32948 11717 33012
rect 11651 32947 11717 32948
rect 12206 32333 12266 35850
rect 12758 35730 12818 37979
rect 12574 35670 12818 35730
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12574 33285 12634 35670
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12571 33284 12637 33285
rect 12571 33220 12572 33284
rect 12636 33220 12637 33284
rect 12571 33219 12637 33220
rect 12203 32332 12269 32333
rect 12203 32268 12204 32332
rect 12268 32268 12269 32332
rect 12203 32267 12269 32268
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 10182 31710 10978 31770
rect 10182 30701 10242 31710
rect 10179 30700 10245 30701
rect 10179 30636 10180 30700
rect 10244 30636 10245 30700
rect 10179 30635 10245 30636
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 8707 19684 8773 19685
rect 8707 19620 8708 19684
rect 8772 19620 8773 19684
rect 8707 19619 8773 19620
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 5395 18188 5461 18189
rect 5395 18124 5396 18188
rect 5460 18124 5461 18188
rect 5395 18123 5461 18124
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 8710 5813 8770 19619
rect 8707 5812 8773 5813
rect 8707 5748 8708 5812
rect 8772 5748 8773 5812
rect 8707 5747 8773 5748
rect 10182 5677 10242 30635
rect 12019 24036 12085 24037
rect 12019 23972 12020 24036
rect 12084 23972 12085 24036
rect 12019 23971 12085 23972
rect 12022 14109 12082 23971
rect 12206 19413 12266 32267
rect 12203 19412 12269 19413
rect 12203 19348 12204 19412
rect 12268 19348 12269 19412
rect 12203 19347 12269 19348
rect 12574 17917 12634 33219
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 14411 32468 14477 32469
rect 14411 32404 14412 32468
rect 14476 32404 14477 32468
rect 14411 32403 14477 32404
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 14414 21725 14474 32403
rect 15699 29068 15765 29069
rect 15699 29004 15700 29068
rect 15764 29004 15765 29068
rect 15699 29003 15765 29004
rect 14963 28252 15029 28253
rect 14963 28188 14964 28252
rect 15028 28188 15029 28252
rect 14963 28187 15029 28188
rect 14411 21724 14477 21725
rect 14411 21660 14412 21724
rect 14476 21660 14477 21724
rect 14411 21659 14477 21660
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 14779 19684 14845 19685
rect 14779 19620 14780 19684
rect 14844 19620 14845 19684
rect 14779 19619 14845 19620
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12571 17916 12637 17917
rect 12571 17852 12572 17916
rect 12636 17852 12637 17916
rect 12571 17851 12637 17852
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12019 14108 12085 14109
rect 12019 14044 12020 14108
rect 12084 14044 12085 14108
rect 12019 14043 12085 14044
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 10179 5676 10245 5677
rect 10179 5612 10180 5676
rect 10244 5612 10245 5676
rect 10179 5611 10245 5612
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 4928 13264 5952
rect 14782 5133 14842 19619
rect 14966 16285 15026 28187
rect 15147 27300 15213 27301
rect 15147 27236 15148 27300
rect 15212 27236 15213 27300
rect 15147 27235 15213 27236
rect 15150 18325 15210 27235
rect 15147 18324 15213 18325
rect 15147 18260 15148 18324
rect 15212 18260 15213 18324
rect 15147 18259 15213 18260
rect 15702 16285 15762 29003
rect 15886 28253 15946 40019
rect 16070 38725 16130 43011
rect 16067 38724 16133 38725
rect 16067 38660 16068 38724
rect 16132 38660 16133 38724
rect 16067 38659 16133 38660
rect 15883 28252 15949 28253
rect 15883 28188 15884 28252
rect 15948 28188 15949 28252
rect 15883 28187 15949 28188
rect 16070 21997 16130 38659
rect 16251 36956 16317 36957
rect 16251 36892 16252 36956
rect 16316 36892 16317 36956
rect 16251 36891 16317 36892
rect 16254 29205 16314 36891
rect 16251 29204 16317 29205
rect 16251 29140 16252 29204
rect 16316 29140 16317 29204
rect 16251 29139 16317 29140
rect 16438 29069 16498 52531
rect 16435 29068 16501 29069
rect 16435 29004 16436 29068
rect 16500 29004 16501 29068
rect 16435 29003 16501 29004
rect 16803 28388 16869 28389
rect 16803 28324 16804 28388
rect 16868 28324 16869 28388
rect 16803 28323 16869 28324
rect 16251 27980 16317 27981
rect 16251 27916 16252 27980
rect 16316 27916 16317 27980
rect 16251 27915 16317 27916
rect 16067 21996 16133 21997
rect 16067 21932 16068 21996
rect 16132 21932 16133 21996
rect 16067 21931 16133 21932
rect 16070 20773 16130 21931
rect 16067 20772 16133 20773
rect 16067 20708 16068 20772
rect 16132 20708 16133 20772
rect 16067 20707 16133 20708
rect 16254 16829 16314 27915
rect 16806 25261 16866 28323
rect 17174 27437 17234 52531
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 23795 52596 23861 52597
rect 23795 52532 23796 52596
rect 23860 52532 23861 52596
rect 23795 52531 23861 52532
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 18643 47700 18709 47701
rect 18643 47636 18644 47700
rect 18708 47636 18709 47700
rect 18643 47635 18709 47636
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17355 39948 17421 39949
rect 17355 39884 17356 39948
rect 17420 39884 17421 39948
rect 17355 39883 17421 39884
rect 17171 27436 17237 27437
rect 17171 27372 17172 27436
rect 17236 27372 17237 27436
rect 17171 27371 17237 27372
rect 16803 25260 16869 25261
rect 16803 25196 16804 25260
rect 16868 25196 16869 25260
rect 16803 25195 16869 25196
rect 17358 20637 17418 39883
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 18646 38861 18706 47635
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 21771 47020 21837 47021
rect 21771 46956 21772 47020
rect 21836 46956 21837 47020
rect 21771 46955 21837 46956
rect 20115 45932 20181 45933
rect 20115 45868 20116 45932
rect 20180 45868 20181 45932
rect 20115 45867 20181 45868
rect 19747 43212 19813 43213
rect 19747 43148 19748 43212
rect 19812 43148 19813 43212
rect 19747 43147 19813 43148
rect 19195 40084 19261 40085
rect 19195 40020 19196 40084
rect 19260 40020 19261 40084
rect 19195 40019 19261 40020
rect 18643 38860 18709 38861
rect 18643 38796 18644 38860
rect 18708 38796 18709 38860
rect 18643 38795 18709 38796
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17355 20636 17421 20637
rect 17355 20572 17356 20636
rect 17420 20572 17421 20636
rect 17355 20571 17421 20572
rect 17944 19616 18264 20640
rect 18646 19957 18706 38795
rect 19198 33149 19258 40019
rect 19750 38453 19810 43147
rect 19747 38452 19813 38453
rect 19747 38388 19748 38452
rect 19812 38388 19813 38452
rect 19747 38387 19813 38388
rect 19195 33148 19261 33149
rect 19195 33084 19196 33148
rect 19260 33084 19261 33148
rect 19195 33083 19261 33084
rect 19563 31924 19629 31925
rect 19563 31860 19564 31924
rect 19628 31860 19629 31924
rect 19563 31859 19629 31860
rect 19566 20637 19626 31859
rect 19750 30837 19810 38387
rect 20118 31245 20178 45867
rect 21587 43076 21653 43077
rect 21587 43012 21588 43076
rect 21652 43012 21653 43076
rect 21587 43011 21653 43012
rect 20115 31244 20181 31245
rect 20115 31180 20116 31244
rect 20180 31180 20181 31244
rect 20115 31179 20181 31180
rect 19747 30836 19813 30837
rect 19747 30772 19748 30836
rect 19812 30772 19813 30836
rect 19747 30771 19813 30772
rect 19747 27844 19813 27845
rect 19747 27780 19748 27844
rect 19812 27780 19813 27844
rect 19747 27779 19813 27780
rect 19750 20773 19810 27779
rect 19747 20772 19813 20773
rect 19747 20708 19748 20772
rect 19812 20708 19813 20772
rect 19747 20707 19813 20708
rect 19563 20636 19629 20637
rect 19563 20572 19564 20636
rect 19628 20572 19629 20636
rect 19563 20571 19629 20572
rect 18643 19956 18709 19957
rect 18643 19892 18644 19956
rect 18708 19892 18709 19956
rect 18643 19891 18709 19892
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 18459 19412 18525 19413
rect 18459 19348 18460 19412
rect 18524 19348 18525 19412
rect 18459 19347 18525 19348
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 16251 16828 16317 16829
rect 16251 16764 16252 16828
rect 16316 16764 16317 16828
rect 16251 16763 16317 16764
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 14963 16284 15029 16285
rect 14963 16220 14964 16284
rect 15028 16220 15029 16284
rect 14963 16219 15029 16220
rect 15699 16284 15765 16285
rect 15699 16220 15700 16284
rect 15764 16220 15765 16284
rect 15699 16219 15765 16220
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 14779 5132 14845 5133
rect 14779 5068 14780 5132
rect 14844 5068 14845 5132
rect 14779 5067 14845 5068
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 18462 4045 18522 19347
rect 20118 18733 20178 31179
rect 20483 29068 20549 29069
rect 20483 29004 20484 29068
rect 20548 29004 20549 29068
rect 20483 29003 20549 29004
rect 20486 20773 20546 29003
rect 21590 28525 21650 43011
rect 21774 31789 21834 46955
rect 22691 46612 22757 46613
rect 22691 46548 22692 46612
rect 22756 46548 22757 46612
rect 22691 46547 22757 46548
rect 21955 45932 22021 45933
rect 21955 45868 21956 45932
rect 22020 45868 22021 45932
rect 21955 45867 22021 45868
rect 21771 31788 21837 31789
rect 21771 31724 21772 31788
rect 21836 31724 21837 31788
rect 21771 31723 21837 31724
rect 21958 30293 22018 45867
rect 22507 36684 22573 36685
rect 22507 36620 22508 36684
rect 22572 36620 22573 36684
rect 22507 36619 22573 36620
rect 22510 33013 22570 36619
rect 22507 33012 22573 33013
rect 22507 32948 22508 33012
rect 22572 32948 22573 33012
rect 22507 32947 22573 32948
rect 21955 30292 22021 30293
rect 21955 30228 21956 30292
rect 22020 30228 22021 30292
rect 21955 30227 22021 30228
rect 21587 28524 21653 28525
rect 21587 28460 21588 28524
rect 21652 28460 21653 28524
rect 21587 28459 21653 28460
rect 22694 28389 22754 46547
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 23798 32605 23858 52531
rect 23795 32604 23861 32605
rect 23795 32540 23796 32604
rect 23860 32540 23861 32604
rect 23795 32539 23861 32540
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22691 28388 22757 28389
rect 22691 28324 22692 28388
rect 22756 28324 22757 28388
rect 22691 28323 22757 28324
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 20483 20772 20549 20773
rect 20483 20708 20484 20772
rect 20548 20708 20549 20772
rect 20483 20707 20549 20708
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 20115 18732 20181 18733
rect 20115 18668 20116 18732
rect 20180 18668 20181 18732
rect 20115 18667 20181 18668
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 18459 4044 18525 4045
rect 18459 3980 18460 4044
rect 18524 3980 18525 4044
rect 18459 3979 18525 3980
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _109_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1679235063
transform 1 0 24564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _111_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1679235063
transform 1 0 23736 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1679235063
transform 1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1679235063
transform 1 0 24656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1679235063
transform 1 0 24564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1679235063
transform 1 0 16008 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1679235063
transform 1 0 23184 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1679235063
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1679235063
transform 1 0 20700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform 1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 21160 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1679235063
transform 1 0 21160 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1679235063
transform 1 0 23276 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1679235063
transform 1 0 21160 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1679235063
transform 1 0 24656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1679235063
transform 1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1679235063
transform 1 0 21896 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1679235063
transform 1 0 23184 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1679235063
transform 1 0 23736 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1679235063
transform 1 0 24564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1679235063
transform 1 0 24564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1679235063
transform 1 0 24564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1679235063
transform 1 0 24564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1679235063
transform 1 0 25024 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1679235063
transform 1 0 24564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1679235063
transform 1 0 22172 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1679235063
transform 1 0 13340 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1679235063
transform 1 0 14076 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform 1 0 13616 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform 1 0 15824 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1679235063
transform 1 0 16836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1679235063
transform 1 0 15272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1679235063
transform 1 0 15548 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1679235063
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1679235063
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1679235063
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1679235063
transform 1 0 17112 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1679235063
transform 1 0 16836 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1679235063
transform 1 0 18400 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1679235063
transform 1 0 18492 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 19504 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform 1 0 20608 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1679235063
transform 1 0 19596 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 20332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1679235063
transform 1 0 21068 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1679235063
transform 1 0 19044 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1679235063
transform 1 0 18676 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1679235063
transform 1 0 20792 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1679235063
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1679235063
transform 1 0 21068 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1679235063
transform 1 0 20240 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1679235063
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1679235063
transform 1 0 3128 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1679235063
transform 1 0 4876 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1679235063
transform 1 0 4140 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1679235063
transform 1 0 6716 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _172_
timestamp 1679235063
transform 1 0 4692 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1679235063
transform 1 0 4968 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1679235063
transform 1 0 6532 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1679235063
transform 1 0 6808 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1679235063
transform 1 0 6624 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1679235063
transform 1 0 6532 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1679235063
transform 1 0 7268 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _179_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7452 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1679235063
transform 1 0 7636 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1679235063
transform 1 0 7912 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1679235063
transform 1 0 8832 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1679235063
transform 1 0 6808 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1679235063
transform 1 0 9108 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1679235063
transform 1 0 8372 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1679235063
transform 1 0 10396 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1679235063
transform 1 0 9200 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1679235063
transform 1 0 11408 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1679235063
transform 1 0 10856 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1679235063
transform 1 0 11408 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1679235063
transform 1 0 9016 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1679235063
transform 1 0 9292 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1679235063
transform 1 0 12236 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1679235063
transform 1 0 10212 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1679235063
transform 1 0 11684 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1679235063
transform 1 0 12604 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1679235063
transform 1 0 12328 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1679235063
transform 1 0 2392 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1679235063
transform 1 0 2024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1679235063
transform 1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1679235063
transform 1 0 2024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1679235063
transform 1 0 2024 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1679235063
transform 1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1679235063
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1679235063
transform 1 0 2024 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 12696 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform -1 0 11408 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 11960 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1679235063
transform 1 0 13708 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1679235063
transform 1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1679235063
transform 1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1679235063
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1679235063
transform 1 0 14904 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1679235063
transform 1 0 17388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1679235063
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1679235063
transform 1 0 16100 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1679235063
transform 1 0 17204 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1679235063
transform 1 0 17112 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1679235063
transform 1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1679235063
transform 1 0 18952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1679235063
transform 1 0 18124 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1679235063
transform 1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1679235063
transform 1 0 20700 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1679235063
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A
timestamp 1679235063
transform 1 0 19596 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 1679235063
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A
timestamp 1679235063
transform 1 0 3680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A
timestamp 1679235063
transform 1 0 5428 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1679235063
transform 1 0 3772 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1679235063
transform 1 0 5244 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1679235063
transform 1 0 5520 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1679235063
transform 1 0 7084 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1679235063
transform 1 0 7176 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1679235063
transform 1 0 6348 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A
timestamp 1679235063
transform 1 0 7084 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1679235063
transform 1 0 8188 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1679235063
transform 1 0 8464 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1679235063
transform 1 0 9384 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1679235063
transform 1 0 9660 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1679235063
transform 1 0 8188 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1679235063
transform 1 0 10212 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1679235063
transform 1 0 11960 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1679235063
transform 1 0 11500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1679235063
transform 1 0 11040 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1679235063
transform 1 0 12052 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 6532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 9384 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11868 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 7728 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14904 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11960 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 10028 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 10672 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12972 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__CLK
timestamp 1679235063
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 8464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 7820 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 15088 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13524 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 13892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 14720 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 13800 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 12420 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 12604 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 11040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 8556 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 12144 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16008 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 14628 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 13708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 12420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 13708 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15088 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 15272 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16192 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 12420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 12604 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 13156 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10028 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 11040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 8556 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 9936 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13156 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 15272 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 13616 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 11776 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 12052 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 10396 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 3956 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 5704 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 2576 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6624 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 4324 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 5980 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
timestamp 1679235063
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 16652 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform 1 0 9200 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 17112 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform 1 0 21528 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform 1 0 17480 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 20332 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 10304 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 10672 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 13156 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 19228 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 21068 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform 1 0 18492 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold6_A
timestamp 1679235063
transform 1 0 23828 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold7_A
timestamp 1679235063
transform 1 0 23368 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold12_A
timestamp 1679235063
transform 1 0 4968 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold13_A
timestamp 1679235063
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold15_A
timestamp 1679235063
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold17_A
timestamp 1679235063
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold19_A
timestamp 1679235063
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold21_A
timestamp 1679235063
transform 1 0 17756 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold22_A
timestamp 1679235063
transform 1 0 14812 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold23_A
timestamp 1679235063
transform 1 0 19872 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold24_A
timestamp 1679235063
transform 1 0 17388 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold25_A
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold26_A
timestamp 1679235063
transform 1 0 21436 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold27_A
timestamp 1679235063
transform 1 0 18584 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold28_A
timestamp 1679235063
transform 1 0 14260 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold29_A
timestamp 1679235063
transform 1 0 7084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold30_A
timestamp 1679235063
transform 1 0 18768 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold31_A
timestamp 1679235063
transform 1 0 14444 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold32_A
timestamp 1679235063
transform 1 0 17572 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold33_A
timestamp 1679235063
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold34_A
timestamp 1679235063
transform 1 0 15180 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold35_A
timestamp 1679235063
transform 1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold36_A
timestamp 1679235063
transform 1 0 25116 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold37_A
timestamp 1679235063
transform 1 0 4600 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold38_A
timestamp 1679235063
transform 1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold39_A
timestamp 1679235063
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold40_A
timestamp 1679235063
transform 1 0 7268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold41_A
timestamp 1679235063
transform 1 0 18860 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold42_A
timestamp 1679235063
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold43_A
timestamp 1679235063
transform 1 0 16376 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold44_A
timestamp 1679235063
transform 1 0 18952 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold45_A
timestamp 1679235063
transform 1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold46_A
timestamp 1679235063
transform 1 0 24012 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold47_A
timestamp 1679235063
transform 1 0 25116 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold48_A
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold49_A
timestamp 1679235063
transform 1 0 21436 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold50_A
timestamp 1679235063
transform 1 0 4784 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold51_A
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold52_A
timestamp 1679235063
transform 1 0 10488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold53_A
timestamp 1679235063
transform 1 0 6440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold54_A
timestamp 1679235063
transform 1 0 7544 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold55_A
timestamp 1679235063
transform 1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold56_A
timestamp 1679235063
transform 1 0 10304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold57_A
timestamp 1679235063
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold58_A
timestamp 1679235063
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold59_A
timestamp 1679235063
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold60_A
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold61_A
timestamp 1679235063
transform 1 0 3956 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold64_A
timestamp 1679235063
transform 1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform 1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 25208 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 24748 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 24472 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 24748 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 24564 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 25392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 25208 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 25392 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 24748 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform 1 0 24748 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform 1 0 24748 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform 1 0 25392 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 23552 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 25392 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 25208 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 24748 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 24748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 24748 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 24748 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 10764 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 12144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1679235063
transform 1 0 11500 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1679235063
transform 1 0 17848 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform 1 0 19320 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform 1 0 20792 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1679235063
transform 1 0 22816 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1679235063
transform 1 0 25300 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1679235063
transform 1 0 23552 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1679235063
transform 1 0 23736 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1679235063
transform 1 0 24380 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1679235063
transform 1 0 14904 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1679235063
transform 1 0 16376 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1679235063
transform 1 0 24656 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1679235063
transform 1 0 24656 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1679235063
transform 1 0 24472 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1679235063
transform 1 0 25392 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1679235063
transform 1 0 24656 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1679235063
transform 1 0 24656 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1679235063
transform 1 0 23920 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1679235063
transform 1 0 24104 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1679235063
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1679235063
transform 1 0 2116 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1679235063
transform 1 0 5060 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1679235063
transform 1 0 3772 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1679235063
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1679235063
transform 1 0 3220 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output145_A
timestamp 1679235063
transform 1 0 18492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output146_A
timestamp 1679235063
transform 1 0 18492 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18492 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 16100 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16284 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 16284 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18492 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21436 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21896 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 22264 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21436 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21068 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 17388 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 17572 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 17940 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20884 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21436 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 23828 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25116 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 25116 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24104 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18216 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 15824 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17112 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16100 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 14904 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17940 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21712 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 20424 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17388 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20792 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24012 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 25392 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 24748 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24564 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 25392 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25300 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23920 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 25208 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24656 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 23736 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 24380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24012 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21344 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21252 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 20332 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20424 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21068 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 18860 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18676 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 17664 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 17112 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16376 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16376 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 15640 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14904 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12420 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 11592 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13248 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14352 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14720 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13156 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11776 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10304 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9752 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8556 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8188 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8372 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8464 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10304 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 8372 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 9108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17388 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18860 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19688 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21712 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24012 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23736 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22908 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21528 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20240 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 6532 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 11500 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 8832 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 9844 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 12236 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 15180 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15364 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 14168 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14260 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 13156 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12972 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 10948 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 10580 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11500 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 8648 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 10488 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 7268 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8648 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 7728 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 7544 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8464 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8464 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 7084 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10304 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 9016 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 10856 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10120 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8096 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 5980 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 7084 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 6900 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 8004 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8188 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1679235063
transform 1 0 8096 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 7912 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 9292 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9476 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12788 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18860 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 18032 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16836 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17020 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 19228 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19044 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 17848 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 12328 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 11592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 12972 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18860 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20056 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 20424 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 16836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19688 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21068 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23000 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 19872 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17480 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18676 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21436 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18124 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 16468 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16744 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18124 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 17940 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 20240 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 18216 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 18032 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 13064 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 14444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18584 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18768 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21528 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 17204 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20516 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20700 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23276 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 19688 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15732 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17296 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 20976 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18032 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18768 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18584 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 13064 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_45.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20424 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15916 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16008 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 10856 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23276 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 22816 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 22632 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23460 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 23276 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 22448 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 22264 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 22264 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 21252 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 21620 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 21436 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23000 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 23920 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24104 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 19412 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 23184 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23000 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 20608 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 21252 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21620 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 22080 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21896 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 18584 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 20608 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21896 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 20976 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 20792 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 15732 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19320 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 20240 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 19044 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19044 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 17848 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 13800 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17664 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 17204 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 12328 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15640 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 14168 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 11592 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13616 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 10028 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16284 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16100 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 12696 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17848 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 11040 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16100 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15088 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 8832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 8556 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12420 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12236 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 7268 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15916 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15272 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12880 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12512 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 6900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16008 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17204 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17296 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18308 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20240 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23276 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 23092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20056 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21068 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_54.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16928 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18308 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8556 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 9108 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 8924 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18308 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 18124 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 13984 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 15548 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 8832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 9016 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18032 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 17848 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 18400 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 12144 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 12328 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 13892 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16192 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14812 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 14628 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 10580 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 10764 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 12144 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8464 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 8648 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 10212 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 18216 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 13616 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 8464 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 9660 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8096 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 8280 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 8464 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 17848 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 12236 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 12420 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 7084 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 8280 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12512 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11776 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 7268 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 7452 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15732 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14536 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 14352 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 18308 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 8924 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 9108 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13156 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 12512 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 4600 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12236 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11040 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 12880 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 7452 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16652 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 11500 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_52.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4048 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9752 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6532 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 5704 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9108 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12604 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9936 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 8004 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9108 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11040 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6624 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 5336 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6532 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9752 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 5796 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 4232 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11684 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 8740 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__256 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 11316 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9936 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform 1 0 8280 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform 1 0 7084 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15640 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 15272 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14812 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 14260 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 11408 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform 1 0 10120 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__257
timestamp 1679235063
transform 1 0 13248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 12052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10488 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10028 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15456 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14444 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14352 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 12972 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10396 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12328 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11776 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 8740 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__258
timestamp 1679235063
transform 1 0 11868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 8924 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 7452 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform 1 0 6256 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4692 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13524 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14260 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 11960 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11684 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 7820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__259
timestamp 1679235063
transform 1 0 9844 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9476 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 6808 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4048 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3956 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4140 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 3680 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 4232 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 3036 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 2944 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 2760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 3956 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 4232 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 3956 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 4508 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 3404 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 3956 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_4  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 3680 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 9016 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9844 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14720 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 8464 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform 1 0 10488 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform 1 0 8004 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 9936 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform 1 0 17480 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 20332 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform 1 0 17848 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 20516 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform 1 0 9108 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform 1 0 10212 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 9292 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 11960 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform 1 0 19412 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 21436 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform 1 0 18860 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform 1 0 21988 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35
timestamp 1679235063
transform 1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49
timestamp 1679235063
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1679235063
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1679235063
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1679235063
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1679235063
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1679235063
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1679235063
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1679235063
transform 1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1679235063
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1679235063
transform 1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1679235063
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1679235063
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1679235063
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1679235063
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1679235063
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_263
timestamp 1679235063
transform 1 0 25300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1679235063
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1679235063
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_33
timestamp 1679235063
transform 1 0 4140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_37
timestamp 1679235063
transform 1 0 4508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_42
timestamp 1679235063
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1679235063
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_60
timestamp 1679235063
transform 1 0 6624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_70
timestamp 1679235063
transform 1 0 7544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1679235063
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1679235063
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1679235063
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1679235063
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1679235063
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1679235063
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1679235063
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1679235063
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_207 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1679235063
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1679235063
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_225 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_231
timestamp 1679235063
transform 1 0 22356 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1679235063
transform 1 0 23184 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_244
timestamp 1679235063
transform 1 0 23552 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_256
timestamp 1679235063
transform 1 0 24656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_260
timestamp 1679235063
transform 1 0 25024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1679235063
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1679235063
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1679235063
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_34
timestamp 1679235063
transform 1 0 4232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_46
timestamp 1679235063
transform 1 0 5336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1679235063
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1679235063
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1679235063
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_91
timestamp 1679235063
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_103
timestamp 1679235063
transform 1 0 10580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1679235063
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1679235063
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1679235063
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1679235063
transform 1 0 14812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1679235063
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1679235063
transform 1 0 18308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1679235063
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1679235063
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1679235063
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_235
timestamp 1679235063
transform 1 0 22724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_241
timestamp 1679235063
transform 1 0 23276 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1679235063
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_263
timestamp 1679235063
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1679235063
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_19
timestamp 1679235063
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1679235063
transform 1 0 3312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp 1679235063
transform 1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1679235063
transform 1 0 5152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1679235063
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_67
timestamp 1679235063
transform 1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_72
timestamp 1679235063
transform 1 0 7728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1679235063
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1679235063
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1679235063
transform 1 0 10120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_104
timestamp 1679235063
transform 1 0 10672 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_107
timestamp 1679235063
transform 1 0 10948 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_123
timestamp 1679235063
transform 1 0 12420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_151
timestamp 1679235063
transform 1 0 14996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_159
timestamp 1679235063
transform 1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1679235063
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1679235063
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1679235063
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1679235063
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1679235063
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1679235063
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_247
timestamp 1679235063
transform 1 0 23828 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1679235063
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1679235063
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1679235063
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_35
timestamp 1679235063
transform 1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_39
timestamp 1679235063
transform 1 0 4692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_46
timestamp 1679235063
transform 1 0 5336 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_54
timestamp 1679235063
transform 1 0 6072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_58
timestamp 1679235063
transform 1 0 6440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp 1679235063
transform 1 0 6900 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_67
timestamp 1679235063
transform 1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_74
timestamp 1679235063
transform 1 0 7912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1679235063
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1679235063
transform 1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_96
timestamp 1679235063
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_102
timestamp 1679235063
transform 1 0 10488 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_114
timestamp 1679235063
transform 1 0 11592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_118
timestamp 1679235063
transform 1 0 11960 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_122
timestamp 1679235063
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1679235063
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1679235063
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1679235063
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_177
timestamp 1679235063
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1679235063
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1679235063
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_235
timestamp 1679235063
transform 1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1679235063
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_259
timestamp 1679235063
transform 1 0 24932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1679235063
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_5
timestamp 1679235063
transform 1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1679235063
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_31
timestamp 1679235063
transform 1 0 3956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1679235063
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_46
timestamp 1679235063
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_65
timestamp 1679235063
transform 1 0 7084 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1679235063
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1679235063
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1679235063
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1679235063
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1679235063
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1679235063
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1679235063
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1679235063
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1679235063
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1679235063
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1679235063
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_11
timestamp 1679235063
transform 1 0 2116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_23
timestamp 1679235063
transform 1 0 3220 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_33
timestamp 1679235063
transform 1 0 4140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_45
timestamp 1679235063
transform 1 0 5244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_57
timestamp 1679235063
transform 1 0 6348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_69
timestamp 1679235063
transform 1 0 7452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1679235063
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1679235063
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1679235063
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1679235063
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1679235063
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1679235063
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_177
timestamp 1679235063
transform 1 0 17388 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1679235063
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_209
timestamp 1679235063
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_227
timestamp 1679235063
transform 1 0 21988 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1679235063
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1679235063
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1679235063
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1679235063
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_10
timestamp 1679235063
transform 1 0 2024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1679235063
transform 1 0 2668 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_29
timestamp 1679235063
transform 1 0 3772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_41
timestamp 1679235063
transform 1 0 4876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1679235063
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1679235063
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1679235063
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1679235063
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1679235063
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1679235063
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1679235063
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1679235063
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1679235063
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 1679235063
transform 1 0 17756 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1679235063
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1679235063
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1679235063
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_243
timestamp 1679235063
transform 1 0 23460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_247
timestamp 1679235063
transform 1 0 23828 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1679235063
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1679235063
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1679235063
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1679235063
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1679235063
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1679235063
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1679235063
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1679235063
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1679235063
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1679235063
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1679235063
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1679235063
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1679235063
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1679235063
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1679235063
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1679235063
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_203
timestamp 1679235063
transform 1 0 19780 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_207
timestamp 1679235063
transform 1 0 20148 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1679235063
transform 1 0 20700 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1679235063
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1679235063
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_259
timestamp 1679235063
transform 1 0 24932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1679235063
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1679235063
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1679235063
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1679235063
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1679235063
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1679235063
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1679235063
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1679235063
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1679235063
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1679235063
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1679235063
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1679235063
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1679235063
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1679235063
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1679235063
transform 1 0 18492 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_195
timestamp 1679235063
transform 1 0 19044 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_203
timestamp 1679235063
transform 1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1679235063
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1679235063
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1679235063
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1679235063
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_55
timestamp 1679235063
transform 1 0 6164 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_61
timestamp 1679235063
transform 1 0 6716 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_73
timestamp 1679235063
transform 1 0 7820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1679235063
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1679235063
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1679235063
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1679235063
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1679235063
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1679235063
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1679235063
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1679235063
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1679235063
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1679235063
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1679235063
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_205
timestamp 1679235063
transform 1 0 19964 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_211
timestamp 1679235063
transform 1 0 20516 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_220
timestamp 1679235063
transform 1 0 21344 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_232
timestamp 1679235063
transform 1 0 22448 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1679235063
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_258
timestamp 1679235063
transform 1 0 24840 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1679235063
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1679235063
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1679235063
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1679235063
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1679235063
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1679235063
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1679235063
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1679235063
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1679235063
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1679235063
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1679235063
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1679235063
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1679235063
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1679235063
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1679235063
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_199
timestamp 1679235063
transform 1 0 19412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_203
timestamp 1679235063
transform 1 0 19780 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_211
timestamp 1679235063
transform 1 0 20516 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 1679235063
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1679235063
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1679235063
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1679235063
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1679235063
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1679235063
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1679235063
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1679235063
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1679235063
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1679235063
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1679235063
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1679235063
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1679235063
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1679235063
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1679235063
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1679235063
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1679235063
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1679235063
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1679235063
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1679235063
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1679235063
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_221
timestamp 1679235063
transform 1 0 21436 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_225
timestamp 1679235063
transform 1 0 21804 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_237
timestamp 1679235063
transform 1 0 22908 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_245
timestamp 1679235063
transform 1 0 23644 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1679235063
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_259
timestamp 1679235063
transform 1 0 24932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1679235063
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1679235063
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1679235063
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1679235063
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_68
timestamp 1679235063
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_80
timestamp 1679235063
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_92
timestamp 1679235063
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1679235063
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1679235063
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1679235063
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1679235063
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1679235063
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1679235063
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_175
timestamp 1679235063
transform 1 0 17204 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_187
timestamp 1679235063
transform 1 0 18308 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_198
timestamp 1679235063
transform 1 0 19320 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_210
timestamp 1679235063
transform 1 0 20424 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1679235063
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_233
timestamp 1679235063
transform 1 0 22540 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_238
timestamp 1679235063
transform 1 0 23000 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_246
timestamp 1679235063
transform 1 0 23736 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1679235063
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1679235063
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1679235063
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1679235063
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1679235063
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1679235063
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1679235063
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1679235063
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1679235063
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1679235063
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1679235063
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1679235063
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1679235063
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_150
timestamp 1679235063
transform 1 0 14904 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_162
timestamp 1679235063
transform 1 0 16008 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_168
timestamp 1679235063
transform 1 0 16560 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_173
timestamp 1679235063
transform 1 0 17020 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_185
timestamp 1679235063
transform 1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1679235063
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_209
timestamp 1679235063
transform 1 0 20332 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1679235063
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_222
timestamp 1679235063
transform 1 0 21528 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_226
timestamp 1679235063
transform 1 0 21896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1679235063
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1679235063
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_259
timestamp 1679235063
transform 1 0 24932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_265
timestamp 1679235063
transform 1 0 25484 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1679235063
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1679235063
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1679235063
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1679235063
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1679235063
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1679235063
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1679235063
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1679235063
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1679235063
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1679235063
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1679235063
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_122
timestamp 1679235063
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_126
timestamp 1679235063
transform 1 0 12696 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_138
timestamp 1679235063
transform 1 0 13800 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_146
timestamp 1679235063
transform 1 0 14536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_150
timestamp 1679235063
transform 1 0 14904 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_156
timestamp 1679235063
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1679235063
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1679235063
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_189
timestamp 1679235063
transform 1 0 18492 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_195
timestamp 1679235063
transform 1 0 19044 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_205
timestamp 1679235063
transform 1 0 19964 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_212
timestamp 1679235063
transform 1 0 20608 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_237
timestamp 1679235063
transform 1 0 22908 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_243
timestamp 1679235063
transform 1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_247
timestamp 1679235063
transform 1 0 23828 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1679235063
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1679235063
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1679235063
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1679235063
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1679235063
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1679235063
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1679235063
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1679235063
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1679235063
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1679235063
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1679235063
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1679235063
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1679235063
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1679235063
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1679235063
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_155
timestamp 1679235063
transform 1 0 15364 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1679235063
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1679235063
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1679235063
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1679235063
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_204
timestamp 1679235063
transform 1 0 19872 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_212
timestamp 1679235063
transform 1 0 20608 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_217
timestamp 1679235063
transform 1 0 21068 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_229
timestamp 1679235063
transform 1 0 22172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_241
timestamp 1679235063
transform 1 0 23276 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1679235063
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_265
timestamp 1679235063
transform 1 0 25484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1679235063
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1679235063
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1679235063
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1679235063
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1679235063
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1679235063
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1679235063
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1679235063
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1679235063
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1679235063
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1679235063
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1679235063
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_160
timestamp 1679235063
transform 1 0 15824 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1679235063
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1679235063
transform 1 0 17204 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_179
timestamp 1679235063
transform 1 0 17572 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1679235063
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp 1679235063
transform 1 0 20056 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1679235063
transform 1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1679235063
transform 1 0 21160 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1679235063
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_237
timestamp 1679235063
transform 1 0 22908 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_257
timestamp 1679235063
transform 1 0 24748 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_265
timestamp 1679235063
transform 1 0 25484 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1679235063
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1679235063
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1679235063
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1679235063
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1679235063
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1679235063
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1679235063
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1679235063
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1679235063
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_133
timestamp 1679235063
transform 1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1679235063
transform 1 0 15272 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_167
timestamp 1679235063
transform 1 0 16468 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_173
timestamp 1679235063
transform 1 0 17020 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_199
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_207
timestamp 1679235063
transform 1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 1679235063
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_226
timestamp 1679235063
transform 1 0 21896 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1679235063
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_244
timestamp 1679235063
transform 1 0 23552 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_265
timestamp 1679235063
transform 1 0 25484 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1679235063
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1679235063
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1679235063
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1679235063
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_69
timestamp 1679235063
transform 1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_86
timestamp 1679235063
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_115
timestamp 1679235063
transform 1 0 11684 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_127
timestamp 1679235063
transform 1 0 12788 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_131
timestamp 1679235063
transform 1 0 13156 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_134
timestamp 1679235063
transform 1 0 13432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1679235063
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_148
timestamp 1679235063
transform 1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1679235063
transform 1 0 15088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_158
timestamp 1679235063
transform 1 0 15640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_164
timestamp 1679235063
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_180
timestamp 1679235063
transform 1 0 17664 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_192
timestamp 1679235063
transform 1 0 18768 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_196
timestamp 1679235063
transform 1 0 19136 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_244
timestamp 1679235063
transform 1 0 23552 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_264
timestamp 1679235063
transform 1 0 25392 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1679235063
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1679235063
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1679235063
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1679235063
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_61
timestamp 1679235063
transform 1 0 6716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1679235063
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_89
timestamp 1679235063
transform 1 0 9292 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1679235063
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_120
timestamp 1679235063
transform 1 0 12144 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1679235063
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1679235063
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1679235063
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1679235063
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1679235063
transform 1 0 16376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_170
timestamp 1679235063
transform 1 0 16744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_174
timestamp 1679235063
transform 1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1679235063
transform 1 0 17572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1679235063
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1679235063
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_212
timestamp 1679235063
transform 1 0 20608 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_215
timestamp 1679235063
transform 1 0 20884 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_221
timestamp 1679235063
transform 1 0 21436 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_224
timestamp 1679235063
transform 1 0 21712 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1679235063
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1679235063
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1679235063
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1679235063
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1679235063
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_69
timestamp 1679235063
transform 1 0 7452 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_95
timestamp 1679235063
transform 1 0 9844 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_99
timestamp 1679235063
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1679235063
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_119
timestamp 1679235063
transform 1 0 12052 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_130
timestamp 1679235063
transform 1 0 13064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_138
timestamp 1679235063
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_142
timestamp 1679235063
transform 1 0 14168 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_154
timestamp 1679235063
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1679235063
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_194
timestamp 1679235063
transform 1 0 18952 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_198
timestamp 1679235063
transform 1 0 19320 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_205
timestamp 1679235063
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_213
timestamp 1679235063
transform 1 0 20700 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1679235063
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_227
timestamp 1679235063
transform 1 0 21988 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_235
timestamp 1679235063
transform 1 0 22724 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_241
timestamp 1679235063
transform 1 0 23276 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_247
timestamp 1679235063
transform 1 0 23828 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1679235063
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1679235063
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1679235063
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1679235063
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1679235063
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1679235063
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1679235063
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1679235063
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1679235063
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1679235063
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_120
timestamp 1679235063
transform 1 0 12144 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_127
timestamp 1679235063
transform 1 0 12788 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_147
timestamp 1679235063
transform 1 0 14628 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1679235063
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_179
timestamp 1679235063
transform 1 0 17572 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_187
timestamp 1679235063
transform 1 0 18308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1679235063
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_202
timestamp 1679235063
transform 1 0 19688 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_207
timestamp 1679235063
transform 1 0 20148 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_235
timestamp 1679235063
transform 1 0 22724 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_239
timestamp 1679235063
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1679235063
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1679235063
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1679235063
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1679235063
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1679235063
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1679235063
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1679235063
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1679235063
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_81
timestamp 1679235063
transform 1 0 8556 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_115
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1679235063
transform 1 0 12420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1679235063
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1679235063
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_151
timestamp 1679235063
transform 1 0 14996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1679235063
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_161
timestamp 1679235063
transform 1 0 15916 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1679235063
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1679235063
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_178
timestamp 1679235063
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_182
timestamp 1679235063
transform 1 0 17848 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1679235063
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_204
timestamp 1679235063
transform 1 0 19872 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_208
timestamp 1679235063
transform 1 0 20240 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1679235063
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_229
timestamp 1679235063
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_233
timestamp 1679235063
transform 1 0 22540 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_239
timestamp 1679235063
transform 1 0 23092 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_243
timestamp 1679235063
transform 1 0 23460 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_247
timestamp 1679235063
transform 1 0 23828 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1679235063
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1679235063
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1679235063
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1679235063
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1679235063
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1679235063
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_77
timestamp 1679235063
transform 1 0 8188 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1679235063
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_100
timestamp 1679235063
transform 1 0 10304 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_106
timestamp 1679235063
transform 1 0 10856 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_129
timestamp 1679235063
transform 1 0 12972 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1679235063
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_152
timestamp 1679235063
transform 1 0 15088 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_164
timestamp 1679235063
transform 1 0 16192 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_174
timestamp 1679235063
transform 1 0 17112 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_185
timestamp 1679235063
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1679235063
transform 1 0 18492 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_208
timestamp 1679235063
transform 1 0 20240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1679235063
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1679235063
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_223
timestamp 1679235063
transform 1 0 21620 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_228
timestamp 1679235063
transform 1 0 22080 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_265
timestamp 1679235063
transform 1 0 25484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_11
timestamp 1679235063
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_18
timestamp 1679235063
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_30
timestamp 1679235063
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_42
timestamp 1679235063
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1679235063
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_80
timestamp 1679235063
transform 1 0 8464 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_84
timestamp 1679235063
transform 1 0 8832 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_94
timestamp 1679235063
transform 1 0 9752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1679235063
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1679235063
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_124
timestamp 1679235063
transform 1 0 12512 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_128
timestamp 1679235063
transform 1 0 12880 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_131
timestamp 1679235063
transform 1 0 13156 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1679235063
transform 1 0 13892 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_145
timestamp 1679235063
transform 1 0 14444 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1679235063
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_157
timestamp 1679235063
transform 1 0 15548 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_164
timestamp 1679235063
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_191
timestamp 1679235063
transform 1 0 18676 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_195
timestamp 1679235063
transform 1 0 19044 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1679235063
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_213
timestamp 1679235063
transform 1 0 20700 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_217
timestamp 1679235063
transform 1 0 21068 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1679235063
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_240
timestamp 1679235063
transform 1 0 23184 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_244
timestamp 1679235063
transform 1 0 23552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1679235063
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1679235063
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1679235063
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1679235063
transform 1 0 4876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_45
timestamp 1679235063
transform 1 0 5244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_66
timestamp 1679235063
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_72
timestamp 1679235063
transform 1 0 7728 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_96
timestamp 1679235063
transform 1 0 9936 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_100
timestamp 1679235063
transform 1 0 10304 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_111
timestamp 1679235063
transform 1 0 11316 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_115
timestamp 1679235063
transform 1 0 11684 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_125
timestamp 1679235063
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1679235063
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_149
timestamp 1679235063
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_152
timestamp 1679235063
transform 1 0 15088 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1679235063
transform 1 0 16100 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_167
timestamp 1679235063
transform 1 0 16468 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_179
timestamp 1679235063
transform 1 0 17572 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1679235063
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1679235063
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_199
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_205
timestamp 1679235063
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1679235063
transform 1 0 20884 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_223
timestamp 1679235063
transform 1 0 21620 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_244
timestamp 1679235063
transform 1 0 23552 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1679235063
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_265
timestamp 1679235063
transform 1 0 25484 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_15
timestamp 1679235063
transform 1 0 2484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_19
timestamp 1679235063
transform 1 0 2852 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_36
timestamp 1679235063
transform 1 0 4416 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1679235063
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_82
timestamp 1679235063
transform 1 0 8648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_92
timestamp 1679235063
transform 1 0 9568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_96
timestamp 1679235063
transform 1 0 9936 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_106
timestamp 1679235063
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_115
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1679235063
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1679235063
transform 1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_154
timestamp 1679235063
transform 1 0 15272 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1679235063
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_174
timestamp 1679235063
transform 1 0 17112 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_200
timestamp 1679235063
transform 1 0 19504 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_204
timestamp 1679235063
transform 1 0 19872 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_213
timestamp 1679235063
transform 1 0 20700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_217
timestamp 1679235063
transform 1 0 21068 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_244
timestamp 1679235063
transform 1 0 23552 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1679235063
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1679235063
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1679235063
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1679235063
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_53
timestamp 1679235063
transform 1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_65
timestamp 1679235063
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_78
timestamp 1679235063
transform 1 0 8280 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_96
timestamp 1679235063
transform 1 0 9936 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_113
timestamp 1679235063
transform 1 0 11500 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_120
timestamp 1679235063
transform 1 0 12144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1679235063
transform 1 0 12788 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1679235063
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_160
timestamp 1679235063
transform 1 0 15824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_173
timestamp 1679235063
transform 1 0 17020 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1679235063
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1679235063
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1679235063
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_203
timestamp 1679235063
transform 1 0 19780 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_224
timestamp 1679235063
transform 1 0 21712 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_248
timestamp 1679235063
transform 1 0 23920 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_259
timestamp 1679235063
transform 1 0 24932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_265
timestamp 1679235063
transform 1 0 25484 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_15
timestamp 1679235063
transform 1 0 2484 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_21
timestamp 1679235063
transform 1 0 3036 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_38
timestamp 1679235063
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1679235063
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_57
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_65
timestamp 1679235063
transform 1 0 7084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_76
timestamp 1679235063
transform 1 0 8096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1679235063
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_95
timestamp 1679235063
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1679235063
transform 1 0 10212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1679235063
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_124
timestamp 1679235063
transform 1 0 12512 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_132
timestamp 1679235063
transform 1 0 13248 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_141
timestamp 1679235063
transform 1 0 14076 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_152
timestamp 1679235063
transform 1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_156
timestamp 1679235063
transform 1 0 15456 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1679235063
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_176
timestamp 1679235063
transform 1 0 17296 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_189
timestamp 1679235063
transform 1 0 18492 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_213
timestamp 1679235063
transform 1 0 20700 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_217
timestamp 1679235063
transform 1 0 21068 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1679235063
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_227
timestamp 1679235063
transform 1 0 21988 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_245
timestamp 1679235063
transform 1 0 23644 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1679235063
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_261
timestamp 1679235063
transform 1 0 25116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_265
timestamp 1679235063
transform 1 0 25484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1679235063
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1679235063
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_47
timestamp 1679235063
transform 1 0 5428 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_59
timestamp 1679235063
transform 1 0 6532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_71
timestamp 1679235063
transform 1 0 7636 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1679235063
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_87
timestamp 1679235063
transform 1 0 9108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_92
timestamp 1679235063
transform 1 0 9568 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1679235063
transform 1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_121
timestamp 1679235063
transform 1 0 12236 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_152
timestamp 1679235063
transform 1 0 15088 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_185
timestamp 1679235063
transform 1 0 18124 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_191
timestamp 1679235063
transform 1 0 18676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_204
timestamp 1679235063
transform 1 0 19872 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_208
timestamp 1679235063
transform 1 0 20240 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_220
timestamp 1679235063
transform 1 0 21344 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1679235063
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_255
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_263
timestamp 1679235063
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_9
timestamp 1679235063
transform 1 0 1932 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_13
timestamp 1679235063
transform 1 0 2300 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_35
timestamp 1679235063
transform 1 0 4324 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_42
timestamp 1679235063
transform 1 0 4968 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1679235063
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1679235063
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_92
timestamp 1679235063
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_104
timestamp 1679235063
transform 1 0 10672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_124
timestamp 1679235063
transform 1 0 12512 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_130
timestamp 1679235063
transform 1 0 13064 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_133
timestamp 1679235063
transform 1 0 13340 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1679235063
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_150
timestamp 1679235063
transform 1 0 14904 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1679235063
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1679235063
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_187
timestamp 1679235063
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_195
timestamp 1679235063
transform 1 0 19044 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_208
timestamp 1679235063
transform 1 0 20240 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_212
timestamp 1679235063
transform 1 0 20608 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1679235063
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_247
timestamp 1679235063
transform 1 0 23828 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_251
timestamp 1679235063
transform 1 0 24196 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_263
timestamp 1679235063
transform 1 0 25300 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1679235063
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1679235063
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_41
timestamp 1679235063
transform 1 0 4876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_46
timestamp 1679235063
transform 1 0 5336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_70
timestamp 1679235063
transform 1 0 7544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_74
timestamp 1679235063
transform 1 0 7912 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_78
timestamp 1679235063
transform 1 0 8280 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1679235063
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1679235063
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_114
timestamp 1679235063
transform 1 0 11592 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_124
timestamp 1679235063
transform 1 0 12512 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_136
timestamp 1679235063
transform 1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_152
timestamp 1679235063
transform 1 0 15088 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_156
timestamp 1679235063
transform 1 0 15456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_168
timestamp 1679235063
transform 1 0 16560 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_178
timestamp 1679235063
transform 1 0 17480 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_184
timestamp 1679235063
transform 1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_188
timestamp 1679235063
transform 1 0 18400 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1679235063
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_199
timestamp 1679235063
transform 1 0 19412 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_207
timestamp 1679235063
transform 1 0 20148 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_210
timestamp 1679235063
transform 1 0 20424 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_222
timestamp 1679235063
transform 1 0 21528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1679235063
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1679235063
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1679235063
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1679235063
transform 1 0 3588 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_51
timestamp 1679235063
transform 1 0 5796 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1679235063
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_79
timestamp 1679235063
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_92
timestamp 1679235063
transform 1 0 9568 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1679235063
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1679235063
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_128
timestamp 1679235063
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1679235063
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_139
timestamp 1679235063
transform 1 0 13892 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1679235063
transform 1 0 14812 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1679235063
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1679235063
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1679235063
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_177
timestamp 1679235063
transform 1 0 17388 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_183
timestamp 1679235063
transform 1 0 17940 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_190
timestamp 1679235063
transform 1 0 18584 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_203
timestamp 1679235063
transform 1 0 19780 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_215
timestamp 1679235063
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1679235063
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_244
timestamp 1679235063
transform 1 0 23552 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1679235063
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_9
timestamp 1679235063
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_13
timestamp 1679235063
transform 1 0 2300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_17
timestamp 1679235063
transform 1 0 2668 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1679235063
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_35
timestamp 1679235063
transform 1 0 4324 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_47
timestamp 1679235063
transform 1 0 5428 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_59
timestamp 1679235063
transform 1 0 6532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1679235063
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_71
timestamp 1679235063
transform 1 0 7636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_93
timestamp 1679235063
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_115
timestamp 1679235063
transform 1 0 11684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_119
timestamp 1679235063
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_131
timestamp 1679235063
transform 1 0 13156 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_135
timestamp 1679235063
transform 1 0 13524 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_153
timestamp 1679235063
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_160
timestamp 1679235063
transform 1 0 15824 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_166
timestamp 1679235063
transform 1 0 16376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_170
timestamp 1679235063
transform 1 0 16744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp 1679235063
transform 1 0 17020 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_184
timestamp 1679235063
transform 1 0 18032 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_190
timestamp 1679235063
transform 1 0 18584 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1679235063
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_203
timestamp 1679235063
transform 1 0 19780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_224
timestamp 1679235063
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_228
timestamp 1679235063
transform 1 0 22080 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_232
timestamp 1679235063
transform 1 0 22448 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_265
timestamp 1679235063
transform 1 0 25484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1679235063
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_33
timestamp 1679235063
transform 1 0 4140 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1679235063
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1679235063
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_74
timestamp 1679235063
transform 1 0 7912 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_87
timestamp 1679235063
transform 1 0 9108 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_100
timestamp 1679235063
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_124
timestamp 1679235063
transform 1 0 12512 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_132
timestamp 1679235063
transform 1 0 13248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_144
timestamp 1679235063
transform 1 0 14352 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_148
timestamp 1679235063
transform 1 0 14720 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_158
timestamp 1679235063
transform 1 0 15640 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1679235063
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_174
timestamp 1679235063
transform 1 0 17112 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_183
timestamp 1679235063
transform 1 0 17940 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_192
timestamp 1679235063
transform 1 0 18768 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_204
timestamp 1679235063
transform 1 0 19872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_208
timestamp 1679235063
transform 1 0 20240 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_211
timestamp 1679235063
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1679235063
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1679235063
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1679235063
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1679235063
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1679235063
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1679235063
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_37
timestamp 1679235063
transform 1 0 4508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_49
timestamp 1679235063
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_61
timestamp 1679235063
transform 1 0 6716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_73
timestamp 1679235063
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1679235063
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1679235063
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_105
timestamp 1679235063
transform 1 0 10764 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_110
timestamp 1679235063
transform 1 0 11224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_121
timestamp 1679235063
transform 1 0 12236 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1679235063
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_129
timestamp 1679235063
transform 1 0 12972 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1679235063
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1679235063
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_163
timestamp 1679235063
transform 1 0 16100 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_169
timestamp 1679235063
transform 1 0 16652 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1679235063
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1679235063
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 1679235063
transform 1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_223
timestamp 1679235063
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_259
timestamp 1679235063
transform 1 0 24932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_265
timestamp 1679235063
transform 1 0 25484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_9
timestamp 1679235063
transform 1 0 1932 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_13
timestamp 1679235063
transform 1 0 2300 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_25
timestamp 1679235063
transform 1 0 3404 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_37
timestamp 1679235063
transform 1 0 4508 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1679235063
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_61
timestamp 1679235063
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_71
timestamp 1679235063
transform 1 0 7636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_86
timestamp 1679235063
transform 1 0 9016 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_90
timestamp 1679235063
transform 1 0 9384 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_96
timestamp 1679235063
transform 1 0 9936 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_99
timestamp 1679235063
transform 1 0 10212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_116
timestamp 1679235063
transform 1 0 11776 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_127
timestamp 1679235063
transform 1 0 12788 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_133
timestamp 1679235063
transform 1 0 13340 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_142
timestamp 1679235063
transform 1 0 14168 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_157
timestamp 1679235063
transform 1 0 15548 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1679235063
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_177
timestamp 1679235063
transform 1 0 17388 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_180
timestamp 1679235063
transform 1 0 17664 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1679235063
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_206
timestamp 1679235063
transform 1 0 20056 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_210
timestamp 1679235063
transform 1 0 20424 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1679235063
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_248
timestamp 1679235063
transform 1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_254
timestamp 1679235063
transform 1 0 24472 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1679235063
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_263
timestamp 1679235063
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_9
timestamp 1679235063
transform 1 0 1932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_13
timestamp 1679235063
transform 1 0 2300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_17
timestamp 1679235063
transform 1 0 2668 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1679235063
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_35
timestamp 1679235063
transform 1 0 4324 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_47
timestamp 1679235063
transform 1 0 5428 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_71
timestamp 1679235063
transform 1 0 7636 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_75
timestamp 1679235063
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1679235063
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_93
timestamp 1679235063
transform 1 0 9660 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_107
timestamp 1679235063
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_120
timestamp 1679235063
transform 1 0 12144 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_127
timestamp 1679235063
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_163
timestamp 1679235063
transform 1 0 16100 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_187
timestamp 1679235063
transform 1 0 18308 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_191
timestamp 1679235063
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1679235063
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_219
timestamp 1679235063
transform 1 0 21252 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_223
timestamp 1679235063
transform 1 0 21620 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_230
timestamp 1679235063
transform 1 0 22264 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_21
timestamp 1679235063
transform 1 0 3036 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_33
timestamp 1679235063
transform 1 0 4140 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1679235063
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_59
timestamp 1679235063
transform 1 0 6532 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_91
timestamp 1679235063
transform 1 0 9476 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_98
timestamp 1679235063
transform 1 0 10120 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_102
timestamp 1679235063
transform 1 0 10488 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1679235063
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_115
timestamp 1679235063
transform 1 0 11684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1679235063
transform 1 0 11960 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_126
timestamp 1679235063
transform 1 0 12696 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_140
timestamp 1679235063
transform 1 0 13984 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_152
timestamp 1679235063
transform 1 0 15088 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1679235063
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_176
timestamp 1679235063
transform 1 0 17296 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1679235063
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_215
timestamp 1679235063
transform 1 0 20884 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_219
timestamp 1679235063
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_257
timestamp 1679235063
transform 1 0 24748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1679235063
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1679235063
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_13
timestamp 1679235063
transform 1 0 2300 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_18
timestamp 1679235063
transform 1 0 2760 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1679235063
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_51
timestamp 1679235063
transform 1 0 5796 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_58
timestamp 1679235063
transform 1 0 6440 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_62
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_74
timestamp 1679235063
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 1679235063
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_99
timestamp 1679235063
transform 1 0 10212 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_103
timestamp 1679235063
transform 1 0 10580 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_114
timestamp 1679235063
transform 1 0 11592 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_127
timestamp 1679235063
transform 1 0 12788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_134
timestamp 1679235063
transform 1 0 13432 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_146
timestamp 1679235063
transform 1 0 14536 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_158
timestamp 1679235063
transform 1 0 15640 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_175
timestamp 1679235063
transform 1 0 17204 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_182
timestamp 1679235063
transform 1 0 17848 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_188
timestamp 1679235063
transform 1 0 18400 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_201
timestamp 1679235063
transform 1 0 19596 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_222
timestamp 1679235063
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_230
timestamp 1679235063
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_264
timestamp 1679235063
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1679235063
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1679235063
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_27
timestamp 1679235063
transform 1 0 3588 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_48
timestamp 1679235063
transform 1 0 5520 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1679235063
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_57
timestamp 1679235063
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_65
timestamp 1679235063
transform 1 0 7084 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1679235063
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_80
timestamp 1679235063
transform 1 0 8464 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_93
timestamp 1679235063
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_100
timestamp 1679235063
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1679235063
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_124
timestamp 1679235063
transform 1 0 12512 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_132
timestamp 1679235063
transform 1 0 13248 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_143
timestamp 1679235063
transform 1 0 14260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_147
timestamp 1679235063
transform 1 0 14628 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1679235063
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1679235063
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1679235063
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_193
timestamp 1679235063
transform 1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_201
timestamp 1679235063
transform 1 0 19596 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_206
timestamp 1679235063
transform 1 0 20056 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1679235063
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1679235063
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1679235063
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_257
timestamp 1679235063
transform 1 0 24748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1679235063
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1679235063
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1679235063
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1679235063
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1679235063
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_34
timestamp 1679235063
transform 1 0 4232 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_46
timestamp 1679235063
transform 1 0 5336 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_58
timestamp 1679235063
transform 1 0 6440 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1679235063
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_87
timestamp 1679235063
transform 1 0 9108 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_93
timestamp 1679235063
transform 1 0 9660 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_106
timestamp 1679235063
transform 1 0 10856 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_110
timestamp 1679235063
transform 1 0 11224 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_121
timestamp 1679235063
transform 1 0 12236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1679235063
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1679235063
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_147
timestamp 1679235063
transform 1 0 14628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_157
timestamp 1679235063
transform 1 0 15548 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_181
timestamp 1679235063
transform 1 0 17756 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_187
timestamp 1679235063
transform 1 0 18308 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1679235063
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1679235063
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_208
timestamp 1679235063
transform 1 0 20240 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_220
timestamp 1679235063
transform 1 0 21344 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_237
timestamp 1679235063
transform 1 0 22908 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_243
timestamp 1679235063
transform 1 0 23460 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1679235063
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1679235063
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_259
timestamp 1679235063
transform 1 0 24932 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_263
timestamp 1679235063
transform 1 0 25300 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1679235063
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_14
timestamp 1679235063
transform 1 0 2392 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_20
timestamp 1679235063
transform 1 0 2944 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_29
timestamp 1679235063
transform 1 0 3772 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1679235063
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1679235063
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1679235063
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1679235063
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_69
timestamp 1679235063
transform 1 0 7452 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_78
timestamp 1679235063
transform 1 0 8280 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_82
timestamp 1679235063
transform 1 0 8648 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_86
timestamp 1679235063
transform 1 0 9016 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_97
timestamp 1679235063
transform 1 0 10028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1679235063
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1679235063
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_117
timestamp 1679235063
transform 1 0 11868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_121
timestamp 1679235063
transform 1 0 12236 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_125
timestamp 1679235063
transform 1 0 12604 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_146
timestamp 1679235063
transform 1 0 14536 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_150
timestamp 1679235063
transform 1 0 14904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_154
timestamp 1679235063
transform 1 0 15272 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1679235063
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1679235063
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_177
timestamp 1679235063
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_200
timestamp 1679235063
transform 1 0 19504 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_213
timestamp 1679235063
transform 1 0 20700 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_217
timestamp 1679235063
transform 1 0 21068 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1679235063
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1679235063
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_236
timestamp 1679235063
transform 1 0 22816 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_244
timestamp 1679235063
transform 1 0 23552 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_264
timestamp 1679235063
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1679235063
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1679235063
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1679235063
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1679235063
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_33
timestamp 1679235063
transform 1 0 4140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_45
timestamp 1679235063
transform 1 0 5244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_57
timestamp 1679235063
transform 1 0 6348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_78
timestamp 1679235063
transform 1 0 8280 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1679235063
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1679235063
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_90
timestamp 1679235063
transform 1 0 9384 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_116
timestamp 1679235063
transform 1 0 11776 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_129
timestamp 1679235063
transform 1 0 12972 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1679235063
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_141
timestamp 1679235063
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_146
timestamp 1679235063
transform 1 0 14536 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_154
timestamp 1679235063
transform 1 0 15272 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_175
timestamp 1679235063
transform 1 0 17204 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_181
timestamp 1679235063
transform 1 0 17756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1679235063
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1679235063
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_208
timestamp 1679235063
transform 1 0 20240 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_232
timestamp 1679235063
transform 1 0 22448 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_245
timestamp 1679235063
transform 1 0 23644 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1679235063
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1679235063
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_259
timestamp 1679235063
transform 1 0 24932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_263
timestamp 1679235063
transform 1 0 25300 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1679235063
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_15
timestamp 1679235063
transform 1 0 2484 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_24
timestamp 1679235063
transform 1 0 3312 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_41
timestamp 1679235063
transform 1 0 4876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1679235063
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1679235063
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_79
timestamp 1679235063
transform 1 0 8372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_92
timestamp 1679235063
transform 1 0 9568 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_100
timestamp 1679235063
transform 1 0 10304 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1679235063
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1679235063
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1679235063
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_118
timestamp 1679235063
transform 1 0 11960 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_144
timestamp 1679235063
transform 1 0 14352 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_157
timestamp 1679235063
transform 1 0 15548 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1679235063
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1679235063
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_177
timestamp 1679235063
transform 1 0 17388 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_188
timestamp 1679235063
transform 1 0 18400 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_209
timestamp 1679235063
transform 1 0 20332 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_216
timestamp 1679235063
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1679235063
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_232
timestamp 1679235063
transform 1 0 22448 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_256
timestamp 1679235063
transform 1 0 24656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_264
timestamp 1679235063
transform 1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1679235063
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1679235063
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1679235063
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1679235063
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1679235063
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_53
timestamp 1679235063
transform 1 0 5980 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_75
timestamp 1679235063
transform 1 0 8004 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1679235063
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1679235063
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1679235063
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_129
timestamp 1679235063
transform 1 0 12972 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1679235063
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1679235063
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 1679235063
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_149
timestamp 1679235063
transform 1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_161
timestamp 1679235063
transform 1 0 15916 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_167
timestamp 1679235063
transform 1 0 16468 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_179
timestamp 1679235063
transform 1 0 17572 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_188
timestamp 1679235063
transform 1 0 18400 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1679235063
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1679235063
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_201
timestamp 1679235063
transform 1 0 19596 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_204
timestamp 1679235063
transform 1 0 19872 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_215
timestamp 1679235063
transform 1 0 20884 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_223
timestamp 1679235063
transform 1 0 21620 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_247
timestamp 1679235063
transform 1 0 23828 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1679235063
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_259
timestamp 1679235063
transform 1 0 24932 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_263
timestamp 1679235063
transform 1 0 25300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 1679235063
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_9
timestamp 1679235063
transform 1 0 1932 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_13
timestamp 1679235063
transform 1 0 2300 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_25
timestamp 1679235063
transform 1 0 3404 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_30
timestamp 1679235063
transform 1 0 3864 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_42
timestamp 1679235063
transform 1 0 4968 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1679235063
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1679235063
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_69
timestamp 1679235063
transform 1 0 7452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_77
timestamp 1679235063
transform 1 0 8188 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_98
timestamp 1679235063
transform 1 0 10120 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_102
timestamp 1679235063
transform 1 0 10488 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1679235063
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1679235063
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_128
timestamp 1679235063
transform 1 0 12880 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_134
timestamp 1679235063
transform 1 0 13432 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_146
timestamp 1679235063
transform 1 0 14536 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_47_154
timestamp 1679235063
transform 1 0 15272 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1679235063
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_175
timestamp 1679235063
transform 1 0 17204 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_180
timestamp 1679235063
transform 1 0 17664 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_191
timestamp 1679235063
transform 1 0 18676 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_204
timestamp 1679235063
transform 1 0 19872 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_208
timestamp 1679235063
transform 1 0 20240 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1679235063
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1679235063
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_248
timestamp 1679235063
transform 1 0 23920 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_252
timestamp 1679235063
transform 1 0 24288 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_259
timestamp 1679235063
transform 1 0 24932 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_265
timestamp 1679235063
transform 1 0 25484 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1679235063
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1679235063
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1679235063
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_29
timestamp 1679235063
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_33
timestamp 1679235063
transform 1 0 4140 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_47
timestamp 1679235063
transform 1 0 5428 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_79
timestamp 1679235063
transform 1 0 8372 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1679235063
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1679235063
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_97
timestamp 1679235063
transform 1 0 10028 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_123
timestamp 1679235063
transform 1 0 12420 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_136
timestamp 1679235063
transform 1 0 13616 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1679235063
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_152
timestamp 1679235063
transform 1 0 15088 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_156
timestamp 1679235063
transform 1 0 15456 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_167
timestamp 1679235063
transform 1 0 16468 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_171
timestamp 1679235063
transform 1 0 16836 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_184
timestamp 1679235063
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1679235063
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_219
timestamp 1679235063
transform 1 0 21252 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_223
timestamp 1679235063
transform 1 0 21620 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_235
timestamp 1679235063
transform 1 0 22724 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1679235063
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1679235063
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_258
timestamp 1679235063
transform 1 0 24840 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1679235063
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1679235063
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1679235063
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1679235063
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1679235063
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1679235063
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1679235063
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_69
timestamp 1679235063
transform 1 0 7452 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_92
timestamp 1679235063
transform 1 0 9568 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_96
timestamp 1679235063
transform 1 0 9936 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1679235063
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1679235063
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_121
timestamp 1679235063
transform 1 0 12236 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_133
timestamp 1679235063
transform 1 0 13340 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1679235063
transform 1 0 14536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_159
timestamp 1679235063
transform 1 0 15732 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_165
timestamp 1679235063
transform 1 0 16284 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1679235063
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_180
timestamp 1679235063
transform 1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_186
timestamp 1679235063
transform 1 0 18216 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_198
timestamp 1679235063
transform 1 0 19320 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_204
timestamp 1679235063
transform 1 0 19872 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_215
timestamp 1679235063
transform 1 0 20884 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_219
timestamp 1679235063
transform 1 0 21252 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1679235063
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_236
timestamp 1679235063
transform 1 0 22816 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_246
timestamp 1679235063
transform 1 0 23736 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_251
timestamp 1679235063
transform 1 0 24196 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_259
timestamp 1679235063
transform 1 0 24932 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1679235063
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1679235063
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1679235063
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_29
timestamp 1679235063
transform 1 0 3772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_33
timestamp 1679235063
transform 1 0 4140 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_47
timestamp 1679235063
transform 1 0 5428 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_59
timestamp 1679235063
transform 1 0 6532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_71
timestamp 1679235063
transform 1 0 7636 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1679235063
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_89
timestamp 1679235063
transform 1 0 9292 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_100
timestamp 1679235063
transform 1 0 10304 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_121
timestamp 1679235063
transform 1 0 12236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_134
timestamp 1679235063
transform 1 0 13432 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1679235063
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1679235063
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_147
timestamp 1679235063
transform 1 0 14628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1679235063
transform 1 0 16560 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_181
timestamp 1679235063
transform 1 0 17756 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1679235063
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_197
timestamp 1679235063
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_210
timestamp 1679235063
transform 1 0 20424 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_214
timestamp 1679235063
transform 1 0 20792 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_218
timestamp 1679235063
transform 1 0 21160 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_231
timestamp 1679235063
transform 1 0 22356 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1679235063
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1679235063
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1679235063
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1679235063
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1679235063
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1679235063
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1679235063
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1679235063
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1679235063
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1679235063
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1679235063
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_81
timestamp 1679235063
transform 1 0 8556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_87
timestamp 1679235063
transform 1 0 9108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_95
timestamp 1679235063
transform 1 0 9844 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_99
timestamp 1679235063
transform 1 0 10212 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1679235063
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1679235063
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_118
timestamp 1679235063
transform 1 0 11960 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1679235063
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_137
timestamp 1679235063
transform 1 0 13708 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1679235063
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1679235063
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_175
timestamp 1679235063
transform 1 0 17204 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_188
timestamp 1679235063
transform 1 0 18400 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_194
timestamp 1679235063
transform 1 0 18952 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_198
timestamp 1679235063
transform 1 0 19320 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_202
timestamp 1679235063
transform 1 0 19688 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1679235063
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1679235063
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1679235063
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_237
timestamp 1679235063
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_241
timestamp 1679235063
transform 1 0 23276 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_262
timestamp 1679235063
transform 1 0 25208 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1679235063
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1679235063
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1679235063
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1679235063
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_44
timestamp 1679235063
transform 1 0 5152 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_56
timestamp 1679235063
transform 1 0 6256 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_68
timestamp 1679235063
transform 1 0 7360 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_52_77
timestamp 1679235063
transform 1 0 8188 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1679235063
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1679235063
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1679235063
transform 1 0 9476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_112
timestamp 1679235063
transform 1 0 11408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_116
timestamp 1679235063
transform 1 0 11776 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_120
timestamp 1679235063
transform 1 0 12144 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_125
timestamp 1679235063
transform 1 0 12604 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_136
timestamp 1679235063
transform 1 0 13616 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1679235063
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_153
timestamp 1679235063
transform 1 0 15180 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_159
timestamp 1679235063
transform 1 0 15732 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_162
timestamp 1679235063
transform 1 0 16008 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_184
timestamp 1679235063
transform 1 0 18032 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_188
timestamp 1679235063
transform 1 0 18400 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1679235063
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_208
timestamp 1679235063
transform 1 0 20240 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_212
timestamp 1679235063
transform 1 0 20608 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_224
timestamp 1679235063
transform 1 0 21712 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_236
timestamp 1679235063
transform 1 0 22816 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_240
timestamp 1679235063
transform 1 0 23184 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_244
timestamp 1679235063
transform 1 0 23552 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1679235063
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_253
timestamp 1679235063
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_259
timestamp 1679235063
transform 1 0 24932 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_264
timestamp 1679235063
transform 1 0 25392 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1679235063
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_21
timestamp 1679235063
transform 1 0 3036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1679235063
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1679235063
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1679235063
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_57
timestamp 1679235063
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_67
timestamp 1679235063
transform 1 0 7268 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_78
timestamp 1679235063
transform 1 0 8280 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_91
timestamp 1679235063
transform 1 0 9476 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_95
timestamp 1679235063
transform 1 0 9844 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1679235063
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1679235063
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1679235063
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_125
timestamp 1679235063
transform 1 0 12604 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_148
timestamp 1679235063
transform 1 0 14720 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_152
timestamp 1679235063
transform 1 0 15088 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1679235063
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_169
timestamp 1679235063
transform 1 0 16652 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_172
timestamp 1679235063
transform 1 0 16928 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_183
timestamp 1679235063
transform 1 0 17940 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1679235063
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_209
timestamp 1679235063
transform 1 0 20332 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_215
timestamp 1679235063
transform 1 0 20884 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1679235063
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_225
timestamp 1679235063
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_249
timestamp 1679235063
transform 1 0 24012 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1679235063
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_260
timestamp 1679235063
transform 1 0 25024 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1679235063
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1679235063
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1679235063
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1679235063
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1679235063
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1679235063
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_53
timestamp 1679235063
transform 1 0 5980 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_75
timestamp 1679235063
transform 1 0 8004 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1679235063
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_85
timestamp 1679235063
transform 1 0 8924 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_88
timestamp 1679235063
transform 1 0 9200 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_110
timestamp 1679235063
transform 1 0 11224 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_114
timestamp 1679235063
transform 1 0 11592 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_126
timestamp 1679235063
transform 1 0 12696 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_134
timestamp 1679235063
transform 1 0 13432 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1679235063
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_152
timestamp 1679235063
transform 1 0 15088 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_164
timestamp 1679235063
transform 1 0 16192 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_175
timestamp 1679235063
transform 1 0 17204 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1679235063
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1679235063
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1679235063
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_208
timestamp 1679235063
transform 1 0 20240 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_221
timestamp 1679235063
transform 1 0 21436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_225
timestamp 1679235063
transform 1 0 21804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_235
timestamp 1679235063
transform 1 0 22724 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_247
timestamp 1679235063
transform 1 0 23828 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1679235063
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1679235063
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_259
timestamp 1679235063
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_264
timestamp 1679235063
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1679235063
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1679235063
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_27
timestamp 1679235063
transform 1 0 3588 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_35
timestamp 1679235063
transform 1 0 4324 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_40
timestamp 1679235063
transform 1 0 4784 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1679235063
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1679235063
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_57
timestamp 1679235063
transform 1 0 6348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_66
timestamp 1679235063
transform 1 0 7176 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_91
timestamp 1679235063
transform 1 0 9476 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_98
timestamp 1679235063
transform 1 0 10120 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_102
timestamp 1679235063
transform 1 0 10488 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1679235063
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_113
timestamp 1679235063
transform 1 0 11500 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_116
timestamp 1679235063
transform 1 0 11776 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_127
timestamp 1679235063
transform 1 0 12788 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_134
timestamp 1679235063
transform 1 0 13432 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1679235063
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1679235063
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_180
timestamp 1679235063
transform 1 0 17664 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_193
timestamp 1679235063
transform 1 0 18860 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_199
timestamp 1679235063
transform 1 0 19412 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_205
timestamp 1679235063
transform 1 0 19964 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_209
timestamp 1679235063
transform 1 0 20332 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1679235063
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_227
timestamp 1679235063
transform 1 0 21988 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_232
timestamp 1679235063
transform 1 0 22448 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_239
timestamp 1679235063
transform 1 0 23092 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_243
timestamp 1679235063
transform 1 0 23460 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_255
timestamp 1679235063
transform 1 0 24564 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_259
timestamp 1679235063
transform 1 0 24932 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_264
timestamp 1679235063
transform 1 0 25392 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1679235063
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_8
timestamp 1679235063
transform 1 0 1840 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_20
timestamp 1679235063
transform 1 0 2944 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1679235063
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_41
timestamp 1679235063
transform 1 0 4876 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_65
timestamp 1679235063
transform 1 0 7084 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_78
timestamp 1679235063
transform 1 0 8280 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_85
timestamp 1679235063
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_89
timestamp 1679235063
transform 1 0 9292 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_99
timestamp 1679235063
transform 1 0 10212 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_107
timestamp 1679235063
transform 1 0 10948 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_118
timestamp 1679235063
transform 1 0 11960 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_122
timestamp 1679235063
transform 1 0 12328 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_134
timestamp 1679235063
transform 1 0 13432 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1679235063
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_152
timestamp 1679235063
transform 1 0 15088 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_158
timestamp 1679235063
transform 1 0 15640 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_161
timestamp 1679235063
transform 1 0 15916 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_172
timestamp 1679235063
transform 1 0 16928 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_178
timestamp 1679235063
transform 1 0 17480 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_184
timestamp 1679235063
transform 1 0 18032 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1679235063
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_201
timestamp 1679235063
transform 1 0 19596 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_212
timestamp 1679235063
transform 1 0 20608 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_225
timestamp 1679235063
transform 1 0 21804 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_232
timestamp 1679235063
transform 1 0 22448 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_238
timestamp 1679235063
transform 1 0 23000 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1679235063
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1679235063
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_259
timestamp 1679235063
transform 1 0 24932 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1679235063
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1679235063
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_13
timestamp 1679235063
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_25
timestamp 1679235063
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_37
timestamp 1679235063
transform 1 0 4508 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_45
timestamp 1679235063
transform 1 0 5244 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1679235063
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1679235063
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_57
timestamp 1679235063
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_67
timestamp 1679235063
transform 1 0 7268 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_79
timestamp 1679235063
transform 1 0 8372 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_91
timestamp 1679235063
transform 1 0 9476 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_97
timestamp 1679235063
transform 1 0 10028 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1679235063
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 1679235063
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_121
timestamp 1679235063
transform 1 0 12236 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_137
timestamp 1679235063
transform 1 0 13708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_161
timestamp 1679235063
transform 1 0 15916 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1679235063
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1679235063
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_181
timestamp 1679235063
transform 1 0 17756 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_204
timestamp 1679235063
transform 1 0 19872 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_217
timestamp 1679235063
transform 1 0 21068 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1679235063
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1679235063
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_230
timestamp 1679235063
transform 1 0 22264 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_237
timestamp 1679235063
transform 1 0 22908 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1679235063
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_5
timestamp 1679235063
transform 1 0 1564 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_17
timestamp 1679235063
transform 1 0 2668 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_25
timestamp 1679235063
transform 1 0 3404 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1679235063
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_41
timestamp 1679235063
transform 1 0 4876 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_47
timestamp 1679235063
transform 1 0 5428 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_68
timestamp 1679235063
transform 1 0 7360 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_74
timestamp 1679235063
transform 1 0 7912 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1679235063
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1679235063
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_96
timestamp 1679235063
transform 1 0 9936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_100
timestamp 1679235063
transform 1 0 10304 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_121
timestamp 1679235063
transform 1 0 12236 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_125
timestamp 1679235063
transform 1 0 12604 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1679235063
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_143
timestamp 1679235063
transform 1 0 14260 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_155
timestamp 1679235063
transform 1 0 15364 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_181
timestamp 1679235063
transform 1 0 17756 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_185
timestamp 1679235063
transform 1 0 18124 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_193
timestamp 1679235063
transform 1 0 18860 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1679235063
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_208
timestamp 1679235063
transform 1 0 20240 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_214
timestamp 1679235063
transform 1 0 20792 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_226
timestamp 1679235063
transform 1 0 21896 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_239
timestamp 1679235063
transform 1 0 23092 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_243
timestamp 1679235063
transform 1 0 23460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1679235063
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1679235063
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_258
timestamp 1679235063
transform 1 0 24840 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1679235063
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1679235063
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1679235063
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1679235063
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1679235063
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1679235063
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1679235063
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_80
timestamp 1679235063
transform 1 0 8464 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_104
timestamp 1679235063
transform 1 0 10672 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1679235063
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1679235063
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_135
timestamp 1679235063
transform 1 0 13524 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_139
timestamp 1679235063
transform 1 0 13892 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_151
timestamp 1679235063
transform 1 0 14996 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1679235063
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1679235063
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1679235063
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1679235063
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_205
timestamp 1679235063
transform 1 0 19964 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_210
timestamp 1679235063
transform 1 0 20424 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1679235063
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1679235063
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_236
timestamp 1679235063
transform 1 0 22816 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_249
timestamp 1679235063
transform 1 0 24012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_256
timestamp 1679235063
transform 1 0 24656 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_260
timestamp 1679235063
transform 1 0 25024 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1679235063
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1679235063
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1679235063
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1679235063
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1679235063
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1679235063
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_53
timestamp 1679235063
transform 1 0 5980 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_74
timestamp 1679235063
transform 1 0 7912 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_78
timestamp 1679235063
transform 1 0 8280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_85
timestamp 1679235063
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_98
timestamp 1679235063
transform 1 0 10120 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_110
timestamp 1679235063
transform 1 0 11224 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_122
timestamp 1679235063
transform 1 0 12328 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_128
timestamp 1679235063
transform 1 0 12880 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1679235063
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1679235063
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_153
timestamp 1679235063
transform 1 0 15180 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_175
timestamp 1679235063
transform 1 0 17204 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_179
timestamp 1679235063
transform 1 0 17572 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_191
timestamp 1679235063
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1679235063
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1679235063
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_219
timestamp 1679235063
transform 1 0 21252 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_226
timestamp 1679235063
transform 1 0 21896 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1679235063
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_255
timestamp 1679235063
transform 1 0 24564 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_264
timestamp 1679235063
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1679235063
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_8
timestamp 1679235063
transform 1 0 1840 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_20
timestamp 1679235063
transform 1 0 2944 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_32
timestamp 1679235063
transform 1 0 4048 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1679235063
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_59
timestamp 1679235063
transform 1 0 6532 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_71
timestamp 1679235063
transform 1 0 7636 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_75
timestamp 1679235063
transform 1 0 8004 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_96
timestamp 1679235063
transform 1 0 9936 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_100
timestamp 1679235063
transform 1 0 10304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1679235063
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_135
timestamp 1679235063
transform 1 0 13524 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_141
timestamp 1679235063
transform 1 0 14076 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_148
timestamp 1679235063
transform 1 0 14720 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_160
timestamp 1679235063
transform 1 0 15824 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_169
timestamp 1679235063
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_177
timestamp 1679235063
transform 1 0 17388 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_199
timestamp 1679235063
transform 1 0 19412 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_212
timestamp 1679235063
transform 1 0 20608 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_216
timestamp 1679235063
transform 1 0 20976 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1679235063
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_231
timestamp 1679235063
transform 1 0 22356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_235
timestamp 1679235063
transform 1 0 22724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_260
timestamp 1679235063
transform 1 0 25024 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1679235063
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_13
timestamp 1679235063
transform 1 0 2300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_25
timestamp 1679235063
transform 1 0 3404 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1679235063
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1679235063
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1679235063
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_65
timestamp 1679235063
transform 1 0 7084 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1679235063
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1679235063
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_96
timestamp 1679235063
transform 1 0 9936 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_108
timestamp 1679235063
transform 1 0 11040 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_124
timestamp 1679235063
transform 1 0 12512 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_135
timestamp 1679235063
transform 1 0 13524 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1679235063
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_152
timestamp 1679235063
transform 1 0 15088 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_158
timestamp 1679235063
transform 1 0 15640 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_161
timestamp 1679235063
transform 1 0 15916 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_172
timestamp 1679235063
transform 1 0 16928 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_179
timestamp 1679235063
transform 1 0 17572 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_191
timestamp 1679235063
transform 1 0 18676 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1679235063
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_208
timestamp 1679235063
transform 1 0 20240 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_223
timestamp 1679235063
transform 1 0 21620 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_235
timestamp 1679235063
transform 1 0 22724 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1679235063
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1679235063
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_259
timestamp 1679235063
transform 1 0 24932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1679235063
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_5
timestamp 1679235063
transform 1 0 1564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_17
timestamp 1679235063
transform 1 0 2668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_29
timestamp 1679235063
transform 1 0 3772 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_51
timestamp 1679235063
transform 1 0 5796 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1679235063
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1679235063
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_78
timestamp 1679235063
transform 1 0 8280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_84
timestamp 1679235063
transform 1 0 8832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_95
timestamp 1679235063
transform 1 0 9844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1679235063
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_115
timestamp 1679235063
transform 1 0 11684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_129
timestamp 1679235063
transform 1 0 12972 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_142
timestamp 1679235063
transform 1 0 14168 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_155
timestamp 1679235063
transform 1 0 15364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1679235063
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1679235063
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_171
timestamp 1679235063
transform 1 0 16836 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_182
timestamp 1679235063
transform 1 0 17848 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_194
timestamp 1679235063
transform 1 0 18952 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_199
timestamp 1679235063
transform 1 0 19412 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_214
timestamp 1679235063
transform 1 0 20792 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_218
timestamp 1679235063
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1679235063
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_233
timestamp 1679235063
transform 1 0 22540 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_256
timestamp 1679235063
transform 1 0 24656 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_260
timestamp 1679235063
transform 1 0 25024 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1679235063
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1679235063
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1679235063
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1679235063
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1679235063
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1679235063
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_53
timestamp 1679235063
transform 1 0 5980 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_61
timestamp 1679235063
transform 1 0 6716 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1679235063
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1679235063
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_98
timestamp 1679235063
transform 1 0 10120 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_104
timestamp 1679235063
transform 1 0 10672 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_108
timestamp 1679235063
transform 1 0 11040 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_119
timestamp 1679235063
transform 1 0 12052 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_126
timestamp 1679235063
transform 1 0 12696 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1679235063
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_141
timestamp 1679235063
transform 1 0 14076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_148
timestamp 1679235063
transform 1 0 14720 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_159
timestamp 1679235063
transform 1 0 15732 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_172
timestamp 1679235063
transform 1 0 16928 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_185
timestamp 1679235063
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_192
timestamp 1679235063
transform 1 0 18768 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1679235063
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_210
timestamp 1679235063
transform 1 0 20424 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_214
timestamp 1679235063
transform 1 0 20792 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_219
timestamp 1679235063
transform 1 0 21252 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_232
timestamp 1679235063
transform 1 0 22448 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_244
timestamp 1679235063
transform 1 0 23552 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_253
timestamp 1679235063
transform 1 0 24380 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_258
timestamp 1679235063
transform 1 0 24840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_264
timestamp 1679235063
transform 1 0 25392 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1679235063
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_8
timestamp 1679235063
transform 1 0 1840 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_20
timestamp 1679235063
transform 1 0 2944 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_32
timestamp 1679235063
transform 1 0 4048 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_44
timestamp 1679235063
transform 1 0 5152 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1679235063
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_57
timestamp 1679235063
transform 1 0 6348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_82
timestamp 1679235063
transform 1 0 8648 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_88
timestamp 1679235063
transform 1 0 9200 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_93
timestamp 1679235063
transform 1 0 9660 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_106
timestamp 1679235063
transform 1 0 10856 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1679235063
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_118
timestamp 1679235063
transform 1 0 11960 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_131
timestamp 1679235063
transform 1 0 13156 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_138
timestamp 1679235063
transform 1 0 13800 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_142
timestamp 1679235063
transform 1 0 14168 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_147
timestamp 1679235063
transform 1 0 14628 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_160
timestamp 1679235063
transform 1 0 15824 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_164
timestamp 1679235063
transform 1 0 16192 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1679235063
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_180
timestamp 1679235063
transform 1 0 17664 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_192
timestamp 1679235063
transform 1 0 18768 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_203
timestamp 1679235063
transform 1 0 19780 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_207
timestamp 1679235063
transform 1 0 20148 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_217
timestamp 1679235063
transform 1 0 21068 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1679235063
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1679235063
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_236
timestamp 1679235063
transform 1 0 22816 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_242
timestamp 1679235063
transform 1 0 23368 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1679235063
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1679235063
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_13
timestamp 1679235063
transform 1 0 2300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_25
timestamp 1679235063
transform 1 0 3404 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1679235063
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_41
timestamp 1679235063
transform 1 0 4876 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_67
timestamp 1679235063
transform 1 0 7268 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_71
timestamp 1679235063
transform 1 0 7636 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1679235063
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_85
timestamp 1679235063
transform 1 0 8924 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_97
timestamp 1679235063
transform 1 0 10028 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_110
timestamp 1679235063
transform 1 0 11224 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_116
timestamp 1679235063
transform 1 0 11776 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_126
timestamp 1679235063
transform 1 0 12696 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_130
timestamp 1679235063
transform 1 0 13064 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_133
timestamp 1679235063
transform 1 0 13340 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_137
timestamp 1679235063
transform 1 0 13708 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_141
timestamp 1679235063
transform 1 0 14076 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_152
timestamp 1679235063
transform 1 0 15088 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_160
timestamp 1679235063
transform 1 0 15824 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_181
timestamp 1679235063
transform 1 0 17756 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1679235063
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1679235063
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_208
timestamp 1679235063
transform 1 0 20240 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_221
timestamp 1679235063
transform 1 0 21436 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_225
timestamp 1679235063
transform 1 0 21804 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_236
timestamp 1679235063
transform 1 0 22816 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_249
timestamp 1679235063
transform 1 0 24012 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1679235063
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1679235063
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_5
timestamp 1679235063
transform 1 0 1564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_17
timestamp 1679235063
transform 1 0 2668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_29
timestamp 1679235063
transform 1 0 3772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_41
timestamp 1679235063
transform 1 0 4876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1679235063
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_57
timestamp 1679235063
transform 1 0 6348 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_65
timestamp 1679235063
transform 1 0 7084 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_69
timestamp 1679235063
transform 1 0 7452 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_75
timestamp 1679235063
transform 1 0 8004 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_84
timestamp 1679235063
transform 1 0 8832 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_96
timestamp 1679235063
transform 1 0 9936 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_100
timestamp 1679235063
transform 1 0 10304 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_110
timestamp 1679235063
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_115
timestamp 1679235063
transform 1 0 11684 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_139
timestamp 1679235063
transform 1 0 13892 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_146
timestamp 1679235063
transform 1 0 14536 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_159
timestamp 1679235063
transform 1 0 15732 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_163
timestamp 1679235063
transform 1 0 16100 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1679235063
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1679235063
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_174
timestamp 1679235063
transform 1 0 17112 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_182
timestamp 1679235063
transform 1 0 17848 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_192
timestamp 1679235063
transform 1 0 18768 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_205
timestamp 1679235063
transform 1 0 19964 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_218
timestamp 1679235063
transform 1 0 21160 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_67_225
timestamp 1679235063
transform 1 0 21804 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_248
timestamp 1679235063
transform 1 0 23920 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_252
timestamp 1679235063
transform 1 0 24288 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_257
timestamp 1679235063
transform 1 0 24748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_264
timestamp 1679235063
transform 1 0 25392 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1679235063
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1679235063
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1679235063
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1679235063
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_61
timestamp 1679235063
transform 1 0 6716 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_67
timestamp 1679235063
transform 1 0 7268 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_79
timestamp 1679235063
transform 1 0 8372 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1679235063
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1679235063
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_90
timestamp 1679235063
transform 1 0 9384 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_103
timestamp 1679235063
transform 1 0 10580 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_127
timestamp 1679235063
transform 1 0 12788 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_133
timestamp 1679235063
transform 1 0 13340 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_137
timestamp 1679235063
transform 1 0 13708 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_141
timestamp 1679235063
transform 1 0 14076 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_153
timestamp 1679235063
transform 1 0 15180 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_166
timestamp 1679235063
transform 1 0 16376 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_178
timestamp 1679235063
transform 1 0 17480 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1679235063
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_208
timestamp 1679235063
transform 1 0 20240 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_212
timestamp 1679235063
transform 1 0 20608 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_218
timestamp 1679235063
transform 1 0 21160 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_228
timestamp 1679235063
transform 1 0 22080 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_232
timestamp 1679235063
transform 1 0 22448 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_243
timestamp 1679235063
transform 1 0 23460 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1679235063
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1679235063
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1679235063
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1679235063
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1679235063
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1679235063
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1679235063
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1679235063
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1679235063
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_57
timestamp 1679235063
transform 1 0 6348 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_65
timestamp 1679235063
transform 1 0 7084 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_76
timestamp 1679235063
transform 1 0 8096 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_103
timestamp 1679235063
transform 1 0 10580 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_110
timestamp 1679235063
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_115
timestamp 1679235063
transform 1 0 11684 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_123
timestamp 1679235063
transform 1 0 12420 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_127
timestamp 1679235063
transform 1 0 12788 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_148
timestamp 1679235063
transform 1 0 14720 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_152
timestamp 1679235063
transform 1 0 15088 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_156
timestamp 1679235063
transform 1 0 15456 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_166
timestamp 1679235063
transform 1 0 16376 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_171
timestamp 1679235063
transform 1 0 16836 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_183
timestamp 1679235063
transform 1 0 17940 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_195
timestamp 1679235063
transform 1 0 19044 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_212
timestamp 1679235063
transform 1 0 20608 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_218
timestamp 1679235063
transform 1 0 21160 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_225
timestamp 1679235063
transform 1 0 21804 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_229
timestamp 1679235063
transform 1 0 22172 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_234
timestamp 1679235063
transform 1 0 22632 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_242
timestamp 1679235063
transform 1 0 23368 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1679235063
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1679235063
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_8
timestamp 1679235063
transform 1 0 1840 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_20
timestamp 1679235063
transform 1 0 2944 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1679235063
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1679235063
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_53
timestamp 1679235063
transform 1 0 5980 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_75
timestamp 1679235063
transform 1 0 8004 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_79
timestamp 1679235063
transform 1 0 8372 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_85
timestamp 1679235063
transform 1 0 8924 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_97
timestamp 1679235063
transform 1 0 10028 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_101
timestamp 1679235063
transform 1 0 10396 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_105
timestamp 1679235063
transform 1 0 10764 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_121
timestamp 1679235063
transform 1 0 12236 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_134
timestamp 1679235063
transform 1 0 13432 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_138
timestamp 1679235063
transform 1 0 13800 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_141
timestamp 1679235063
transform 1 0 14076 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_151
timestamp 1679235063
transform 1 0 14996 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_162
timestamp 1679235063
transform 1 0 16008 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_166
timestamp 1679235063
transform 1 0 16376 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_178
timestamp 1679235063
transform 1 0 17480 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_190
timestamp 1679235063
transform 1 0 18584 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_197
timestamp 1679235063
transform 1 0 19228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_205
timestamp 1679235063
transform 1 0 19964 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_210
timestamp 1679235063
transform 1 0 20424 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_214
timestamp 1679235063
transform 1 0 20792 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_224
timestamp 1679235063
transform 1 0 21712 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_230
timestamp 1679235063
transform 1 0 22264 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_241
timestamp 1679235063
transform 1 0 23276 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_247
timestamp 1679235063
transform 1 0 23828 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_259
timestamp 1679235063
transform 1 0 24932 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_264
timestamp 1679235063
transform 1 0 25392 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1679235063
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_13
timestamp 1679235063
transform 1 0 2300 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_21
timestamp 1679235063
transform 1 0 3036 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_26
timestamp 1679235063
transform 1 0 3496 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_30
timestamp 1679235063
transform 1 0 3864 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_42
timestamp 1679235063
transform 1 0 4968 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_54
timestamp 1679235063
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1679235063
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_69
timestamp 1679235063
transform 1 0 7452 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_71_77
timestamp 1679235063
transform 1 0 8188 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_105
timestamp 1679235063
transform 1 0 10764 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_109
timestamp 1679235063
transform 1 0 11132 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_113
timestamp 1679235063
transform 1 0 11500 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_124
timestamp 1679235063
transform 1 0 12512 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_156
timestamp 1679235063
transform 1 0 15456 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_160
timestamp 1679235063
transform 1 0 15824 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_169
timestamp 1679235063
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_191
timestamp 1679235063
transform 1 0 18676 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_197
timestamp 1679235063
transform 1 0 19228 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_208
timestamp 1679235063
transform 1 0 20240 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_212
timestamp 1679235063
transform 1 0 20608 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1679235063
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_225
timestamp 1679235063
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_230
timestamp 1679235063
transform 1 0 22264 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_236
timestamp 1679235063
transform 1 0 22816 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_257
timestamp 1679235063
transform 1 0 24748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1679235063
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_5
timestamp 1679235063
transform 1 0 1564 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_17
timestamp 1679235063
transform 1 0 2668 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_25
timestamp 1679235063
transform 1 0 3404 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1679235063
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_41
timestamp 1679235063
transform 1 0 4876 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_46
timestamp 1679235063
transform 1 0 5336 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_50
timestamp 1679235063
transform 1 0 5704 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_72
timestamp 1679235063
transform 1 0 7728 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_78
timestamp 1679235063
transform 1 0 8280 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_85
timestamp 1679235063
transform 1 0 8924 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_100
timestamp 1679235063
transform 1 0 10304 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_113
timestamp 1679235063
transform 1 0 11500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_117
timestamp 1679235063
transform 1 0 11868 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_129
timestamp 1679235063
transform 1 0 12972 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1679235063
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1679235063
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1679235063
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_153
timestamp 1679235063
transform 1 0 15180 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_161
timestamp 1679235063
transform 1 0 15916 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_173
timestamp 1679235063
transform 1 0 17020 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_177
timestamp 1679235063
transform 1 0 17388 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 1679235063
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_197
timestamp 1679235063
transform 1 0 19228 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_219
timestamp 1679235063
transform 1 0 21252 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_232
timestamp 1679235063
transform 1 0 22448 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_245
timestamp 1679235063
transform 1 0 23644 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_249
timestamp 1679235063
transform 1 0 24012 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_259
timestamp 1679235063
transform 1 0 24932 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1679235063
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1679235063
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1679235063
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_27
timestamp 1679235063
transform 1 0 3588 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_31
timestamp 1679235063
transform 1 0 3956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_37
timestamp 1679235063
transform 1 0 4508 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_45
timestamp 1679235063
transform 1 0 5244 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_49
timestamp 1679235063
transform 1 0 5612 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1679235063
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_57
timestamp 1679235063
transform 1 0 6348 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_63
timestamp 1679235063
transform 1 0 6900 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_67
timestamp 1679235063
transform 1 0 7268 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_89
timestamp 1679235063
transform 1 0 9292 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_102
timestamp 1679235063
transform 1 0 10488 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_106
timestamp 1679235063
transform 1 0 10856 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_73_113
timestamp 1679235063
transform 1 0 11500 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_125
timestamp 1679235063
transform 1 0 12604 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_138
timestamp 1679235063
transform 1 0 13800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_145
timestamp 1679235063
transform 1 0 14444 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_153
timestamp 1679235063
transform 1 0 15180 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_164
timestamp 1679235063
transform 1 0 16192 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_169
timestamp 1679235063
transform 1 0 16652 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_180
timestamp 1679235063
transform 1 0 17664 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_186
timestamp 1679235063
transform 1 0 18216 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_191
timestamp 1679235063
transform 1 0 18676 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_204
timestamp 1679235063
transform 1 0 19872 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_217
timestamp 1679235063
transform 1 0 21068 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_221
timestamp 1679235063
transform 1 0 21436 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1679235063
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_238
timestamp 1679235063
transform 1 0 23000 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_242
timestamp 1679235063
transform 1 0 23368 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_263
timestamp 1679235063
transform 1 0 25300 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1679235063
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_9
timestamp 1679235063
transform 1 0 1932 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_21
timestamp 1679235063
transform 1 0 3036 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1679235063
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_29
timestamp 1679235063
transform 1 0 3772 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_37
timestamp 1679235063
transform 1 0 4508 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_43
timestamp 1679235063
transform 1 0 5060 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_47
timestamp 1679235063
transform 1 0 5428 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_59
timestamp 1679235063
transform 1 0 6532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_71
timestamp 1679235063
transform 1 0 7636 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_79
timestamp 1679235063
transform 1 0 8372 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1679235063
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_93
timestamp 1679235063
transform 1 0 9660 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_101
timestamp 1679235063
transform 1 0 10396 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_125
timestamp 1679235063
transform 1 0 12604 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_129
timestamp 1679235063
transform 1 0 12972 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_137
timestamp 1679235063
transform 1 0 13708 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_141
timestamp 1679235063
transform 1 0 14076 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_145
timestamp 1679235063
transform 1 0 14444 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_169
timestamp 1679235063
transform 1 0 16652 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_173
timestamp 1679235063
transform 1 0 17020 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_183
timestamp 1679235063
transform 1 0 17940 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1679235063
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1679235063
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_197
timestamp 1679235063
transform 1 0 19228 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_220
timestamp 1679235063
transform 1 0 21344 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_224
timestamp 1679235063
transform 1 0 21712 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_234
timestamp 1679235063
transform 1 0 22632 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1679235063
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_255
timestamp 1679235063
transform 1 0 24564 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_265
timestamp 1679235063
transform 1 0 25484 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1679235063
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_13
timestamp 1679235063
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_25
timestamp 1679235063
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_37
timestamp 1679235063
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1679235063
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1679235063
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1679235063
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_69
timestamp 1679235063
transform 1 0 7452 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_75
timestamp 1679235063
transform 1 0 8004 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_83
timestamp 1679235063
transform 1 0 8740 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_96
timestamp 1679235063
transform 1 0 9936 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_100
timestamp 1679235063
transform 1 0 10304 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_105
timestamp 1679235063
transform 1 0 10764 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_110
timestamp 1679235063
transform 1 0 11224 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_113
timestamp 1679235063
transform 1 0 11500 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_121
timestamp 1679235063
transform 1 0 12236 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_143
timestamp 1679235063
transform 1 0 14260 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_156
timestamp 1679235063
transform 1 0 15456 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_160
timestamp 1679235063
transform 1 0 15824 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_171
timestamp 1679235063
transform 1 0 16836 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_182
timestamp 1679235063
transform 1 0 17848 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_186
timestamp 1679235063
transform 1 0 18216 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_207
timestamp 1679235063
transform 1 0 20148 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_211
timestamp 1679235063
transform 1 0 20516 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_219
timestamp 1679235063
transform 1 0 21252 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_225
timestamp 1679235063
transform 1 0 21804 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_236
timestamp 1679235063
transform 1 0 22816 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1679235063
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_5
timestamp 1679235063
transform 1 0 1564 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_17
timestamp 1679235063
transform 1 0 2668 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_25
timestamp 1679235063
transform 1 0 3404 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1679235063
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1679235063
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_53
timestamp 1679235063
transform 1 0 5980 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_59
timestamp 1679235063
transform 1 0 6532 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_64
timestamp 1679235063
transform 1 0 6992 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_68
timestamp 1679235063
transform 1 0 7360 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_76
timestamp 1679235063
transform 1 0 8096 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_82
timestamp 1679235063
transform 1 0 8648 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_85
timestamp 1679235063
transform 1 0 8924 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_108
timestamp 1679235063
transform 1 0 11040 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_116
timestamp 1679235063
transform 1 0 11776 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_120
timestamp 1679235063
transform 1 0 12144 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_132
timestamp 1679235063
transform 1 0 13248 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1679235063
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1679235063
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1679235063
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_177
timestamp 1679235063
transform 1 0 17388 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_181
timestamp 1679235063
transform 1 0 17756 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_184
timestamp 1679235063
transform 1 0 18032 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1679235063
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1679235063
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_221
timestamp 1679235063
transform 1 0 21436 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_76_236
timestamp 1679235063
transform 1 0 22816 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_240
timestamp 1679235063
transform 1 0 23184 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_248
timestamp 1679235063
transform 1 0 23920 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_253
timestamp 1679235063
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_261
timestamp 1679235063
transform 1 0 25116 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1679235063
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1679235063
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1679235063
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1679235063
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_54
timestamp 1679235063
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_57
timestamp 1679235063
transform 1 0 6348 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_63
timestamp 1679235063
transform 1 0 6900 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_71
timestamp 1679235063
transform 1 0 7636 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_78
timestamp 1679235063
transform 1 0 8280 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_88
timestamp 1679235063
transform 1 0 9200 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_92
timestamp 1679235063
transform 1 0 9568 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_104
timestamp 1679235063
transform 1 0 10672 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_110
timestamp 1679235063
transform 1 0 11224 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_115
timestamp 1679235063
transform 1 0 11684 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_126
timestamp 1679235063
transform 1 0 12696 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_130
timestamp 1679235063
transform 1 0 13064 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_151
timestamp 1679235063
transform 1 0 14996 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_157
timestamp 1679235063
transform 1 0 15548 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_165
timestamp 1679235063
transform 1 0 16284 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_169
timestamp 1679235063
transform 1 0 16652 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_191
timestamp 1679235063
transform 1 0 18676 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_195
timestamp 1679235063
transform 1 0 19044 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_199
timestamp 1679235063
transform 1 0 19412 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_220
timestamp 1679235063
transform 1 0 21344 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_225
timestamp 1679235063
transform 1 0 21804 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_229
timestamp 1679235063
transform 1 0 22172 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_250
timestamp 1679235063
transform 1 0 24104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1679235063
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1679235063
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1679235063
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1679235063
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1679235063
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1679235063
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_53
timestamp 1679235063
transform 1 0 5980 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_59
timestamp 1679235063
transform 1 0 6532 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_67
timestamp 1679235063
transform 1 0 7268 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_75
timestamp 1679235063
transform 1 0 8004 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_79
timestamp 1679235063
transform 1 0 8372 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1679235063
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1679235063
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_91
timestamp 1679235063
transform 1 0 9476 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_95
timestamp 1679235063
transform 1 0 9844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_107
timestamp 1679235063
transform 1 0 10948 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_110
timestamp 1679235063
transform 1 0 11224 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_116
timestamp 1679235063
transform 1 0 11776 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_120
timestamp 1679235063
transform 1 0 12144 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_125
timestamp 1679235063
transform 1 0 12604 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_138
timestamp 1679235063
transform 1 0 13800 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_141
timestamp 1679235063
transform 1 0 14076 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_149
timestamp 1679235063
transform 1 0 14812 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_172
timestamp 1679235063
transform 1 0 16928 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_176
timestamp 1679235063
transform 1 0 17296 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_188
timestamp 1679235063
transform 1 0 18400 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_197
timestamp 1679235063
transform 1 0 19228 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_220
timestamp 1679235063
transform 1 0 21344 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_224
timestamp 1679235063
transform 1 0 21712 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_250
timestamp 1679235063
transform 1 0 24104 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_255
timestamp 1679235063
transform 1 0 24564 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_263
timestamp 1679235063
transform 1 0 25300 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_5
timestamp 1679235063
transform 1 0 1564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_17
timestamp 1679235063
transform 1 0 2668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_29
timestamp 1679235063
transform 1 0 3772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_41
timestamp 1679235063
transform 1 0 4876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_53
timestamp 1679235063
transform 1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1679235063
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1679235063
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_81
timestamp 1679235063
transform 1 0 8556 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_86
timestamp 1679235063
transform 1 0 9016 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_108
timestamp 1679235063
transform 1 0 11040 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_115
timestamp 1679235063
transform 1 0 11684 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_121
timestamp 1679235063
transform 1 0 12236 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_133
timestamp 1679235063
transform 1 0 13340 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_141
timestamp 1679235063
transform 1 0 14076 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_164
timestamp 1679235063
transform 1 0 16192 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1679235063
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_181
timestamp 1679235063
transform 1 0 17756 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_187
timestamp 1679235063
transform 1 0 18308 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_208
timestamp 1679235063
transform 1 0 20240 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_212
timestamp 1679235063
transform 1 0 20608 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_225
timestamp 1679235063
transform 1 0 21804 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_247
timestamp 1679235063
transform 1 0 23828 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_251
timestamp 1679235063
transform 1 0 24196 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_264
timestamp 1679235063
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1679235063
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1679235063
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1679235063
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1679235063
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1679235063
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1679235063
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_65
timestamp 1679235063
transform 1 0 7084 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_73
timestamp 1679235063
transform 1 0 7820 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_78
timestamp 1679235063
transform 1 0 8280 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1679235063
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_85
timestamp 1679235063
transform 1 0 8924 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_90
timestamp 1679235063
transform 1 0 9384 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_96
timestamp 1679235063
transform 1 0 9936 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_100
timestamp 1679235063
transform 1 0 10304 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_113
timestamp 1679235063
transform 1 0 11500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_138
timestamp 1679235063
transform 1 0 13800 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_143
timestamp 1679235063
transform 1 0 14260 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_155
timestamp 1679235063
transform 1 0 15364 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_163
timestamp 1679235063
transform 1 0 16100 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_168
timestamp 1679235063
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_180
timestamp 1679235063
transform 1 0 17664 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_188
timestamp 1679235063
transform 1 0 18400 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_193
timestamp 1679235063
transform 1 0 18860 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_197
timestamp 1679235063
transform 1 0 19228 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_200
timestamp 1679235063
transform 1 0 19504 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_211
timestamp 1679235063
transform 1 0 20516 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_224
timestamp 1679235063
transform 1 0 21712 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_228
timestamp 1679235063
transform 1 0 22080 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_250
timestamp 1679235063
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_255
timestamp 1679235063
transform 1 0 24564 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_263
timestamp 1679235063
transform 1 0 25300 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1679235063
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1679235063
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1679235063
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1679235063
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1679235063
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1679235063
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_57
timestamp 1679235063
transform 1 0 6348 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_65
timestamp 1679235063
transform 1 0 7084 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1679235063
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1679235063
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1679235063
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_105
timestamp 1679235063
transform 1 0 10764 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_109
timestamp 1679235063
transform 1 0 11132 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_113
timestamp 1679235063
transform 1 0 11500 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_121
timestamp 1679235063
transform 1 0 12236 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_142
timestamp 1679235063
transform 1 0 14168 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1679235063
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1679235063
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_191
timestamp 1679235063
transform 1 0 18676 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_215
timestamp 1679235063
transform 1 0 20884 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_219
timestamp 1679235063
transform 1 0 21252 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1679235063
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_225
timestamp 1679235063
transform 1 0 21804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_229
timestamp 1679235063
transform 1 0 22172 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_239
timestamp 1679235063
transform 1 0 23092 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_245
timestamp 1679235063
transform 1 0 23644 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_253
timestamp 1679235063
transform 1 0 24380 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1679235063
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1679235063
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1679235063
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1679235063
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1679235063
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1679235063
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1679235063
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1679235063
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1679235063
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1679235063
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_85
timestamp 1679235063
transform 1 0 8924 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_93
timestamp 1679235063
transform 1 0 9660 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_97
timestamp 1679235063
transform 1 0 10028 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_119
timestamp 1679235063
transform 1 0 12052 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_123
timestamp 1679235063
transform 1 0 12420 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1679235063
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1679235063
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_141
timestamp 1679235063
transform 1 0 14076 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_144
timestamp 1679235063
transform 1 0 14352 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_156
timestamp 1679235063
transform 1 0 15456 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_178
timestamp 1679235063
transform 1 0 17480 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_182
timestamp 1679235063
transform 1 0 17848 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1679235063
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_199
timestamp 1679235063
transform 1 0 19412 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_211
timestamp 1679235063
transform 1 0 20516 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_225
timestamp 1679235063
transform 1 0 21804 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_236
timestamp 1679235063
transform 1 0 22816 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_248
timestamp 1679235063
transform 1 0 23920 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_253
timestamp 1679235063
transform 1 0 24380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_259
timestamp 1679235063
transform 1 0 24932 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_264
timestamp 1679235063
transform 1 0 25392 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1679235063
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1679235063
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1679235063
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1679235063
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1679235063
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1679235063
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1679235063
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1679235063
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_81
timestamp 1679235063
transform 1 0 8556 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_90
timestamp 1679235063
transform 1 0 9384 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_102
timestamp 1679235063
transform 1 0 10488 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_110
timestamp 1679235063
transform 1 0 11224 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1679235063
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1679235063
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1679235063
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1679235063
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1679235063
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1679235063
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_169
timestamp 1679235063
transform 1 0 16652 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_180
timestamp 1679235063
transform 1 0 17664 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_193
timestamp 1679235063
transform 1 0 18860 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_197
timestamp 1679235063
transform 1 0 19228 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_209
timestamp 1679235063
transform 1 0 20332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_221
timestamp 1679235063
transform 1 0 21436 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1679235063
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1679235063
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_249
timestamp 1679235063
transform 1 0 24012 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_253
timestamp 1679235063
transform 1 0 24380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1679235063
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1679235063
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_9
timestamp 1679235063
transform 1 0 1932 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_13
timestamp 1679235063
transform 1 0 2300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_25
timestamp 1679235063
transform 1 0 3404 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1679235063
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1679235063
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1679235063
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1679235063
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1679235063
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1679235063
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1679235063
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1679235063
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1679235063
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1679235063
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1679235063
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1679235063
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1679235063
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1679235063
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1679235063
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_177
timestamp 1679235063
transform 1 0 17388 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_182
timestamp 1679235063
transform 1 0 17848 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_194
timestamp 1679235063
transform 1 0 18952 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1679235063
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1679235063
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1679235063
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1679235063
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1679235063
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1679235063
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_253
timestamp 1679235063
transform 1 0 24380 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_259
timestamp 1679235063
transform 1 0 24932 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1679235063
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1679235063
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1679235063
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1679235063
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1679235063
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1679235063
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1679235063
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1679235063
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1679235063
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1679235063
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1679235063
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1679235063
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1679235063
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1679235063
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_125
timestamp 1679235063
transform 1 0 12604 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_129
timestamp 1679235063
transform 1 0 12972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_141
timestamp 1679235063
transform 1 0 14076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_153
timestamp 1679235063
transform 1 0 15180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_165
timestamp 1679235063
transform 1 0 16284 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1679235063
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1679235063
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1679235063
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1679235063
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1679235063
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1679235063
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1679235063
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1679235063
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1679235063
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_261
timestamp 1679235063
transform 1 0 25116 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1679235063
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_21
timestamp 1679235063
transform 1 0 3036 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_86_25
timestamp 1679235063
transform 1 0 3404 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1679235063
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1679235063
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1679235063
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1679235063
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1679235063
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1679235063
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1679235063
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1679235063
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_109
timestamp 1679235063
transform 1 0 11132 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_113
timestamp 1679235063
transform 1 0 11500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_117
timestamp 1679235063
transform 1 0 11868 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_129
timestamp 1679235063
transform 1 0 12972 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_137
timestamp 1679235063
transform 1 0 13708 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1679235063
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1679235063
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1679235063
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1679235063
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1679235063
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1679235063
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1679235063
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1679235063
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1679235063
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1679235063
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1679235063
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1679235063
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_253
timestamp 1679235063
transform 1 0 24380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_259
timestamp 1679235063
transform 1 0 24932 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1679235063
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_87_3
timestamp 1679235063
transform 1 0 1380 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_87_25
timestamp 1679235063
transform 1 0 3404 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_87_54
timestamp 1679235063
transform 1 0 6072 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_61
timestamp 1679235063
transform 1 0 6716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_73
timestamp 1679235063
transform 1 0 7820 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_85
timestamp 1679235063
transform 1 0 8924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_90
timestamp 1679235063
transform 1 0 9384 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_102
timestamp 1679235063
transform 1 0 10488 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_110
timestamp 1679235063
transform 1 0 11224 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1679235063
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1679235063
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1679235063
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1679235063
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1679235063
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1679235063
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1679235063
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1679235063
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1679235063
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1679235063
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1679235063
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1679235063
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1679235063
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1679235063
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1679235063
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1679235063
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_88_3
timestamp 1679235063
transform 1 0 1380 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_9
timestamp 1679235063
transform 1 0 1932 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1679235063
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_29
timestamp 1679235063
transform 1 0 3772 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_41
timestamp 1679235063
transform 1 0 4876 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_45
timestamp 1679235063
transform 1 0 5244 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_57
timestamp 1679235063
transform 1 0 6348 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_61
timestamp 1679235063
transform 1 0 6716 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1679235063
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1679235063
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1679235063
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_88_85
timestamp 1679235063
transform 1 0 8924 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_91
timestamp 1679235063
transform 1 0 9476 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_103
timestamp 1679235063
transform 1 0 10580 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_115
timestamp 1679235063
transform 1 0 11684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_127
timestamp 1679235063
transform 1 0 12788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1679235063
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1679235063
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1679235063
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1679235063
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1679235063
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1679235063
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1679235063
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1679235063
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1679235063
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1679235063
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1679235063
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1679235063
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1679235063
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_253
timestamp 1679235063
transform 1 0 24380 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_261
timestamp 1679235063
transform 1 0 25116 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1679235063
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_8
timestamp 1679235063
transform 1 0 1840 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_12
timestamp 1679235063
transform 1 0 2208 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_29
timestamp 1679235063
transform 1 0 3772 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_49
timestamp 1679235063
transform 1 0 5612 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1679235063
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_57
timestamp 1679235063
transform 1 0 6348 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_65
timestamp 1679235063
transform 1 0 7084 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_79
timestamp 1679235063
transform 1 0 8372 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_87
timestamp 1679235063
transform 1 0 9108 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1679235063
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1679235063
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1679235063
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1679235063
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1679235063
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1679235063
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1679235063
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1679235063
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1679235063
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1679235063
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1679235063
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1679235063
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1679235063
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1679235063
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1679235063
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1679235063
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1679235063
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_249
timestamp 1679235063
transform 1 0 24012 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_255
timestamp 1679235063
transform 1 0 24564 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_258
timestamp 1679235063
transform 1 0 24840 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1679235063
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_3
timestamp 1679235063
transform 1 0 1380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_9
timestamp 1679235063
transform 1 0 1932 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_26
timestamp 1679235063
transform 1 0 3496 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_29
timestamp 1679235063
transform 1 0 3772 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_39
timestamp 1679235063
transform 1 0 4692 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_61
timestamp 1679235063
transform 1 0 6716 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1679235063
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1679235063
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_97
timestamp 1679235063
transform 1 0 10028 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_102
timestamp 1679235063
transform 1 0 10488 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_114
timestamp 1679235063
transform 1 0 11592 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_126
timestamp 1679235063
transform 1 0 12696 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_138
timestamp 1679235063
transform 1 0 13800 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1679235063
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1679235063
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1679235063
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1679235063
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1679235063
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1679235063
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1679235063
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1679235063
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1679235063
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1679235063
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1679235063
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1679235063
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_90_253
timestamp 1679235063
transform 1 0 24380 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_90_258
timestamp 1679235063
transform 1 0 24840 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1679235063
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_91_3
timestamp 1679235063
transform 1 0 1380 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_14
timestamp 1679235063
transform 1 0 2392 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_34
timestamp 1679235063
transform 1 0 4232 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_54
timestamp 1679235063
transform 1 0 6072 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_57
timestamp 1679235063
transform 1 0 6348 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_61
timestamp 1679235063
transform 1 0 6716 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_66
timestamp 1679235063
transform 1 0 7176 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_72
timestamp 1679235063
transform 1 0 7728 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_89
timestamp 1679235063
transform 1 0 9292 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_91_109
timestamp 1679235063
transform 1 0 11132 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_113
timestamp 1679235063
transform 1 0 11500 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_118
timestamp 1679235063
transform 1 0 11960 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1679235063
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_141
timestamp 1679235063
transform 1 0 14076 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_148
timestamp 1679235063
transform 1 0 14720 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_91_152
timestamp 1679235063
transform 1 0 15088 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_160
timestamp 1679235063
transform 1 0 15824 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_164
timestamp 1679235063
transform 1 0 16192 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_91_169
timestamp 1679235063
transform 1 0 16652 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_180
timestamp 1679235063
transform 1 0 17664 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_91_184
timestamp 1679235063
transform 1 0 18032 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_192
timestamp 1679235063
transform 1 0 18768 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_196
timestamp 1679235063
transform 1 0 19136 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_200
timestamp 1679235063
transform 1 0 19504 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_91_206
timestamp 1679235063
transform 1 0 20056 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_212
timestamp 1679235063
transform 1 0 20608 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_216
timestamp 1679235063
transform 1 0 20976 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_220
timestamp 1679235063
transform 1 0 21344 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1679235063
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1679235063
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_237
timestamp 1679235063
transform 1 0 22908 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_242
timestamp 1679235063
transform 1 0 23368 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_246
timestamp 1679235063
transform 1 0 23736 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_251
timestamp 1679235063
transform 1 0 24196 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_255
timestamp 1679235063
transform 1 0 24564 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_258
timestamp 1679235063
transform 1 0 24840 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_264
timestamp 1679235063
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_92_3
timestamp 1679235063
transform 1 0 1380 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_9
timestamp 1679235063
transform 1 0 1932 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_26
timestamp 1679235063
transform 1 0 3496 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_29
timestamp 1679235063
transform 1 0 3772 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_41
timestamp 1679235063
transform 1 0 4876 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_45
timestamp 1679235063
transform 1 0 5244 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_62
timestamp 1679235063
transform 1 0 6808 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1679235063
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1679235063
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_97
timestamp 1679235063
transform 1 0 10028 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_92_121
timestamp 1679235063
transform 1 0 12236 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_128
timestamp 1679235063
transform 1 0 12880 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_132
timestamp 1679235063
transform 1 0 13248 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_92_137
timestamp 1679235063
transform 1 0 13708 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_92_141
timestamp 1679235063
transform 1 0 14076 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_147
timestamp 1679235063
transform 1 0 14628 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_151
timestamp 1679235063
transform 1 0 14996 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_155
timestamp 1679235063
transform 1 0 15364 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_161
timestamp 1679235063
transform 1 0 15916 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_165
timestamp 1679235063
transform 1 0 16284 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_92_168
timestamp 1679235063
transform 1 0 16560 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_175
timestamp 1679235063
transform 1 0 17204 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_183
timestamp 1679235063
transform 1 0 17940 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_191
timestamp 1679235063
transform 1 0 18676 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1679235063
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_197
timestamp 1679235063
transform 1 0 19228 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_203
timestamp 1679235063
transform 1 0 19780 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_211
timestamp 1679235063
transform 1 0 20516 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_219
timestamp 1679235063
transform 1 0 21252 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_227
timestamp 1679235063
transform 1 0 21988 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_234
timestamp 1679235063
transform 1 0 22632 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_92_238
timestamp 1679235063
transform 1 0 23000 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_92_244
timestamp 1679235063
transform 1 0 23552 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_253
timestamp 1679235063
transform 1 0 24380 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_258
timestamp 1679235063
transform 1 0 24840 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1679235063
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_93_3
timestamp 1679235063
transform 1 0 1380 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_14
timestamp 1679235063
transform 1 0 2392 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_34
timestamp 1679235063
transform 1 0 4232 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1679235063
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_57
timestamp 1679235063
transform 1 0 6348 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_67
timestamp 1679235063
transform 1 0 7268 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_73
timestamp 1679235063
transform 1 0 7820 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_90
timestamp 1679235063
transform 1 0 9384 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1679235063
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_115
timestamp 1679235063
transform 1 0 11684 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_133
timestamp 1679235063
transform 1 0 13340 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_145
timestamp 1679235063
transform 1 0 14444 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_157
timestamp 1679235063
transform 1 0 15548 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_93_165
timestamp 1679235063
transform 1 0 16284 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_169
timestamp 1679235063
transform 1 0 16652 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_175
timestamp 1679235063
transform 1 0 17204 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_183
timestamp 1679235063
transform 1 0 17940 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_193
timestamp 1679235063
transform 1 0 18860 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_201
timestamp 1679235063
transform 1 0 19596 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_205
timestamp 1679235063
transform 1 0 19964 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_214
timestamp 1679235063
transform 1 0 20792 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_222
timestamp 1679235063
transform 1 0 21528 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_225
timestamp 1679235063
transform 1 0 21804 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_231
timestamp 1679235063
transform 1 0 22356 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_239
timestamp 1679235063
transform 1 0 23092 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_247
timestamp 1679235063
transform 1 0 23828 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_251
timestamp 1679235063
transform 1 0 24196 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_256
timestamp 1679235063
transform 1 0 24656 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_264
timestamp 1679235063
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1679235063
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_9
timestamp 1679235063
transform 1 0 1932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1679235063
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_29
timestamp 1679235063
transform 1 0 3772 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_39
timestamp 1679235063
transform 1 0 4692 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_45
timestamp 1679235063
transform 1 0 5244 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_62
timestamp 1679235063
transform 1 0 6808 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_82
timestamp 1679235063
transform 1 0 8648 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1679235063
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_97
timestamp 1679235063
transform 1 0 10028 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_117
timestamp 1679235063
transform 1 0 11868 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_94_137
timestamp 1679235063
transform 1 0 13708 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_141
timestamp 1679235063
transform 1 0 14076 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_151
timestamp 1679235063
transform 1 0 14996 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_163
timestamp 1679235063
transform 1 0 16100 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_167
timestamp 1679235063
transform 1 0 16468 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_176
timestamp 1679235063
transform 1 0 17296 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_188
timestamp 1679235063
transform 1 0 18400 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_197
timestamp 1679235063
transform 1 0 19228 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_207
timestamp 1679235063
transform 1 0 20148 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_219
timestamp 1679235063
transform 1 0 21252 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_231
timestamp 1679235063
transform 1 0 22356 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_243
timestamp 1679235063
transform 1 0 23460 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1679235063
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_253
timestamp 1679235063
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_259
timestamp 1679235063
transform 1 0 24932 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_265
timestamp 1679235063
transform 1 0 25484 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1679235063
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1679235063
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1679235063
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_33
timestamp 1679235063
transform 1 0 4140 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1679235063
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1679235063
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1679235063
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1679235063
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1679235063
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_85
timestamp 1679235063
transform 1 0 8924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_93
timestamp 1679235063
transform 1 0 9660 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1679235063
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_113
timestamp 1679235063
transform 1 0 11500 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_118
timestamp 1679235063
transform 1 0 11960 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_138
timestamp 1679235063
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_147
timestamp 1679235063
transform 1 0 14628 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_157
timestamp 1679235063
transform 1 0 15548 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_95_165
timestamp 1679235063
transform 1 0 16284 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1679235063
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_179
timestamp 1679235063
transform 1 0 17572 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_191
timestamp 1679235063
transform 1 0 18676 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_195
timestamp 1679235063
transform 1 0 19044 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1679235063
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_207
timestamp 1679235063
transform 1 0 20148 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_219
timestamp 1679235063
transform 1 0 21252 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1679235063
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1679235063
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_235
timestamp 1679235063
transform 1 0 22724 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_247
timestamp 1679235063
transform 1 0 23828 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_251
timestamp 1679235063
transform 1 0 24196 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_253
timestamp 1679235063
transform 1 0 24380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_259
timestamp 1679235063
transform 1 0 24932 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_263
timestamp 1679235063
transform 1 0 25300 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23276 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 24564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold5
timestamp 1679235063
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  hold6
timestamp 1679235063
transform 1 0 22172 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 22448 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform 1 0 6532 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 3956 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1679235063
transform 1 0 1564 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 3036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 1564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold14
timestamp 1679235063
transform 1 0 2852 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1679235063
transform 1 0 1564 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold16
timestamp 1679235063
transform 1 0 3956 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1679235063
transform 1 0 1564 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold18
timestamp 1679235063
transform 1 0 3128 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1679235063
transform 1 0 1564 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold20
timestamp 1679235063
transform 1 0 2944 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1679235063
transform 1 0 18124 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1679235063
transform 1 0 14812 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform 1 0 20056 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform 1 0 16836 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 1656 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 21620 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 20516 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 13708 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 6532 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1679235063
transform 1 0 19412 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 14812 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 17664 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 15364 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform 1 0 23092 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 3680 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 7912 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform 1 0 14260 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform 1 0 6532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1679235063
transform 1 0 17940 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1679235063
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform 1 0 16560 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1679235063
transform 1 0 19412 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1679235063
transform 1 0 1656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1679235063
transform 1 0 21988 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform 1 0 22724 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1679235063
transform 1 0 2116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1679235063
transform 1 0 20516 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1679235063
transform 1 0 4600 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1679235063
transform 1 0 7912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1679235063
transform 1 0 9844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1679235063
transform 1 0 6808 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1679235063
transform 1 0 6808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 9384 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1679235063
transform 1 0 9200 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1679235063
transform 1 0 11684 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1679235063
transform 1 0 5704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1679235063
transform 1 0 1564 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1679235063
transform 1 0 1748 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1679235063
transform 1 0 3956 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold62
timestamp 1679235063
transform 1 0 1656 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1679235063
transform 1 0 1656 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold65
timestamp 1679235063
transform 1 0 1748 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1679235063
transform 1 0 2484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 1564 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 2392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 25116 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1679235063
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1679235063
transform 1 0 25116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1679235063
transform 1 0 25116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1679235063
transform 1 0 25116 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 25116 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1679235063
transform 1 0 24472 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 25116 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1679235063
transform 1 0 25116 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 25116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1679235063
transform 1 0 23184 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1679235063
transform 1 0 24472 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1679235063
transform 1 0 24472 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1679235063
transform 1 0 24472 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1679235063
transform 1 0 23184 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1679235063
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1679235063
transform 1 0 24472 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1679235063
transform 1 0 25116 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1679235063
transform 1 0 25116 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1679235063
transform 1 0 25116 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1679235063
transform 1 0 23920 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1679235063
transform 1 0 23828 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1679235063
transform 1 0 25116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1679235063
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 25116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1679235063
transform 1 0 25116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1679235063
transform 1 0 25116 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1679235063
transform 1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1679235063
transform 1 0 5704 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1679235063
transform 1 0 6532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1679235063
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1679235063
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1679235063
transform 1 0 7636 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1679235063
transform 1 0 7912 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1679235063
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1679235063
transform 1 0 8280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1679235063
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1679235063
transform 1 0 9016 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1679235063
transform 1 0 8648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1679235063
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1679235063
transform 1 0 9568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1679235063
transform 1 0 10304 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1679235063
transform 1 0 10948 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1679235063
transform 1 0 11684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1679235063
transform 1 0 11684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1679235063
transform 1 0 10304 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1679235063
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1679235063
transform 1 0 2852 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1679235063
transform 1 0 3220 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1679235063
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1679235063
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1679235063
transform 1 0 3956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1679235063
transform 1 0 4692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1679235063
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1679235063
transform 1 0 11684 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1679235063
transform 1 0 16836 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1679235063
transform 1 0 17572 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1679235063
transform 1 0 17388 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1679235063
transform 1 0 19228 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1679235063
transform 1 0 18308 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1679235063
transform 1 0 20148 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1679235063
transform 1 0 18860 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1679235063
transform 1 0 19412 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1679235063
transform 1 0 20884 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1679235063
transform 1 0 21160 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1679235063
transform 1 0 13340 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1679235063
transform 1 0 20332 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1679235063
transform 1 0 21620 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1679235063
transform 1 0 21988 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1679235063
transform 1 0 22724 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1679235063
transform 1 0 22356 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1679235063
transform 1 0 23828 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input81
timestamp 1679235063
transform 1 0 23460 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1679235063
transform 1 0 23092 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1679235063
transform 1 0 23276 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1679235063
transform 1 0 23920 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1679235063
transform 1 0 13708 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1679235063
transform 1 0 14260 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1679235063
transform 1 0 14444 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input88
timestamp 1679235063
transform 1 0 15916 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input89
timestamp 1679235063
transform 1 0 15548 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1679235063
transform 1 0 15916 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1679235063
transform 1 0 15916 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1679235063
transform 1 0 16836 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1679235063
transform 1 0 1564 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1679235063
transform 1 0 1564 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1679235063
transform 1 0 1564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1679235063
transform 1 0 1564 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1679235063
transform 1 0 1564 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1679235063
transform 1 0 25116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1679235063
transform 1 0 25024 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input100
timestamp 1679235063
transform 1 0 25024 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1679235063
transform 1 0 25024 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1679235063
transform 1 0 25024 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1679235063
transform 1 0 25024 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1679235063
transform 1 0 24288 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input105
timestamp 1679235063
transform 1 0 24564 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1679235063
transform 1 0 24564 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input107
timestamp 1679235063
transform 1 0 1564 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1679235063
transform 1 0 1564 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input109
timestamp 1679235063
transform 1 0 3956 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input110
timestamp 1679235063
transform 1 0 3956 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__conb_1  left_tile_210
timestamp 1679235063
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 18216 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 1564 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 22632 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 22080 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 23920 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 22632 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 23920 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 20056 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform 1 0 22080 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform 1 0 23920 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform 1 0 23920 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform 1 0 22632 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform 1 0 22080 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform 1 0 23920 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform 1 0 22632 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 23920 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform 1 0 17572 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform 1 0 23920 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1679235063
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1679235063
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1679235063
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1679235063
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1679235063
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1679235063
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1679235063
transform 1 0 19412 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1679235063
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1679235063
transform 1 0 19412 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1679235063
transform 1 0 21252 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1679235063
transform 1 0 12420 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1679235063
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1679235063
transform 1 0 20516 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1679235063
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1679235063
transform 1 0 17480 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1679235063
transform 1 0 22356 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1679235063
transform 1 0 21988 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1679235063
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1679235063
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1679235063
transform 1 0 20792 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1679235063
transform 1 0 17480 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1679235063
transform 1 0 13524 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1679235063
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1679235063
transform 1 0 14260 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1679235063
transform 1 0 14628 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1679235063
transform 1 0 14996 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1679235063
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1679235063
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1679235063
transform 1 0 16836 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1679235063
transform 1 0 1932 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1679235063
transform 1 0 2024 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1679235063
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1679235063
transform 1 0 4600 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1679235063
transform 1 0 5336 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1679235063
transform 1 0 7084 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1679235063
transform 1 0 5336 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1679235063
transform 1 0 7176 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1679235063
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1679235063
transform 1 0 7820 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1679235063
transform 1 0 7176 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1679235063
transform 1 0 2024 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1679235063
transform 1 0 7912 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1679235063
transform 1 0 9660 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1679235063
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1679235063
transform 1 0 9752 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1679235063
transform 1 0 10764 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1679235063
transform 1 0 10396 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1679235063
transform 1 0 9752 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1679235063
transform 1 0 11868 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1679235063
transform 1 0 12236 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1679235063
transform 1 0 12328 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1679235063
transform 1 0 2300 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1679235063
transform 1 0 2024 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1679235063
transform 1 0 2760 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1679235063
transform 1 0 2024 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1679235063
transform 1 0 4140 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1679235063
transform 1 0 2760 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1679235063
transform 1 0 4600 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1679235063
transform 1 0 5244 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1679235063
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1679235063
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1679235063
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1679235063
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1679235063
transform 1 0 1564 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1679235063
transform 1 0 1564 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1679235063
transform 1 0 1564 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1679235063
transform 1 0 1564 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1679235063
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1679235063
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1679235063
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1679235063
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1679235063
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1679235063
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1679235063
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1679235063
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1679235063
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1679235063
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1679235063
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1679235063
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1679235063
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1679235063
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1679235063
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1679235063
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1679235063
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1679235063
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1679235063
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1679235063
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1679235063
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1679235063
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1679235063
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1679235063
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1679235063
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1679235063
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1679235063
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1679235063
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1679235063
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1679235063
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1679235063
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1679235063
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1679235063
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1679235063
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1679235063
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1679235063
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1679235063
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1679235063
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1679235063
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1679235063
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1679235063
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1679235063
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1679235063
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1679235063
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1679235063
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1679235063
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1679235063
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1679235063
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1679235063
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1679235063
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1679235063
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1679235063
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1679235063
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1679235063
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1679235063
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1679235063
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1679235063
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1679235063
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1679235063
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1679235063
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1679235063
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1679235063
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1679235063
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1679235063
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1679235063
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1679235063
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1679235063
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1679235063
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1679235063
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1679235063
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1679235063
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1679235063
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1679235063
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1679235063
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1679235063
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1679235063
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1679235063
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1679235063
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1679235063
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1679235063
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1679235063
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1679235063
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1679235063
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1679235063
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1679235063
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1679235063
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1679235063
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1679235063
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1679235063
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1679235063
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1679235063
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1679235063
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1679235063
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1679235063
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1679235063
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1679235063
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1679235063
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1679235063
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1679235063
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1679235063
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1679235063
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1679235063
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1679235063
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1679235063
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1679235063
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1679235063
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1679235063
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1679235063
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1679235063
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1679235063
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16192 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16468 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19872 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22908 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18768 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15364 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 15916 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17572 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 20608 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21896 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22816 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 22908 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16192 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 14444 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14076 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 12880 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15916 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 18032 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15364 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9108 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17572 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22172 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23368 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23460 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22908 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23552 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23460 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22080 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 22264 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23092 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22816 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 23552 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23460 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 22264 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19504 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19412 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19504 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19504 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 18308 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18400 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19044 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 16836 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15640 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 15088 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14536 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14352 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 13616 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12880 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12052 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 11684 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10396 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 9568 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10580 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12512 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12696 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11132 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9936 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8280 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7728 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6532 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6164 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6532 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6440 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6808 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7636 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11500 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12788 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14536 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15364 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17664 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18860 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19872 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22080 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21712 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20884 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18216 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 3956 0 -1 50048
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9200 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 10212 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11868 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13156 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 12328 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12328 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10948 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 8924 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8464 0 -1 40256
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6808 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 5428 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6532 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 5520 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 4232 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6532 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6164 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 5244 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7544 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9384 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 8832 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8096 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6072 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 3956 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 4876 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6164 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 5888 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7452 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10764 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14812 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 15916 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18032 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 11960 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15364 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1__260
timestamp 1679235063
transform 1 0 13892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 13524 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 14720 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19044 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1__211
timestamp 1679235063
transform 1 0 17664 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17204 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 18952 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19596 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20056 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21988 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_2_
timestamp 1679235063
transform 1 0 20240 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22816 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1_
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1__214
timestamp 1679235063
transform 1 0 21988 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l3_in_0_
timestamp 1679235063
transform 1 0 22080 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17848 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20608 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_2_
timestamp 1679235063
transform 1 0 18032 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3__216
timestamp 1679235063
transform 1 0 17020 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3_
timestamp 1679235063
transform 1 0 16836 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_1_
timestamp 1679235063
transform 1 0 18032 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19228 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17112 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_2_
timestamp 1679235063
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3_
timestamp 1679235063
transform 1 0 13432 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3__261
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17204 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14720 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16376 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17572 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20700 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_2_
timestamp 1679235063
transform 1 0 17572 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19596 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1__262
timestamp 1679235063
transform 1 0 20700 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1_
timestamp 1679235063
transform 1 0 19504 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19872 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18492 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19504 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_2_
timestamp 1679235063
transform 1 0 20056 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21528 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1__263
timestamp 1679235063
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1_
timestamp 1679235063
transform 1 0 22080 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l3_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23184 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16100 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19964 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_2_
timestamp 1679235063
transform 1 0 18124 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1__264
timestamp 1679235063
transform 1 0 16928 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1_
timestamp 1679235063
transform 1 0 16836 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l3_in_0_
timestamp 1679235063
transform 1 0 15640 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15548 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17940 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19780 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12788 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1__212
timestamp 1679235063
transform 1 0 12604 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l3_in_0_
timestamp 1679235063
transform 1 0 13708 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13064 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20332 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20792 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1_
timestamp 1679235063
transform 1 0 21068 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1__213
timestamp 1679235063
transform 1 0 22632 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18308 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14904 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1__215
timestamp 1679235063
transform 1 0 14352 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14996 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11224 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10396 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20976 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21896 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_0.mux_l2_in_1__217
timestamp 1679235063
transform 1 0 20884 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 22908 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22264 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21252 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 20240 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22816 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_2.mux_l2_in_1__223
timestamp 1679235063
transform 1 0 23828 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 22632 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23184 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_4.mux_l2_in_1__234
timestamp 1679235063
transform 1 0 21988 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 19780 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 22264 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23644 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_2_
timestamp 1679235063
transform 1 0 20240 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_6.mux_l2_in_1__243
timestamp 1679235063
transform 1 0 22448 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 23184 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20884 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_2_
timestamp 1679235063
transform 1 0 18952 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21804 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_1_
timestamp 1679235063
transform 1 0 21620 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_8.mux_l2_in_1__244
timestamp 1679235063
transform 1 0 21988 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l3_in_0_
timestamp 1679235063
transform 1 0 22448 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20884 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19780 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20240 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_10.mux_l2_in_1__218
timestamp 1679235063
transform 1 0 17296 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 16100 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 20608 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 22172 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19688 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_12.mux_l2_in_1__219
timestamp 1679235063
transform 1 0 18492 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_1_
timestamp 1679235063
transform 1 0 17020 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 22816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_14.mux_l2_in_1__220
timestamp 1679235063
transform 1 0 16836 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_1_
timestamp 1679235063
transform 1 0 16836 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l3_in_0_
timestamp 1679235063
transform 1 0 18216 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 22172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18032 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17020 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14352 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_16.mux_l2_in_1__221
timestamp 1679235063
transform 1 0 14260 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16652 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20056 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16192 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_18.mux_l2_in_1__222
timestamp 1679235063
transform 1 0 13524 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12880 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16100 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14628 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13340 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_20.mux_l2_in_1__224
timestamp 1679235063
transform 1 0 13156 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11960 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l3_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12604 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_22.mux_l2_in_1__225
timestamp 1679235063
transform 1 0 11684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_1_
timestamp 1679235063
transform 1 0 10396 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l3_in_0_
timestamp 1679235063
transform 1 0 12604 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17572 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15088 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12604 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_24.mux_l1_in_1__226
timestamp 1679235063
transform 1 0 13156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14812 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_26.mux_l1_in_1__227
timestamp 1679235063
transform 1 0 11960 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_1_
timestamp 1679235063
transform 1 0 11408 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14720 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_1_
timestamp 1679235063
transform 1 0 9200 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_28.mux_l1_in_1__228
timestamp 1679235063
transform 1 0 9384 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12144 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12512 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_1_
timestamp 1679235063
transform 1 0 8740 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_30.mux_l1_in_1__229
timestamp 1679235063
transform 1 0 9108 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16008 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11408 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_32.mux_l1_in_1__230
timestamp 1679235063
transform 1 0 8004 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_1_
timestamp 1679235063
transform 1 0 7636 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10028 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15456 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14904 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_34.mux_l1_in_1__231
timestamp 1679235063
transform 1 0 10028 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_1_
timestamp 1679235063
transform 1 0 8832 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10764 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 7268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_36.mux_l2_in_1__232
timestamp 1679235063
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_1_
timestamp 1679235063
transform 1 0 6532 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l3_in_0_
timestamp 1679235063
transform 1 0 8188 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14628 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12236 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14996 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_38.mux_l2_in_0__233
timestamp 1679235063
transform 1 0 14720 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14168 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_40.mux_l2_in_0__235
timestamp 1679235063
transform 1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16192 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_44.mux_l2_in_0__236
timestamp 1679235063
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18400 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20424 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17480 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20056 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_46.mux_l2_in_0__237
timestamp 1679235063
transform 1 0 20424 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 22632 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_48.mux_l2_in_0__238
timestamp 1679235063
transform 1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23276 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_50.mux_l1_in_1__239
timestamp 1679235063
transform 1 0 20424 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19228 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23000 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_52.mux_l2_in_0__240
timestamp 1679235063
transform 1 0 21988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21068 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 22724 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17756 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_54.mux_l2_in_0__241
timestamp 1679235063
transform 1 0 19596 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19136 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21528 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17296 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_56.mux_l2_in_0__242
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 9108 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 17112 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14904 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 10028 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_0.mux_l1_in_3__245
timestamp 1679235063
transform 1 0 9384 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11868 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11684 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10672 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11592 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 12696 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15364 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_2.mux_l2_in_1__248
timestamp 1679235063
transform 1 0 14168 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 12972 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12696 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15180 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_2_
timestamp 1679235063
transform 1 0 11132 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 10396 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_4.mux_l2_in_1__252
timestamp 1679235063
transform 1 0 11684 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10672 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 9200 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18124 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_2_
timestamp 1679235063
transform 1 0 14260 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_6.mux_l1_in_3__255
timestamp 1679235063
transform 1 0 9844 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_3_
timestamp 1679235063
transform 1 0 8648 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9752 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9292 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 7268 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 9108 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 17296 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_2_
timestamp 1679235063
transform 1 0 12788 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_10.mux_l1_in_3__246
timestamp 1679235063
transform 1 0 7912 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_3_
timestamp 1679235063
transform 1 0 7452 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9200 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9108 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 7452 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8004 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12144 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_1_
timestamp 1679235063
transform 1 0 16376 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_2_
timestamp 1679235063
transform 1 0 7820 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_1_
timestamp 1679235063
transform 1 0 7452 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_12.mux_l2_in_1__247
timestamp 1679235063
transform 1 0 6900 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l3_in_0_
timestamp 1679235063
transform 1 0 7636 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7728 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14536 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_1_
timestamp 1679235063
transform 1 0 18308 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_2_
timestamp 1679235063
transform 1 0 9476 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_20.mux_l2_in_1__249
timestamp 1679235063
transform 1 0 9752 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9384 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9016 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8372 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12328 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12880 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_28.mux_l2_in_1__250
timestamp 1679235063
transform 1 0 5336 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_1_
timestamp 1679235063
transform 1 0 4968 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l3_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5796 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l1_in_0_
timestamp 1679235063
transform -1 0 12236 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11868 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_36.mux_l2_in_1__251
timestamp 1679235063
transform 1 0 9108 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_1_
timestamp 1679235063
transform 1 0 7820 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9660 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7176 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_44.mux_l1_in_1__253
timestamp 1679235063
transform 1 0 10948 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10396 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19136 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_52.mux_l2_in_1__254
timestamp 1679235063
transform 1 0 14444 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l3_in_0_
timestamp 1679235063
transform 1 0 15548 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10028 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1679235063
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1679235063
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1679235063
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1679235063
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1679235063
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1679235063
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1679235063
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1679235063
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1679235063
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1679235063
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1679235063
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1679235063
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1679235063
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1679235063
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1679235063
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1679235063
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1679235063
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1679235063
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1679235063
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1679235063
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1679235063
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1679235063
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1679235063
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1679235063
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1679235063
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1679235063
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1679235063
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1679235063
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1679235063
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1679235063
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1679235063
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1679235063
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1679235063
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1679235063
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1679235063
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1679235063
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1679235063
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1679235063
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1679235063
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1679235063
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1679235063
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1679235063
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1679235063
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1679235063
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1679235063
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1679235063
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1679235063
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1679235063
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1679235063
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1679235063
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1679235063
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1679235063
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1679235063
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1679235063
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1679235063
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1679235063
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1679235063
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1679235063
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1679235063
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1679235063
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1679235063
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1679235063
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1679235063
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1679235063
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1679235063
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1679235063
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1679235063
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1679235063
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1679235063
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1679235063
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1679235063
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1679235063
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1679235063
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1679235063
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1679235063
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1679235063
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1679235063
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1679235063
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1679235063
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1679235063
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1679235063
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1679235063
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1679235063
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1679235063
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1679235063
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1679235063
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1679235063
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1679235063
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1679235063
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1679235063
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1679235063
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1679235063
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1679235063
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1679235063
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1679235063
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1679235063
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1679235063
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1679235063
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1679235063
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1679235063
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1679235063
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1679235063
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1679235063
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1679235063
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1679235063
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1679235063
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1679235063
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1679235063
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1679235063
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1679235063
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1679235063
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1679235063
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1679235063
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1679235063
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1679235063
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1679235063
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1679235063
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1679235063
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1679235063
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1679235063
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1679235063
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1679235063
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1679235063
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1679235063
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1679235063
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1679235063
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1679235063
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1679235063
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1679235063
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1679235063
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1679235063
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1679235063
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1679235063
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1679235063
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1679235063
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1679235063
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1679235063
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1679235063
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1679235063
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1679235063
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1679235063
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1679235063
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1679235063
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1679235063
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1679235063
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1679235063
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1679235063
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1679235063
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1679235063
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1679235063
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1679235063
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1679235063
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1679235063
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1679235063
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1679235063
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1679235063
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1679235063
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1679235063
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1679235063
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1679235063
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1679235063
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1679235063
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1679235063
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1679235063
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 55360 800 55480 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1490 56200 1546 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1674 0 1730 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 66 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 67 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 68 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 69 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 70 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 71 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 72 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 73 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 74 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 75 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 76 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 77 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 chany_bottom_in[20]
port 78 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 chany_bottom_in[21]
port 79 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 chany_bottom_in[22]
port 80 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_in[23]
port 81 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 chany_bottom_in[24]
port 82 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_in[25]
port 83 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 chany_bottom_in[26]
port 84 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 chany_bottom_in[27]
port 85 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 chany_bottom_in[28]
port 86 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 chany_bottom_in[29]
port 87 nsew signal input
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 88 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 89 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 90 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 91 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 92 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 93 nsew signal input
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 94 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 95 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 96 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 97 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 98 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 99 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 100 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 101 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 102 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 103 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 104 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 105 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 106 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 107 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 chany_bottom_out[20]
port 108 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 chany_bottom_out[21]
port 109 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 chany_bottom_out[22]
port 110 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 chany_bottom_out[23]
port 111 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 chany_bottom_out[24]
port 112 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 chany_bottom_out[25]
port 113 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 chany_bottom_out[26]
port 114 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 chany_bottom_out[27]
port 115 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 chany_bottom_out[28]
port 116 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 chany_bottom_out[29]
port 117 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 118 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 119 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 120 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 121 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 122 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 123 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 124 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 125 nsew signal tristate
flabel metal2 s 12898 56200 12954 57000 0 FreeSans 224 90 0 0 chany_top_in_0[0]
port 126 nsew signal input
flabel metal2 s 16578 56200 16634 57000 0 FreeSans 224 90 0 0 chany_top_in_0[10]
port 127 nsew signal input
flabel metal2 s 16946 56200 17002 57000 0 FreeSans 224 90 0 0 chany_top_in_0[11]
port 128 nsew signal input
flabel metal2 s 17314 56200 17370 57000 0 FreeSans 224 90 0 0 chany_top_in_0[12]
port 129 nsew signal input
flabel metal2 s 17682 56200 17738 57000 0 FreeSans 224 90 0 0 chany_top_in_0[13]
port 130 nsew signal input
flabel metal2 s 18050 56200 18106 57000 0 FreeSans 224 90 0 0 chany_top_in_0[14]
port 131 nsew signal input
flabel metal2 s 18418 56200 18474 57000 0 FreeSans 224 90 0 0 chany_top_in_0[15]
port 132 nsew signal input
flabel metal2 s 18786 56200 18842 57000 0 FreeSans 224 90 0 0 chany_top_in_0[16]
port 133 nsew signal input
flabel metal2 s 19154 56200 19210 57000 0 FreeSans 224 90 0 0 chany_top_in_0[17]
port 134 nsew signal input
flabel metal2 s 19522 56200 19578 57000 0 FreeSans 224 90 0 0 chany_top_in_0[18]
port 135 nsew signal input
flabel metal2 s 19890 56200 19946 57000 0 FreeSans 224 90 0 0 chany_top_in_0[19]
port 136 nsew signal input
flabel metal2 s 13266 56200 13322 57000 0 FreeSans 224 90 0 0 chany_top_in_0[1]
port 137 nsew signal input
flabel metal2 s 20258 56200 20314 57000 0 FreeSans 224 90 0 0 chany_top_in_0[20]
port 138 nsew signal input
flabel metal2 s 20626 56200 20682 57000 0 FreeSans 224 90 0 0 chany_top_in_0[21]
port 139 nsew signal input
flabel metal2 s 20994 56200 21050 57000 0 FreeSans 224 90 0 0 chany_top_in_0[22]
port 140 nsew signal input
flabel metal2 s 21362 56200 21418 57000 0 FreeSans 224 90 0 0 chany_top_in_0[23]
port 141 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 chany_top_in_0[24]
port 142 nsew signal input
flabel metal2 s 22098 56200 22154 57000 0 FreeSans 224 90 0 0 chany_top_in_0[25]
port 143 nsew signal input
flabel metal2 s 22466 56200 22522 57000 0 FreeSans 224 90 0 0 chany_top_in_0[26]
port 144 nsew signal input
flabel metal2 s 22834 56200 22890 57000 0 FreeSans 224 90 0 0 chany_top_in_0[27]
port 145 nsew signal input
flabel metal2 s 23202 56200 23258 57000 0 FreeSans 224 90 0 0 chany_top_in_0[28]
port 146 nsew signal input
flabel metal2 s 23570 56200 23626 57000 0 FreeSans 224 90 0 0 chany_top_in_0[29]
port 147 nsew signal input
flabel metal2 s 13634 56200 13690 57000 0 FreeSans 224 90 0 0 chany_top_in_0[2]
port 148 nsew signal input
flabel metal2 s 14002 56200 14058 57000 0 FreeSans 224 90 0 0 chany_top_in_0[3]
port 149 nsew signal input
flabel metal2 s 14370 56200 14426 57000 0 FreeSans 224 90 0 0 chany_top_in_0[4]
port 150 nsew signal input
flabel metal2 s 14738 56200 14794 57000 0 FreeSans 224 90 0 0 chany_top_in_0[5]
port 151 nsew signal input
flabel metal2 s 15106 56200 15162 57000 0 FreeSans 224 90 0 0 chany_top_in_0[6]
port 152 nsew signal input
flabel metal2 s 15474 56200 15530 57000 0 FreeSans 224 90 0 0 chany_top_in_0[7]
port 153 nsew signal input
flabel metal2 s 15842 56200 15898 57000 0 FreeSans 224 90 0 0 chany_top_in_0[8]
port 154 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 chany_top_in_0[9]
port 155 nsew signal input
flabel metal2 s 1858 56200 1914 57000 0 FreeSans 224 90 0 0 chany_top_out_0[0]
port 156 nsew signal tristate
flabel metal2 s 5538 56200 5594 57000 0 FreeSans 224 90 0 0 chany_top_out_0[10]
port 157 nsew signal tristate
flabel metal2 s 5906 56200 5962 57000 0 FreeSans 224 90 0 0 chany_top_out_0[11]
port 158 nsew signal tristate
flabel metal2 s 6274 56200 6330 57000 0 FreeSans 224 90 0 0 chany_top_out_0[12]
port 159 nsew signal tristate
flabel metal2 s 6642 56200 6698 57000 0 FreeSans 224 90 0 0 chany_top_out_0[13]
port 160 nsew signal tristate
flabel metal2 s 7010 56200 7066 57000 0 FreeSans 224 90 0 0 chany_top_out_0[14]
port 161 nsew signal tristate
flabel metal2 s 7378 56200 7434 57000 0 FreeSans 224 90 0 0 chany_top_out_0[15]
port 162 nsew signal tristate
flabel metal2 s 7746 56200 7802 57000 0 FreeSans 224 90 0 0 chany_top_out_0[16]
port 163 nsew signal tristate
flabel metal2 s 8114 56200 8170 57000 0 FreeSans 224 90 0 0 chany_top_out_0[17]
port 164 nsew signal tristate
flabel metal2 s 8482 56200 8538 57000 0 FreeSans 224 90 0 0 chany_top_out_0[18]
port 165 nsew signal tristate
flabel metal2 s 8850 56200 8906 57000 0 FreeSans 224 90 0 0 chany_top_out_0[19]
port 166 nsew signal tristate
flabel metal2 s 2226 56200 2282 57000 0 FreeSans 224 90 0 0 chany_top_out_0[1]
port 167 nsew signal tristate
flabel metal2 s 9218 56200 9274 57000 0 FreeSans 224 90 0 0 chany_top_out_0[20]
port 168 nsew signal tristate
flabel metal2 s 9586 56200 9642 57000 0 FreeSans 224 90 0 0 chany_top_out_0[21]
port 169 nsew signal tristate
flabel metal2 s 9954 56200 10010 57000 0 FreeSans 224 90 0 0 chany_top_out_0[22]
port 170 nsew signal tristate
flabel metal2 s 10322 56200 10378 57000 0 FreeSans 224 90 0 0 chany_top_out_0[23]
port 171 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 chany_top_out_0[24]
port 172 nsew signal tristate
flabel metal2 s 11058 56200 11114 57000 0 FreeSans 224 90 0 0 chany_top_out_0[25]
port 173 nsew signal tristate
flabel metal2 s 11426 56200 11482 57000 0 FreeSans 224 90 0 0 chany_top_out_0[26]
port 174 nsew signal tristate
flabel metal2 s 11794 56200 11850 57000 0 FreeSans 224 90 0 0 chany_top_out_0[27]
port 175 nsew signal tristate
flabel metal2 s 12162 56200 12218 57000 0 FreeSans 224 90 0 0 chany_top_out_0[28]
port 176 nsew signal tristate
flabel metal2 s 12530 56200 12586 57000 0 FreeSans 224 90 0 0 chany_top_out_0[29]
port 177 nsew signal tristate
flabel metal2 s 2594 56200 2650 57000 0 FreeSans 224 90 0 0 chany_top_out_0[2]
port 178 nsew signal tristate
flabel metal2 s 2962 56200 3018 57000 0 FreeSans 224 90 0 0 chany_top_out_0[3]
port 179 nsew signal tristate
flabel metal2 s 3330 56200 3386 57000 0 FreeSans 224 90 0 0 chany_top_out_0[4]
port 180 nsew signal tristate
flabel metal2 s 3698 56200 3754 57000 0 FreeSans 224 90 0 0 chany_top_out_0[5]
port 181 nsew signal tristate
flabel metal2 s 4066 56200 4122 57000 0 FreeSans 224 90 0 0 chany_top_out_0[6]
port 182 nsew signal tristate
flabel metal2 s 4434 56200 4490 57000 0 FreeSans 224 90 0 0 chany_top_out_0[7]
port 183 nsew signal tristate
flabel metal2 s 4802 56200 4858 57000 0 FreeSans 224 90 0 0 chany_top_out_0[8]
port 184 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 chany_top_out_0[9]
port 185 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal3 s 0 35776 800 35896 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal3 s 0 38224 800 38344 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal3 s 0 25984 800 26104 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal3 s 0 43120 800 43240 0 FreeSans 480 0 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 prog_reset
port 200 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 reset
port 201 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 202 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 203 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 204 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 205 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 206 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 207 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 208 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 209 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 210 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 211 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 212 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 213 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 test_enable
port 214 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal input
flabel metal3 s 0 48016 800 48136 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal input
flabel metal3 s 0 50464 800 50584 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal input
flabel metal3 s 0 52912 800 53032 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal2 6026 24276 6026 24276 0 cby_0__1_.cby_0__1_.ccff_tail
rlabel metal2 6210 25092 6210 25092 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 4370 23154 4370 23154 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 4600 19482 4600 19482 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 3450 20978 3450 20978 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 7498 19720 7498 19720 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 13156 14450 13156 14450 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 11592 18598 11592 18598 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal2 8326 20060 8326 20060 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal2 9430 16388 9430 16388 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 16008 16626 16008 16626 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 13156 18802 13156 18802 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 10810 14246 10810 14246 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 6900 17102 6900 17102 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal1 14398 20978 14398 20978 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal2 12834 14348 12834 14348 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal2 8418 16354 8418 16354 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 14352 19278 14352 19278 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal2 12282 19822 12282 19822 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 8878 21590 8878 21590 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal1 12880 14586 12880 14586 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7912 21658 7912 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 6762 24174 6762 24174 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 13570 16864 13570 16864 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14260 18938 14260 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12742 23222 12742 23222 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11730 19448 11730 19448 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11638 16218 11638 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 11730 20230 11730 20230 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 8786 20876 8786 20876 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 9246 21658 9246 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9476 20570 9476 20570 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15226 15334 15226 15334 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9798 17306 9798 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 8280 17850 8280 17850 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14996 15470 14996 15470 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13662 18734 13662 18734 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13846 18394 13846 18394 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 11454 19040 11454 19040 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 11730 16048 11730 16048 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 13018 18632 13018 18632 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10350 16218 10350 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 11270 17238 11270 17238 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10350 16762 10350 16762 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13432 13226 13432 13226 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7084 17578 7084 17578 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 6302 18598 6302 18598 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13616 13294 13616 13294 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14306 18734 14306 18734 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12742 17034 12742 17034 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9338 19482 9338 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12236 13498 12236 13498 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10580 16150 10580 16150 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8372 17646 8372 17646 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8878 16762 8878 16762 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8142 16218 8142 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 12190 16660 12190 16660 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 6256 22746 6256 22746 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 4784 22406 4784 22406 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 12466 18734 12466 18734 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13984 20026 13984 20026 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12052 21658 12052 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10442 18190 10442 18190 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11408 18394 11408 18394 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10810 21658 10810 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7590 21114 7590 21114 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8326 22746 8326 22746 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8694 21386 8694 21386 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 4278 24956 4278 24956 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 3036 25806 3036 25806 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 3404 25738 3404 25738 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel via1 3795 28186 3795 28186 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 4324 20502 4324 20502 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 2254 20876 2254 20876 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 3036 23290 3036 23290 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 3335 27098 3335 27098 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 5796 20230 5796 20230 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 2254 19380 2254 19380 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 2254 23052 2254 23052 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 4071 25126 4071 25126 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 3542 20910 3542 20910 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 3036 21114 3036 21114 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 4301 23086 4301 23086 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal3 2338 55420 2338 55420 0 ccff_head
rlabel metal3 2062 1564 2062 1564 0 ccff_head_0
rlabel metal2 24978 2363 24978 2363 0 ccff_tail
rlabel metal1 1794 49266 1794 49266 0 ccff_tail_0
rlabel metal2 25346 24871 25346 24871 0 chanx_right_in[0]
rlabel via2 25346 34187 25346 34187 0 chanx_right_in[10]
rlabel via2 25346 35037 25346 35037 0 chanx_right_in[11]
rlabel metal2 25346 35989 25346 35989 0 chanx_right_in[12]
rlabel metal2 25346 36703 25346 36703 0 chanx_right_in[13]
rlabel metal2 25346 37349 25346 37349 0 chanx_right_in[14]
rlabel metal2 25346 38607 25346 38607 0 chanx_right_in[15]
rlabel metal1 24794 38930 24794 38930 0 chanx_right_in[16]
rlabel metal1 25070 40494 25070 40494 0 chanx_right_in[17]
rlabel metal1 24794 41514 24794 41514 0 chanx_right_in[18]
rlabel via2 25346 41565 25346 41565 0 chanx_right_in[19]
rlabel metal2 25530 26163 25530 26163 0 chanx_right_in[1]
rlabel metal1 24702 42534 24702 42534 0 chanx_right_in[20]
rlabel metal2 25346 43401 25346 43401 0 chanx_right_in[21]
rlabel metal2 25530 44353 25530 44353 0 chanx_right_in[22]
rlabel metal3 25952 44812 25952 44812 0 chanx_right_in[23]
rlabel metal1 24702 45798 24702 45798 0 chanx_right_in[24]
rlabel metal1 24840 46954 24840 46954 0 chanx_right_in[25]
rlabel metal2 25530 47889 25530 47889 0 chanx_right_in[26]
rlabel via2 25346 48093 25346 48093 0 chanx_right_in[27]
rlabel metal2 25346 49045 25346 49045 0 chanx_right_in[28]
rlabel metal2 25346 49759 25346 49759 0 chanx_right_in[29]
rlabel metal2 24150 28407 24150 28407 0 chanx_right_in[2]
rlabel metal1 24058 28492 24058 28492 0 chanx_right_in[3]
rlabel via2 25530 29291 25530 29291 0 chanx_right_in[4]
rlabel metal2 25346 29869 25346 29869 0 chanx_right_in[5]
rlabel metal2 25346 31127 25346 31127 0 chanx_right_in[6]
rlabel via2 25346 31773 25346 31773 0 chanx_right_in[7]
rlabel metal2 25346 32725 25346 32725 0 chanx_right_in[8]
rlabel metal1 25392 32402 25392 32402 0 chanx_right_in[9]
rlabel metal3 25676 9724 25676 9724 0 chanx_right_out[10]
rlabel metal2 24702 9469 24702 9469 0 chanx_right_out[11]
rlabel metal1 23920 9486 23920 9486 0 chanx_right_out[12]
rlabel metal2 24794 11373 24794 11373 0 chanx_right_out[13]
rlabel metal3 25952 12988 25952 12988 0 chanx_right_out[14]
rlabel metal2 23322 13311 23322 13311 0 chanx_right_out[15]
rlabel metal2 24794 13685 24794 13685 0 chanx_right_out[16]
rlabel metal3 25676 15436 25676 15436 0 chanx_right_out[17]
rlabel metal2 24702 15045 24702 15045 0 chanx_right_out[18]
rlabel metal2 24794 15997 24794 15997 0 chanx_right_out[19]
rlabel metal3 23882 2380 23882 2380 0 chanx_right_out[1]
rlabel metal1 24104 17238 24104 17238 0 chanx_right_out[20]
rlabel metal1 23920 16014 23920 16014 0 chanx_right_out[21]
rlabel metal1 23874 17102 23874 17102 0 chanx_right_out[22]
rlabel metal1 24426 19890 24426 19890 0 chanx_right_out[23]
rlabel metal1 23368 20502 23368 20502 0 chanx_right_out[24]
rlabel metal1 24380 20978 24380 20978 0 chanx_right_out[25]
rlabel metal3 25538 22780 25538 22780 0 chanx_right_out[26]
rlabel metal2 23874 23375 23874 23375 0 chanx_right_out[27]
rlabel metal1 24380 24242 24380 24242 0 chanx_right_out[28]
rlabel metal2 25162 25517 25162 25517 0 chanx_right_out[29]
rlabel metal3 24848 3196 24848 3196 0 chanx_right_out[2]
rlabel metal2 22126 4063 22126 4063 0 chanx_right_out[3]
rlabel metal3 25446 4828 25446 4828 0 chanx_right_out[4]
rlabel metal2 24794 4845 24794 4845 0 chanx_right_out[5]
rlabel metal3 25722 6460 25722 6460 0 chanx_right_out[6]
rlabel metal2 24656 6732 24656 6732 0 chanx_right_out[7]
rlabel metal3 25584 8092 25584 8092 0 chanx_right_out[8]
rlabel metal2 25162 8177 25162 8177 0 chanx_right_out[9]
rlabel metal1 1610 4998 1610 4998 0 chany_bottom_in[0]
rlabel metal2 5382 4556 5382 4556 0 chany_bottom_in[10]
rlabel metal1 5934 2278 5934 2278 0 chany_bottom_in[11]
rlabel metal1 5474 3026 5474 3026 0 chany_bottom_in[12]
rlabel metal2 6486 1761 6486 1761 0 chany_bottom_in[13]
rlabel metal2 6854 3706 6854 3706 0 chany_bottom_in[14]
rlabel metal1 7038 3026 7038 3026 0 chany_bottom_in[15]
rlabel metal1 7636 2414 7636 2414 0 chany_bottom_in[16]
rlabel metal2 7912 1972 7912 1972 0 chany_bottom_in[17]
rlabel metal1 7498 2380 7498 2380 0 chany_bottom_in[18]
rlabel metal2 8694 1761 8694 1761 0 chany_bottom_in[19]
rlabel metal1 1886 3502 1886 3502 0 chany_bottom_in[1]
rlabel metal2 9062 3774 9062 3774 0 chany_bottom_in[20]
rlabel metal1 9890 4114 9890 4114 0 chany_bottom_in[21]
rlabel metal1 9982 3502 9982 3502 0 chany_bottom_in[22]
rlabel metal1 9752 2414 9752 2414 0 chany_bottom_in[23]
rlabel metal2 10350 3502 10350 3502 0 chany_bottom_in[24]
rlabel metal1 10948 3570 10948 3570 0 chany_bottom_in[25]
rlabel metal1 11500 4114 11500 4114 0 chany_bottom_in[26]
rlabel metal1 11776 4590 11776 4590 0 chany_bottom_in[27]
rlabel metal1 11914 2448 11914 2448 0 chany_bottom_in[28]
rlabel metal1 10350 2516 10350 2516 0 chany_bottom_in[29]
rlabel metal2 2162 4318 2162 4318 0 chany_bottom_in[2]
rlabel metal2 2806 3230 2806 3230 0 chany_bottom_in[3]
rlabel metal2 3266 2618 3266 2618 0 chany_bottom_in[4]
rlabel metal1 1702 2448 1702 2448 0 chany_bottom_in[5]
rlabel metal1 4186 4114 4186 4114 0 chany_bottom_in[6]
rlabel metal1 2806 2380 2806 2380 0 chany_bottom_in[7]
rlabel metal2 4646 1588 4646 1588 0 chany_bottom_in[8]
rlabel metal1 4830 3502 4830 3502 0 chany_bottom_in[9]
rlabel metal1 12788 3570 12788 3570 0 chany_bottom_out[0]
rlabel metal1 16882 4046 16882 4046 0 chany_bottom_out[10]
rlabel metal1 18952 2482 18952 2482 0 chany_bottom_out[11]
rlabel metal1 18170 2890 18170 2890 0 chany_bottom_out[12]
rlabel metal1 18354 4046 18354 4046 0 chany_bottom_out[13]
rlabel metal1 18906 3570 18906 3570 0 chany_bottom_out[14]
rlabel metal2 18262 959 18262 959 0 chany_bottom_out[15]
rlabel metal1 19274 3366 19274 3366 0 chany_bottom_out[16]
rlabel metal1 20378 3638 20378 3638 0 chany_bottom_out[17]
rlabel metal1 19872 5270 19872 5270 0 chany_bottom_out[18]
rlabel metal1 20746 3434 20746 3434 0 chany_bottom_out[19]
rlabel metal2 13110 823 13110 823 0 chany_bottom_out[1]
rlabel metal2 20102 2404 20102 2404 0 chany_bottom_out[20]
rlabel metal1 20746 5746 20746 5746 0 chany_bottom_out[21]
rlabel metal2 22494 3978 22494 3978 0 chany_bottom_out[22]
rlabel metal1 19964 5610 19964 5610 0 chany_bottom_out[23]
rlabel metal2 21574 3254 21574 3254 0 chany_bottom_out[24]
rlabel metal2 21942 3492 21942 3492 0 chany_bottom_out[25]
rlabel metal1 22448 7310 22448 7310 0 chany_bottom_out[26]
rlabel metal2 22678 1962 22678 1962 0 chany_bottom_out[27]
rlabel metal2 23046 1639 23046 1639 0 chany_bottom_out[28]
rlabel metal2 23414 1860 23414 1860 0 chany_bottom_out[29]
rlabel metal1 13754 4046 13754 4046 0 chany_bottom_out[2]
rlabel metal2 13846 1554 13846 1554 0 chany_bottom_out[3]
rlabel metal1 14490 2958 14490 2958 0 chany_bottom_out[4]
rlabel metal2 14582 1622 14582 1622 0 chany_bottom_out[5]
rlabel metal1 15226 3570 15226 3570 0 chany_bottom_out[6]
rlabel metal2 15318 1622 15318 1622 0 chany_bottom_out[7]
rlabel metal1 16514 2958 16514 2958 0 chany_bottom_out[8]
rlabel metal1 16698 3570 16698 3570 0 chany_bottom_out[9]
rlabel metal1 11914 54196 11914 54196 0 chany_top_in_0[0]
rlabel metal2 17986 53958 17986 53958 0 chany_top_in_0[10]
rlabel metal1 17342 53550 17342 53550 0 chany_top_in_0[11]
rlabel metal1 17480 51986 17480 51986 0 chany_top_in_0[12]
rlabel metal1 18262 53686 18262 53686 0 chany_top_in_0[13]
rlabel metal2 18262 56236 18262 56236 0 chany_top_in_0[14]
rlabel metal1 18722 53754 18722 53754 0 chany_top_in_0[15]
rlabel metal2 18814 55711 18814 55711 0 chany_top_in_0[16]
rlabel metal1 20562 54128 20562 54128 0 chany_top_in_0[17]
rlabel metal1 20056 53550 20056 53550 0 chany_top_in_0[18]
rlabel metal1 20010 53074 20010 53074 0 chany_top_in_0[19]
rlabel metal2 13294 55711 13294 55711 0 chany_top_in_0[1]
rlabel metal1 20424 51986 20424 51986 0 chany_top_in_0[20]
rlabel metal2 20654 55711 20654 55711 0 chany_top_in_0[21]
rlabel metal1 21344 53550 21344 53550 0 chany_top_in_0[22]
rlabel metal1 23138 54128 23138 54128 0 chany_top_in_0[23]
rlabel metal1 22586 52496 22586 52496 0 chany_top_in_0[24]
rlabel metal2 22126 55711 22126 55711 0 chany_top_in_0[25]
rlabel metal1 22770 53584 22770 53584 0 chany_top_in_0[26]
rlabel metal1 23092 51986 23092 51986 0 chany_top_in_0[27]
rlabel metal2 23230 55711 23230 55711 0 chany_top_in_0[28]
rlabel metal1 23920 51986 23920 51986 0 chany_top_in_0[29]
rlabel metal1 13984 54230 13984 54230 0 chany_top_in_0[2]
rlabel metal1 14076 54298 14076 54298 0 chany_top_in_0[3]
rlabel metal2 14582 56236 14582 56236 0 chany_top_in_0[4]
rlabel metal1 14674 54298 14674 54298 0 chany_top_in_0[5]
rlabel metal1 15272 53550 15272 53550 0 chany_top_in_0[6]
rlabel metal1 17158 54162 17158 54162 0 chany_top_in_0[7]
rlabel metal1 16008 51986 16008 51986 0 chany_top_in_0[8]
rlabel metal1 16330 52666 16330 52666 0 chany_top_in_0[9]
rlabel metal1 2714 52666 2714 52666 0 chany_top_out_0[0]
rlabel metal1 5566 53652 5566 53652 0 chany_top_out_0[10]
rlabel metal1 4600 54094 4600 54094 0 chany_top_out_0[11]
rlabel metal1 6072 53142 6072 53142 0 chany_top_out_0[12]
rlabel metal1 6624 52462 6624 52462 0 chany_top_out_0[13]
rlabel metal1 7314 51442 7314 51442 0 chany_top_out_0[14]
rlabel metal1 6992 53618 6992 53618 0 chany_top_out_0[15]
rlabel metal2 7774 54376 7774 54376 0 chany_top_out_0[16]
rlabel metal2 7958 56236 7958 56236 0 chany_top_out_0[17]
rlabel metal2 8510 54070 8510 54070 0 chany_top_out_0[18]
rlabel metal1 8648 53618 8648 53618 0 chany_top_out_0[19]
rlabel metal1 2852 53686 2852 53686 0 chany_top_out_0[1]
rlabel metal1 9200 53142 9200 53142 0 chany_top_out_0[20]
rlabel metal2 9706 53550 9706 53550 0 chany_top_out_0[21]
rlabel metal1 9982 54264 9982 54264 0 chany_top_out_0[22]
rlabel metal2 10350 54614 10350 54614 0 chany_top_out_0[23]
rlabel metal1 10994 52530 10994 52530 0 chany_top_out_0[24]
rlabel metal2 11086 54920 11086 54920 0 chany_top_out_0[25]
rlabel metal1 11224 54230 11224 54230 0 chany_top_out_0[26]
rlabel metal1 12098 53006 12098 53006 0 chany_top_out_0[27]
rlabel metal1 12466 53618 12466 53618 0 chany_top_out_0[28]
rlabel metal1 12696 54094 12696 54094 0 chany_top_out_0[29]
rlabel metal2 2714 52972 2714 52972 0 chany_top_out_0[2]
rlabel metal2 2990 55711 2990 55711 0 chany_top_out_0[3]
rlabel metal2 3358 54070 3358 54070 0 chany_top_out_0[4]
rlabel metal1 3496 52530 3496 52530 0 chany_top_out_0[5]
rlabel metal2 4232 52972 4232 52972 0 chany_top_out_0[6]
rlabel metal1 4232 53142 4232 53142 0 chany_top_out_0[7]
rlabel metal2 4830 55711 4830 55711 0 chany_top_out_0[8]
rlabel metal2 5382 56236 5382 56236 0 chany_top_out_0[9]
rlabel metal1 19688 42058 19688 42058 0 clknet_0_prog_clk
rlabel metal1 8004 13362 8004 13362 0 clknet_4_0_0_prog_clk
rlabel metal1 6026 39474 6026 39474 0 clknet_4_10_0_prog_clk
rlabel metal1 9200 41242 9200 41242 0 clknet_4_11_0_prog_clk
rlabel metal1 19826 35122 19826 35122 0 clknet_4_12_0_prog_clk
rlabel metal1 22862 33490 22862 33490 0 clknet_4_13_0_prog_clk
rlabel metal1 19458 42126 19458 42126 0 clknet_4_14_0_prog_clk
rlabel metal1 23184 42126 23184 42126 0 clknet_4_15_0_prog_clk
rlabel metal2 11362 17340 11362 17340 0 clknet_4_1_0_prog_clk
rlabel metal1 9016 19890 9016 19890 0 clknet_4_2_0_prog_clk
rlabel metal1 9890 20842 9890 20842 0 clknet_4_3_0_prog_clk
rlabel metal1 18630 18190 18630 18190 0 clknet_4_4_0_prog_clk
rlabel metal1 19044 12750 19044 12750 0 clknet_4_5_0_prog_clk
rlabel metal2 15410 26180 15410 26180 0 clknet_4_6_0_prog_clk
rlabel metal1 19688 20978 19688 20978 0 clknet_4_7_0_prog_clk
rlabel metal1 6854 37162 6854 37162 0 clknet_4_8_0_prog_clk
rlabel metal1 12926 31178 12926 31178 0 clknet_4_9_0_prog_clk
rlabel metal3 1004 13804 1004 13804 0 gfpga_pad_io_soc_dir[0]
rlabel metal3 1004 16252 1004 16252 0 gfpga_pad_io_soc_dir[1]
rlabel metal3 1004 18700 1004 18700 0 gfpga_pad_io_soc_dir[2]
rlabel metal3 1004 21148 1004 21148 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 1426 33490 1426 33490 0 gfpga_pad_io_soc_in[0]
rlabel metal2 1610 36346 1610 36346 0 gfpga_pad_io_soc_in[1]
rlabel metal1 1472 38318 1472 38318 0 gfpga_pad_io_soc_in[2]
rlabel metal1 1472 41106 1472 41106 0 gfpga_pad_io_soc_in[3]
rlabel metal3 1004 23596 1004 23596 0 gfpga_pad_io_soc_out[0]
rlabel metal2 2806 26163 2806 26163 0 gfpga_pad_io_soc_out[1]
rlabel metal3 1004 28492 1004 28492 0 gfpga_pad_io_soc_out[2]
rlabel metal3 1004 30940 1004 30940 0 gfpga_pad_io_soc_out[3]
rlabel metal1 1426 43282 1426 43282 0 isol_n
rlabel metal1 1656 51034 1656 51034 0 net1
rlabel metal1 20194 38318 20194 38318 0 net10
rlabel metal1 18860 41446 18860 41446 0 net100
rlabel metal2 17434 43520 17434 43520 0 net101
rlabel metal1 24334 42670 24334 42670 0 net102
rlabel metal1 25530 51782 25530 51782 0 net103
rlabel metal1 24242 52870 24242 52870 0 net104
rlabel metal2 23736 45540 23736 45540 0 net105
rlabel metal1 25438 53550 25438 53550 0 net106
rlabel metal1 10810 40494 10810 40494 0 net107
rlabel metal1 14904 37434 14904 37434 0 net108
rlabel metal1 15272 40426 15272 40426 0 net109
rlabel metal1 20148 35734 20148 35734 0 net11
rlabel metal1 7682 52496 7682 52496 0 net110
rlabel metal1 18124 6290 18124 6290 0 net111
rlabel metal2 10902 37995 10902 37995 0 net112
rlabel metal1 22678 9996 22678 9996 0 net113
rlabel metal2 23966 9758 23966 9758 0 net114
rlabel metal1 23966 9588 23966 9588 0 net115
rlabel metal1 23828 10642 23828 10642 0 net116
rlabel metal2 21758 15164 21758 15164 0 net117
rlabel metal1 22402 12818 22402 12818 0 net118
rlabel metal2 21482 15504 21482 15504 0 net119
rlabel metal1 21022 41106 21022 41106 0 net12
rlabel metal1 23552 15470 23552 15470 0 net120
rlabel metal1 23920 13906 23920 13906 0 net121
rlabel metal2 24150 18496 24150 18496 0 net122
rlabel metal1 20286 7344 20286 7344 0 net123
rlabel metal2 22172 23052 22172 23052 0 net124
rlabel metal1 24150 16116 24150 16116 0 net125
rlabel metal2 23966 21148 23966 21148 0 net126
rlabel metal1 24242 19822 24242 19822 0 net127
rlabel metal1 22954 20434 22954 20434 0 net128
rlabel metal2 22678 21495 22678 21495 0 net129
rlabel metal2 16054 39746 16054 39746 0 net13
rlabel metal1 24702 20434 24702 20434 0 net130
rlabel metal1 22862 23052 22862 23052 0 net131
rlabel metal1 23092 24174 23092 24174 0 net132
rlabel metal1 23920 25874 23920 25874 0 net133
rlabel metal1 23782 4726 23782 4726 0 net134
rlabel metal2 17802 4998 17802 4998 0 net135
rlabel metal1 23184 7854 23184 7854 0 net136
rlabel metal2 24702 5372 24702 5372 0 net137
rlabel metal1 22678 7718 22678 7718 0 net138
rlabel metal1 24426 9894 24426 9894 0 net139
rlabel metal1 18078 24718 18078 24718 0 net14
rlabel metal2 22586 5100 22586 5100 0 net140
rlabel metal1 23690 7378 23690 7378 0 net141
rlabel metal2 12696 13838 12696 13838 0 net142
rlabel metal1 16238 14790 16238 14790 0 net143
rlabel metal2 19550 2587 19550 2587 0 net144
rlabel metal1 18722 2618 18722 2618 0 net145
rlabel via3 18469 19380 18469 19380 0 net146
rlabel metal1 17526 14858 17526 14858 0 net147
rlabel metal1 19872 2550 19872 2550 0 net148
rlabel metal1 19044 4590 19044 4590 0 net149
rlabel metal1 23598 42670 23598 42670 0 net15
rlabel metal1 20194 14586 20194 14586 0 net150
rlabel metal1 19642 18598 19642 18598 0 net151
rlabel metal2 21298 6460 21298 6460 0 net152
rlabel metal1 13938 13770 13938 13770 0 net153
rlabel metal1 22310 4114 22310 4114 0 net154
rlabel metal1 20516 13838 20516 13838 0 net155
rlabel metal2 22218 6051 22218 6051 0 net156
rlabel metal2 17710 7514 17710 7514 0 net157
rlabel metal2 20654 6460 20654 6460 0 net158
rlabel metal2 22034 8942 22034 8942 0 net159
rlabel metal3 22287 43180 22287 43180 0 net16
rlabel metal2 20746 7854 20746 7854 0 net160
rlabel metal1 20700 6290 20700 6290 0 net161
rlabel metal2 20838 7242 20838 7242 0 net162
rlabel metal1 18032 4590 18032 4590 0 net163
rlabel metal1 13708 13838 13708 13838 0 net164
rlabel metal2 12466 6460 12466 6460 0 net165
rlabel metal1 14122 12682 14122 12682 0 net166
rlabel metal2 14674 7548 14674 7548 0 net167
rlabel metal1 15824 15878 15824 15878 0 net168
rlabel metal2 16882 6154 16882 6154 0 net169
rlabel metal1 24748 45390 24748 45390 0 net17
rlabel metal2 17066 7276 17066 7276 0 net170
rlabel metal1 16192 3434 16192 3434 0 net171
rlabel metal2 1978 45526 1978 45526 0 net172
rlabel via2 2254 53533 2254 53533 0 net173
rlabel metal1 2300 54162 2300 54162 0 net174
rlabel metal1 6348 44982 6348 44982 0 net175
rlabel metal1 5704 52462 5704 52462 0 net176
rlabel metal1 8142 44438 8142 44438 0 net177
rlabel metal1 6210 53550 6210 53550 0 net178
rlabel metal1 8326 45050 8326 45050 0 net179
rlabel metal1 24518 46546 24518 46546 0 net18
rlabel metal1 6670 43350 6670 43350 0 net180
rlabel metal1 8050 51918 8050 51918 0 net181
rlabel metal1 8004 53550 8004 53550 0 net182
rlabel metal1 2254 50252 2254 50252 0 net183
rlabel metal1 7774 53074 7774 53074 0 net184
rlabel metal1 10396 44506 10396 44506 0 net185
rlabel metal1 7406 54128 7406 54128 0 net186
rlabel metal1 9568 53074 9568 53074 0 net187
rlabel metal1 10212 52462 10212 52462 0 net188
rlabel metal1 11362 53550 11362 53550 0 net189
rlabel metal1 23782 45934 23782 45934 0 net19
rlabel metal1 10120 51578 10120 51578 0 net190
rlabel metal1 11822 52122 11822 52122 0 net191
rlabel metal2 12650 53108 12650 53108 0 net192
rlabel metal2 12374 53142 12374 53142 0 net193
rlabel metal1 2898 50830 2898 50830 0 net194
rlabel metal1 3082 51374 3082 51374 0 net195
rlabel metal1 3404 51986 3404 51986 0 net196
rlabel metal1 3726 52462 3726 52462 0 net197
rlabel metal1 4876 50898 4876 50898 0 net198
rlabel metal1 3772 53074 3772 53074 0 net199
rlabel metal2 2530 5882 2530 5882 0 net2
rlabel metal2 19090 39712 19090 39712 0 net20
rlabel metal2 7222 51646 7222 51646 0 net200
rlabel metal1 5474 51340 5474 51340 0 net201
rlabel metal2 1794 14892 1794 14892 0 net202
rlabel metal1 1794 19482 1794 19482 0 net203
rlabel metal2 1794 19754 1794 19754 0 net204
rlabel metal1 1840 21522 1840 21522 0 net205
rlabel metal1 1932 22746 1932 22746 0 net206
rlabel metal1 1932 26350 1932 26350 0 net207
rlabel metal1 1978 26010 1978 26010 0 net208
rlabel metal1 2024 28186 2024 28186 0 net209
rlabel metal1 24610 47634 24610 47634 0 net21
rlabel metal1 24472 2482 24472 2482 0 net210
rlabel metal2 17618 21182 17618 21182 0 net211
rlabel metal1 12926 28186 12926 28186 0 net212
rlabel metal2 21482 33728 21482 33728 0 net213
rlabel metal1 24242 23086 24242 23086 0 net214
rlabel metal1 14904 37842 14904 37842 0 net215
rlabel metal1 17158 21998 17158 21998 0 net216
rlabel metal2 20930 29376 20930 29376 0 net217
rlabel metal1 16928 36074 16928 36074 0 net218
rlabel metal1 17986 36890 17986 36890 0 net219
rlabel metal1 19182 42330 19182 42330 0 net22
rlabel metal1 17066 37978 17066 37978 0 net220
rlabel metal1 14536 39066 14536 39066 0 net221
rlabel metal1 13432 37230 13432 37230 0 net222
rlabel metal1 23460 39338 23460 39338 0 net223
rlabel metal1 12788 32402 12788 32402 0 net224
rlabel metal1 11270 30226 11270 30226 0 net225
rlabel metal1 13018 24242 13018 24242 0 net226
rlabel metal2 11822 25534 11822 25534 0 net227
rlabel metal2 9430 25602 9430 25602 0 net228
rlabel metal2 9154 26690 9154 26690 0 net229
rlabel metal1 18032 42670 18032 42670 0 net23
rlabel metal1 7958 24922 7958 24922 0 net230
rlabel metal1 10074 24820 10074 24820 0 net231
rlabel metal1 6394 9554 6394 9554 0 net232
rlabel metal1 14950 11186 14950 11186 0 net233
rlabel metal1 20700 32878 20700 32878 0 net234
rlabel metal2 17250 13056 17250 13056 0 net235
rlabel metal1 18768 15130 18768 15130 0 net236
rlabel metal2 20470 16830 20470 16830 0 net237
rlabel metal1 22356 15130 22356 15130 0 net238
rlabel metal1 20056 16082 20056 16082 0 net239
rlabel metal1 23092 49946 23092 49946 0 net24
rlabel metal1 21758 12206 21758 12206 0 net240
rlabel metal1 19596 10778 19596 10778 0 net241
rlabel metal1 19642 13294 19642 13294 0 net242
rlabel metal1 23046 34646 23046 34646 0 net243
rlabel metal2 22034 41344 22034 41344 0 net244
rlabel metal1 9936 37842 9936 37842 0 net245
rlabel metal1 7912 30770 7912 30770 0 net246
rlabel metal1 7406 32538 7406 32538 0 net247
rlabel metal1 13800 42194 13800 42194 0 net248
rlabel metal2 9798 33150 9798 33150 0 net249
rlabel metal1 15042 30634 15042 30634 0 net25
rlabel metal2 5382 32980 5382 32980 0 net250
rlabel metal1 8280 38318 8280 38318 0 net251
rlabel metal1 11270 37978 11270 37978 0 net252
rlabel metal1 10902 39066 10902 39066 0 net253
rlabel metal1 14582 35802 14582 35802 0 net254
rlabel metal1 9476 31450 9476 31450 0 net255
rlabel metal2 11730 23358 11730 23358 0 net256
rlabel metal1 12880 20570 12880 20570 0 net257
rlabel metal1 9568 16558 9568 16558 0 net258
rlabel metal1 9844 23834 9844 23834 0 net259
rlabel metal1 16790 31926 16790 31926 0 net26
rlabel metal2 13938 22100 13938 22100 0 net260
rlabel metal1 14076 24242 14076 24242 0 net261
rlabel metal1 20332 26962 20332 26962 0 net262
rlabel metal2 21298 25534 21298 25534 0 net263
rlabel metal2 17250 29716 17250 29716 0 net264
rlabel metal2 24610 2890 24610 2890 0 net265
rlabel metal1 24242 41446 24242 41446 0 net266
rlabel metal1 24334 3502 24334 3502 0 net267
rlabel metal1 25300 2618 25300 2618 0 net268
rlabel metal1 23092 11730 23092 11730 0 net269
rlabel metal1 19734 36006 19734 36006 0 net27
rlabel metal2 20746 17408 20746 17408 0 net270
rlabel metal2 23138 3332 23138 3332 0 net271
rlabel metal1 1702 53006 1702 53006 0 net272
rlabel metal1 4462 51238 4462 51238 0 net273
rlabel metal2 1794 4284 1794 4284 0 net274
rlabel metal1 4048 6426 4048 6426 0 net275
rlabel metal1 5106 3162 5106 3162 0 net276
rlabel metal2 1794 33082 1794 33082 0 net277
rlabel metal1 3082 19380 3082 19380 0 net278
rlabel metal1 2024 36006 2024 36006 0 net279
rlabel metal1 19596 38250 19596 38250 0 net28
rlabel metal1 4646 18734 4646 18734 0 net280
rlabel metal2 1794 38012 1794 38012 0 net281
rlabel metal1 4324 18258 4324 18258 0 net282
rlabel metal2 1794 40698 1794 40698 0 net283
rlabel metal1 3910 17170 3910 17170 0 net284
rlabel metal1 18630 52462 18630 52462 0 net285
rlabel metal1 14030 52394 14030 52394 0 net286
rlabel metal1 21022 53074 21022 53074 0 net287
rlabel metal2 17526 53550 17526 53550 0 net288
rlabel metal1 2116 3706 2116 3706 0 net289
rlabel metal1 18906 35802 18906 35802 0 net29
rlabel metal2 22034 53244 22034 53244 0 net290
rlabel metal1 19458 52496 19458 52496 0 net291
rlabel metal1 14122 52054 14122 52054 0 net292
rlabel metal2 7222 4352 7222 4352 0 net293
rlabel metal2 19366 53550 19366 53550 0 net294
rlabel metal1 15732 54162 15732 54162 0 net295
rlabel metal2 17618 52938 17618 52938 0 net296
rlabel metal1 3726 2618 3726 2618 0 net297
rlabel metal2 15594 52938 15594 52938 0 net298
rlabel metal1 3174 3706 3174 3706 0 net299
rlabel metal1 20010 24718 20010 24718 0 net3
rlabel metal1 21528 33966 21528 33966 0 net30
rlabel metal1 22770 53108 22770 53108 0 net300
rlabel metal1 2990 4080 2990 4080 0 net301
rlabel metal1 8464 3162 8464 3162 0 net302
rlabel metal2 14306 52938 14306 52938 0 net303
rlabel metal1 7452 2550 7452 2550 0 net304
rlabel metal1 17296 53074 17296 53074 0 net305
rlabel metal2 6026 4658 6026 4658 0 net306
rlabel metal2 16882 52938 16882 52938 0 net307
rlabel metal2 20194 52938 20194 52938 0 net308
rlabel metal2 2346 3876 2346 3876 0 net309
rlabel metal1 16238 37638 16238 37638 0 net31
rlabel metal1 21896 52462 21896 52462 0 net310
rlabel metal2 23506 53244 23506 53244 0 net311
rlabel metal1 1702 6256 1702 6256 0 net312
rlabel metal2 20930 52938 20930 52938 0 net313
rlabel metal1 5152 3706 5152 3706 0 net314
rlabel metal2 8602 3910 8602 3910 0 net315
rlabel metal1 9154 3468 9154 3468 0 net316
rlabel metal1 4922 2550 4922 2550 0 net317
rlabel metal2 4646 3196 4646 3196 0 net318
rlabel metal1 8694 4080 8694 4080 0 net319
rlabel metal2 20194 32351 20194 32351 0 net32
rlabel metal1 9752 4590 9752 4590 0 net320
rlabel metal2 11730 3468 11730 3468 0 net321
rlabel metal1 6072 3706 6072 3706 0 net322
rlabel metal1 1978 42670 1978 42670 0 net323
rlabel metal1 4554 5236 4554 5236 0 net324
rlabel metal2 6578 53244 6578 53244 0 net325
rlabel metal2 1794 51884 1794 51884 0 net326
rlabel metal2 4002 51578 4002 51578 0 net327
rlabel metal1 1610 4624 1610 4624 0 net328
rlabel metal2 2438 5202 2438 5202 0 net329
rlabel metal1 4416 5338 4416 5338 0 net33
rlabel metal1 3266 5882 3266 5882 0 net330
rlabel metal2 10304 18292 10304 18292 0 net34
rlabel metal4 12604 37150 12604 37150 0 net35
rlabel metal2 16146 3876 16146 3876 0 net36
rlabel metal1 12926 37298 12926 37298 0 net37
rlabel metal2 13846 38777 13846 38777 0 net38
rlabel metal1 4186 2312 4186 2312 0 net39
rlabel metal2 20148 33660 20148 33660 0 net4
rlabel metal1 12788 2278 12788 2278 0 net40
rlabel via2 16698 36771 16698 36771 0 net41
rlabel metal1 15732 36074 15732 36074 0 net42
rlabel metal1 19044 37842 19044 37842 0 net43
rlabel metal1 5980 18054 5980 18054 0 net44
rlabel via2 14766 19669 14766 19669 0 net45
rlabel metal1 13984 21114 13984 21114 0 net46
rlabel metal1 14398 20230 14398 20230 0 net47
rlabel metal1 13248 18122 13248 18122 0 net48
rlabel metal2 19366 16762 19366 16762 0 net49
rlabel metal2 20470 30940 20470 30940 0 net5
rlabel metal1 15364 16626 15364 16626 0 net50
rlabel metal2 12466 43724 12466 43724 0 net51
rlabel metal1 18216 15062 18216 15062 0 net52
rlabel metal1 13846 2618 13846 2618 0 net53
rlabel metal1 11638 2346 11638 2346 0 net54
rlabel metal1 2024 20842 2024 20842 0 net55
rlabel metal1 8924 19346 8924 19346 0 net56
rlabel metal1 10304 15334 10304 15334 0 net57
rlabel via2 8694 19669 8694 19669 0 net58
rlabel metal1 3864 3910 3864 3910 0 net59
rlabel metal1 21436 31722 21436 31722 0 net6
rlabel metal2 9430 17850 9430 17850 0 net60
rlabel metal1 5014 2516 5014 2516 0 net61
rlabel metal1 12926 36006 12926 36006 0 net62
rlabel metal1 12236 53958 12236 53958 0 net63
rlabel metal2 16974 43180 16974 43180 0 net64
rlabel metal1 15824 43078 15824 43078 0 net65
rlabel metal2 18446 49810 18446 49810 0 net66
rlabel metal1 18630 48246 18630 48246 0 net67
rlabel metal2 18538 50048 18538 50048 0 net68
rlabel metal1 16882 44846 16882 44846 0 net69
rlabel metal2 20102 36822 20102 36822 0 net7
rlabel metal2 18630 49436 18630 49436 0 net70
rlabel metal1 19550 46138 19550 46138 0 net71
rlabel metal1 21206 45934 21206 45934 0 net72
rlabel metal2 21666 50082 21666 50082 0 net73
rlabel metal1 13616 52462 13616 52462 0 net74
rlabel metal2 20194 48892 20194 48892 0 net75
rlabel via2 21666 43061 21666 43061 0 net76
rlabel metal1 22448 43622 22448 43622 0 net77
rlabel metal1 22632 46682 22632 46682 0 net78
rlabel metal2 21390 49334 21390 49334 0 net79
rlabel metal2 20838 37808 20838 37808 0 net8
rlabel metal1 22586 47022 22586 47022 0 net80
rlabel metal3 23759 52564 23759 52564 0 net81
rlabel metal1 22448 43418 22448 43418 0 net82
rlabel metal1 22908 52598 22908 52598 0 net83
rlabel metal2 22770 49266 22770 49266 0 net84
rlabel metal1 14076 51850 14076 51850 0 net85
rlabel metal2 13570 14025 13570 14025 0 net86
rlabel metal1 14766 51850 14766 51850 0 net87
rlabel metal1 15732 53958 15732 53958 0 net88
rlabel metal1 14444 12886 14444 12886 0 net89
rlabel metal1 21390 36040 21390 36040 0 net9
rlabel via3 16445 52564 16445 52564 0 net90
rlabel metal2 17250 49810 17250 49810 0 net91
rlabel via3 17181 52564 17181 52564 0 net92
rlabel metal2 1610 29886 1610 29886 0 net93
rlabel metal1 2852 35462 2852 35462 0 net94
rlabel metal1 2162 37638 2162 37638 0 net95
rlabel metal1 1748 40358 1748 40358 0 net96
rlabel metal2 8786 17340 8786 17340 0 net97
rlabel metal1 25024 3162 25024 3162 0 net98
rlabel metal1 25484 50694 25484 50694 0 net99
rlabel via2 16790 28373 16790 28373 0 prog_clk
rlabel metal1 23828 2822 23828 2822 0 prog_reset
rlabel metal2 25070 50711 25070 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel via2 25070 51357 25070 51357 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 24932 52462 24932 52462 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 25070 53023 25070 53023 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 24702 52887 24702 52887 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 24794 53635 24794 53635 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 25538 55420 25538 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel metal3 25492 56236 25492 56236 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal1 18170 24854 18170 24854 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 16882 20638 16882 20638 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 16284 21862 16284 21862 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1303 11356 1303 11356 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 18676 14042 18676 14042 0 sb_0__1_.mem_bottom_track_1.ccff_head
rlabel metal1 16100 22066 16100 22066 0 sb_0__1_.mem_bottom_track_1.ccff_tail
rlabel metal1 18170 18938 18170 18938 0 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
rlabel metal2 14582 21692 14582 21692 0 sb_0__1_.mem_bottom_track_1.mem_out\[1\]
rlabel metal1 19458 22542 19458 22542 0 sb_0__1_.mem_bottom_track_11.ccff_head
rlabel metal1 17388 25126 17388 25126 0 sb_0__1_.mem_bottom_track_11.ccff_tail
rlabel metal1 19550 34034 19550 34034 0 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
rlabel metal1 17480 26554 17480 26554 0 sb_0__1_.mem_bottom_track_11.mem_out\[1\]
rlabel metal1 20562 25840 20562 25840 0 sb_0__1_.mem_bottom_track_13.ccff_tail
rlabel metal1 20424 34442 20424 34442 0 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
rlabel metal2 21206 29206 21206 29206 0 sb_0__1_.mem_bottom_track_13.mem_out\[1\]
rlabel metal2 24702 26350 24702 26350 0 sb_0__1_.mem_bottom_track_21.ccff_tail
rlabel metal1 20654 31178 20654 31178 0 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
rlabel metal2 22678 25959 22678 25959 0 sb_0__1_.mem_bottom_track_21.mem_out\[1\]
rlabel metal1 15548 30158 15548 30158 0 sb_0__1_.mem_bottom_track_29.ccff_tail
rlabel metal1 17618 32946 17618 32946 0 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
rlabel metal1 17756 30566 17756 30566 0 sb_0__1_.mem_bottom_track_29.mem_out\[1\]
rlabel metal2 21666 20570 21666 20570 0 sb_0__1_.mem_bottom_track_3.ccff_tail
rlabel metal1 19872 27982 19872 27982 0 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 19780 20842 19780 20842 0 sb_0__1_.mem_bottom_track_3.mem_out\[1\]
rlabel metal1 15456 31450 15456 31450 0 sb_0__1_.mem_bottom_track_37.ccff_tail
rlabel metal1 20378 35530 20378 35530 0 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
rlabel metal1 14720 33286 14720 33286 0 sb_0__1_.mem_bottom_track_37.mem_out\[1\]
rlabel metal1 19872 33626 19872 33626 0 sb_0__1_.mem_bottom_track_45.ccff_tail
rlabel metal1 19872 34986 19872 34986 0 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
rlabel metal1 21528 34034 21528 34034 0 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
rlabel metal1 23966 21454 23966 21454 0 sb_0__1_.mem_bottom_track_5.ccff_tail
rlabel metal1 20654 29104 20654 29104 0 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 24610 23630 24610 23630 0 sb_0__1_.mem_bottom_track_5.mem_out\[1\]
rlabel metal1 15916 37774 15916 37774 0 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
rlabel metal1 19366 31994 19366 31994 0 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
rlabel metal1 19218 22202 19218 22202 0 sb_0__1_.mem_bottom_track_7.mem_out\[1\]
rlabel metal1 17756 38182 17756 38182 0 sb_0__1_.mem_right_track_0.ccff_head
rlabel metal1 23690 29682 23690 29682 0 sb_0__1_.mem_right_track_0.ccff_tail
rlabel metal2 21574 34306 21574 34306 0 sb_0__1_.mem_right_track_0.mem_out\[0\]
rlabel metal1 23046 31858 23046 31858 0 sb_0__1_.mem_right_track_0.mem_out\[1\]
rlabel metal1 23736 44710 23736 44710 0 sb_0__1_.mem_right_track_10.ccff_head
rlabel metal1 21022 41786 21022 41786 0 sb_0__1_.mem_right_track_10.ccff_tail
rlabel metal1 20095 42874 20095 42874 0 sb_0__1_.mem_right_track_10.mem_out\[0\]
rlabel metal1 20286 42126 20286 42126 0 sb_0__1_.mem_right_track_10.mem_out\[1\]
rlabel metal2 20102 44404 20102 44404 0 sb_0__1_.mem_right_track_12.ccff_tail
rlabel metal2 19826 44642 19826 44642 0 sb_0__1_.mem_right_track_12.mem_out\[0\]
rlabel metal1 19320 43214 19320 43214 0 sb_0__1_.mem_right_track_12.mem_out\[1\]
rlabel metal1 18722 44166 18722 44166 0 sb_0__1_.mem_right_track_14.ccff_tail
rlabel metal2 19366 46036 19366 46036 0 sb_0__1_.mem_right_track_14.mem_out\[0\]
rlabel metal1 18906 41650 18906 41650 0 sb_0__1_.mem_right_track_14.mem_out\[1\]
rlabel metal1 17066 44710 17066 44710 0 sb_0__1_.mem_right_track_16.ccff_tail
rlabel metal1 18538 47566 18538 47566 0 sb_0__1_.mem_right_track_16.mem_out\[0\]
rlabel metal1 17480 43214 17480 43214 0 sb_0__1_.mem_right_track_16.mem_out\[1\]
rlabel metal1 15916 40970 15916 40970 0 sb_0__1_.mem_right_track_18.ccff_tail
rlabel metal1 17434 47532 17434 47532 0 sb_0__1_.mem_right_track_18.mem_out\[0\]
rlabel metal2 16146 43452 16146 43452 0 sb_0__1_.mem_right_track_18.mem_out\[1\]
rlabel metal1 25300 43078 25300 43078 0 sb_0__1_.mem_right_track_2.ccff_tail
rlabel metal2 22172 44540 22172 44540 0 sb_0__1_.mem_right_track_2.mem_out\[0\]
rlabel metal1 23460 41650 23460 41650 0 sb_0__1_.mem_right_track_2.mem_out\[1\]
rlabel metal1 14168 34510 14168 34510 0 sb_0__1_.mem_right_track_20.ccff_tail
rlabel metal1 15088 43146 15088 43146 0 sb_0__1_.mem_right_track_20.mem_out\[0\]
rlabel metal2 14030 37706 14030 37706 0 sb_0__1_.mem_right_track_20.mem_out\[1\]
rlabel metal1 12811 29682 12811 29682 0 sb_0__1_.mem_right_track_22.ccff_tail
rlabel metal1 13478 40562 13478 40562 0 sb_0__1_.mem_right_track_22.mem_out\[0\]
rlabel metal1 12880 34170 12880 34170 0 sb_0__1_.mem_right_track_22.mem_out\[1\]
rlabel metal1 14352 26758 14352 26758 0 sb_0__1_.mem_right_track_24.ccff_tail
rlabel metal2 12834 27268 12834 27268 0 sb_0__1_.mem_right_track_24.mem_out\[0\]
rlabel metal2 12926 27200 12926 27200 0 sb_0__1_.mem_right_track_26.ccff_tail
rlabel metal2 14490 27744 14490 27744 0 sb_0__1_.mem_right_track_26.mem_out\[0\]
rlabel metal1 12581 26418 12581 26418 0 sb_0__1_.mem_right_track_28.ccff_tail
rlabel metal2 14858 27438 14858 27438 0 sb_0__1_.mem_right_track_28.mem_out\[0\]
rlabel metal1 9108 28662 9108 28662 0 sb_0__1_.mem_right_track_30.ccff_tail
rlabel metal1 12742 29070 12742 29070 0 sb_0__1_.mem_right_track_30.mem_out\[0\]
rlabel metal1 9016 26826 9016 26826 0 sb_0__1_.mem_right_track_32.ccff_tail
rlabel metal1 7912 27574 7912 27574 0 sb_0__1_.mem_right_track_32.mem_out\[0\]
rlabel metal2 8602 24718 8602 24718 0 sb_0__1_.mem_right_track_34.ccff_tail
rlabel metal1 15502 29138 15502 29138 0 sb_0__1_.mem_right_track_34.mem_out\[0\]
rlabel metal2 8786 12954 8786 12954 0 sb_0__1_.mem_right_track_36.ccff_tail
rlabel metal1 8142 23834 8142 23834 0 sb_0__1_.mem_right_track_36.mem_out\[0\]
rlabel metal2 7866 18666 7866 18666 0 sb_0__1_.mem_right_track_36.mem_out\[1\]
rlabel metal1 13110 11832 13110 11832 0 sb_0__1_.mem_right_track_38.ccff_tail
rlabel metal1 12834 13804 12834 13804 0 sb_0__1_.mem_right_track_38.mem_out\[0\]
rlabel metal2 23414 34816 23414 34816 0 sb_0__1_.mem_right_track_4.ccff_tail
rlabel metal1 24288 42330 24288 42330 0 sb_0__1_.mem_right_track_4.mem_out\[0\]
rlabel metal1 23782 38726 23782 38726 0 sb_0__1_.mem_right_track_4.mem_out\[1\]
rlabel metal1 16146 13498 16146 13498 0 sb_0__1_.mem_right_track_40.ccff_tail
rlabel metal2 14858 14076 14858 14076 0 sb_0__1_.mem_right_track_40.mem_out\[0\]
rlabel metal2 18630 16660 18630 16660 0 sb_0__1_.mem_right_track_44.ccff_tail
rlabel metal1 17112 16150 17112 16150 0 sb_0__1_.mem_right_track_44.mem_out\[0\]
rlabel metal2 20194 17816 20194 17816 0 sb_0__1_.mem_right_track_46.ccff_tail
rlabel metal2 19182 18802 19182 18802 0 sb_0__1_.mem_right_track_46.mem_out\[0\]
rlabel metal1 23230 17850 23230 17850 0 sb_0__1_.mem_right_track_48.ccff_tail
rlabel metal1 21160 17850 21160 17850 0 sb_0__1_.mem_right_track_48.mem_out\[0\]
rlabel metal2 21942 19040 21942 19040 0 sb_0__1_.mem_right_track_50.ccff_tail
rlabel metal1 19918 15980 19918 15980 0 sb_0__1_.mem_right_track_50.mem_out\[0\]
rlabel metal1 21436 12682 21436 12682 0 sb_0__1_.mem_right_track_52.ccff_tail
rlabel metal2 21206 15436 21206 15436 0 sb_0__1_.mem_right_track_52.mem_out\[0\]
rlabel metal2 20010 12070 20010 12070 0 sb_0__1_.mem_right_track_54.ccff_tail
rlabel metal1 19182 13362 19182 13362 0 sb_0__1_.mem_right_track_54.mem_out\[0\]
rlabel metal2 17434 14756 17434 14756 0 sb_0__1_.mem_right_track_56.mem_out\[0\]
rlabel metal1 24932 37774 24932 37774 0 sb_0__1_.mem_right_track_6.ccff_tail
rlabel metal2 22448 40188 22448 40188 0 sb_0__1_.mem_right_track_6.mem_out\[0\]
rlabel metal1 24242 36686 24242 36686 0 sb_0__1_.mem_right_track_6.mem_out\[1\]
rlabel metal1 20102 37774 20102 37774 0 sb_0__1_.mem_right_track_8.mem_out\[0\]
rlabel metal2 22586 44642 22586 44642 0 sb_0__1_.mem_right_track_8.mem_out\[1\]
rlabel metal2 12190 46444 12190 46444 0 sb_0__1_.mem_top_track_0.ccff_tail
rlabel metal2 18170 42942 18170 42942 0 sb_0__1_.mem_top_track_0.mem_out\[0\]
rlabel metal1 12466 44268 12466 44268 0 sb_0__1_.mem_top_track_0.mem_out\[1\]
rlabel metal1 7544 38386 7544 38386 0 sb_0__1_.mem_top_track_10.ccff_head
rlabel metal2 6026 36244 6026 36244 0 sb_0__1_.mem_top_track_10.ccff_tail
rlabel via1 9706 38845 9706 38845 0 sb_0__1_.mem_top_track_10.mem_out\[0\]
rlabel metal1 9476 34034 9476 34034 0 sb_0__1_.mem_top_track_10.mem_out\[1\]
rlabel metal1 7728 32334 7728 32334 0 sb_0__1_.mem_top_track_12.ccff_tail
rlabel metal2 13754 33592 13754 33592 0 sb_0__1_.mem_top_track_12.mem_out\[0\]
rlabel metal1 8234 32946 8234 32946 0 sb_0__1_.mem_top_track_12.mem_out\[1\]
rlabel metal1 13110 44914 13110 44914 0 sb_0__1_.mem_top_track_2.ccff_tail
rlabel metal1 17710 42126 17710 42126 0 sb_0__1_.mem_top_track_2.mem_out\[0\]
rlabel metal1 14582 44302 14582 44302 0 sb_0__1_.mem_top_track_2.mem_out\[1\]
rlabel metal2 9614 35700 9614 35700 0 sb_0__1_.mem_top_track_20.ccff_tail
rlabel metal2 9154 30668 9154 30668 0 sb_0__1_.mem_top_track_20.mem_out\[0\]
rlabel metal1 9929 34374 9929 34374 0 sb_0__1_.mem_top_track_20.mem_out\[1\]
rlabel metal2 5842 38522 5842 38522 0 sb_0__1_.mem_top_track_28.ccff_tail
rlabel metal2 13478 34612 13478 34612 0 sb_0__1_.mem_top_track_28.mem_out\[0\]
rlabel metal1 7636 35258 7636 35258 0 sb_0__1_.mem_top_track_28.mem_out\[1\]
rlabel metal1 10258 42092 10258 42092 0 sb_0__1_.mem_top_track_36.ccff_tail
rlabel metal1 7130 40562 7130 40562 0 sb_0__1_.mem_top_track_36.mem_out\[0\]
rlabel metal1 12466 38352 12466 38352 0 sb_0__1_.mem_top_track_36.mem_out\[1\]
rlabel metal1 10534 40902 10534 40902 0 sb_0__1_.mem_top_track_4.ccff_tail
rlabel metal1 14076 43078 14076 43078 0 sb_0__1_.mem_top_track_4.mem_out\[0\]
rlabel metal1 14858 38420 14858 38420 0 sb_0__1_.mem_top_track_4.mem_out\[1\]
rlabel metal1 12558 42568 12558 42568 0 sb_0__1_.mem_top_track_44.ccff_tail
rlabel metal2 13754 39440 13754 39440 0 sb_0__1_.mem_top_track_44.mem_out\[0\]
rlabel metal1 16652 42534 16652 42534 0 sb_0__1_.mem_top_track_52.mem_out\[0\]
rlabel metal1 15962 38250 15962 38250 0 sb_0__1_.mem_top_track_52.mem_out\[1\]
rlabel metal1 18538 37978 18538 37978 0 sb_0__1_.mem_top_track_6.mem_out\[0\]
rlabel metal2 8602 37944 8602 37944 0 sb_0__1_.mem_top_track_6.mem_out\[1\]
rlabel metal1 14950 14586 14950 14586 0 sb_0__1_.mux_bottom_track_1.out
rlabel metal1 15732 26010 15732 26010 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18216 32198 18216 32198 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14030 22066 14030 22066 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15180 22746 15180 22746 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13708 21658 13708 21658 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15180 22406 15180 22406 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 16882 14693 16882 14693 0 sb_0__1_.mux_bottom_track_11.out
rlabel metal1 17434 28594 17434 28594 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18676 34102 18676 34102 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16882 25024 16882 25024 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14214 24650 14214 24650 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16928 24242 16928 24242 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 16790 24820 16790 24820 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 17112 17170 17112 17170 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 18814 19686 18814 19686 0 sb_0__1_.mux_bottom_track_13.out
rlabel metal1 20102 29716 20102 29716 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20792 34714 20792 34714 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18814 27098 18814 27098 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20378 27744 20378 27744 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19918 26010 19918 26010 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18814 19822 18814 19822 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 21022 8534 21022 8534 0 sb_0__1_.mux_bottom_track_21.out
rlabel metal1 21758 29478 21758 29478 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21988 29614 21988 29614 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21114 27336 21114 27336 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 25392 24174 25392 24174 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 24978 24786 24978 24786 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23506 14994 23506 14994 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 14536 17578 14536 17578 0 sb_0__1_.mux_bottom_track_29.out
rlabel metal1 17342 32300 17342 32300 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17250 34510 17250 34510 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17434 29274 17434 29274 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16790 32198 16790 32198 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16468 28526 16468 28526 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15732 28390 15732 28390 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 19734 14790 19734 14790 0 sb_0__1_.mux_bottom_track_3.out
rlabel metal1 19504 25330 19504 25330 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19642 25262 19642 25262 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19504 20570 19504 20570 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19366 20808 19366 20808 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19826 17612 19826 17612 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13248 21862 13248 21862 0 sb_0__1_.mux_bottom_track_37.out
rlabel metal1 16330 34646 16330 34646 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17894 34714 17894 34714 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14904 29274 14904 29274 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13478 28730 13478 28730 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13478 21998 13478 21998 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 18768 15028 18768 15028 0 sb_0__1_.mux_bottom_track_45.out
rlabel metal1 20838 36210 20838 36210 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20424 31790 20424 31790 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20930 33830 20930 33830 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal3 19067 20604 19067 20604 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20608 10540 20608 10540 0 sb_0__1_.mux_bottom_track_5.out
rlabel metal1 21114 29036 21114 29036 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21896 26554 21896 26554 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24840 23154 24840 23154 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22724 26486 22724 26486 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22908 21522 22908 21522 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 21298 18394 21298 18394 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9798 16422 9798 16422 0 sb_0__1_.mux_bottom_track_53.out
rlabel metal1 13662 38760 13662 38760 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13202 37196 13202 37196 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10902 27030 10902 27030 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19136 19210 19136 19210 0 sb_0__1_.mux_bottom_track_7.out
rlabel metal1 18906 26418 18906 26418 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20470 31926 20470 31926 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18308 24582 18308 24582 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17664 21930 17664 21930 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19734 24582 19734 24582 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18722 21998 18722 21998 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 19044 19414 19044 19414 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 22632 26962 22632 26962 0 sb_0__1_.mux_right_track_0.out
rlabel metal1 21988 31858 21988 31858 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22126 32742 22126 32742 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22678 31926 22678 31926 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23322 29240 23322 29240 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 24794 29138 24794 29138 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23460 31994 23460 31994 0 sb_0__1_.mux_right_track_10.out
rlabel metal1 20838 45798 20838 45798 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19688 39882 19688 39882 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20700 42262 20700 42262 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17480 36346 17480 36346 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22034 32436 22034 32436 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 22816 32198 22816 32198 0 sb_0__1_.mux_right_track_12.out
rlabel metal1 19826 45798 19826 45798 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19688 39474 19688 39474 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17066 38114 17066 38114 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19688 39270 19688 39270 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23966 25262 23966 25262 0 sb_0__1_.mux_right_track_14.out
rlabel metal1 18584 41650 18584 41650 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18308 41446 18308 41446 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17434 37638 17434 37638 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal4 19228 36584 19228 36584 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22356 25942 22356 25942 0 sb_0__1_.mux_right_track_16.out
rlabel metal1 17802 47430 17802 47430 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17112 40562 17112 40562 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15134 39542 15134 39542 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20286 32368 20286 32368 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21896 24174 21896 24174 0 sb_0__1_.mux_right_track_18.out
rlabel metal1 16652 41582 16652 41582 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16422 37298 16422 37298 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15318 37230 15318 37230 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16284 37094 16284 37094 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24656 29206 24656 29206 0 sb_0__1_.mux_right_track_2.out
rlabel metal1 23046 41650 23046 41650 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22770 41514 22770 41514 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20240 37638 20240 37638 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23966 41718 23966 41718 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24472 39338 24472 39338 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 24794 36618 24794 36618 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 19872 27574 19872 27574 0 sb_0__1_.mux_right_track_20.out
rlabel metal1 14444 43078 14444 43078 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14536 32946 14536 32946 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14674 32640 14674 32640 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18032 27438 18032 27438 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19734 19890 19734 19890 0 sb_0__1_.mux_right_track_22.out
rlabel metal1 13064 34034 13064 34034 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12926 33830 12926 33830 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 10442 29818 10442 29818 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17802 24140 17802 24140 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21482 20808 21482 20808 0 sb_0__1_.mux_right_track_24.out
rlabel metal1 15180 24786 15180 24786 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13938 24922 13938 24922 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17526 20978 17526 20978 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21298 18224 21298 18224 0 sb_0__1_.mux_right_track_26.out
rlabel metal1 15180 27098 15180 27098 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14214 26214 14214 26214 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16744 21658 16744 21658 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21206 21080 21206 21080 0 sb_0__1_.mux_right_track_28.out
rlabel metal1 13478 26350 13478 26350 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9246 26282 9246 26282 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17066 21556 17066 21556 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21298 17068 21298 17068 0 sb_0__1_.mux_right_track_30.out
rlabel metal2 10902 27506 10902 27506 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10672 26010 10672 26010 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16238 21284 16238 21284 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20930 16082 20930 16082 0 sb_0__1_.mux_right_track_32.out
rlabel metal1 10672 25262 10672 25262 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8050 24650 8050 24650 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14582 20434 14582 20434 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21850 15538 21850 15538 0 sb_0__1_.mux_right_track_34.out
rlabel metal2 13570 26622 13570 26622 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11178 24378 11178 24378 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15962 19346 15962 19346 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17756 10506 17756 10506 0 sb_0__1_.mux_right_track_36.out
rlabel metal1 7682 18394 7682 18394 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8234 12954 8234 12954 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7590 12818 7590 12818 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 14858 11696 14858 11696 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22218 10064 22218 10064 0 sb_0__1_.mux_right_track_38.out
rlabel metal1 15318 11866 15318 11866 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18400 10642 18400 10642 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 25162 28798 25162 28798 0 sb_0__1_.mux_right_track_4.out
rlabel metal1 21988 43622 21988 43622 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22816 38250 22816 38250 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21942 36108 21942 36108 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22494 33456 22494 33456 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23092 34102 23092 34102 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23414 10676 23414 10676 0 sb_0__1_.mux_right_track_40.out
rlabel metal2 17342 14042 17342 14042 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20194 12614 20194 12614 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23736 9962 23736 9962 0 sb_0__1_.mux_right_track_44.out
rlabel metal2 18906 16354 18906 16354 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18676 14790 18676 14790 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24886 10642 24886 10642 0 sb_0__1_.mux_right_track_46.out
rlabel metal1 20562 16626 20562 16626 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 12172 22862 12172 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24932 6766 24932 6766 0 sb_0__1_.mux_right_track_48.out
rlabel metal2 20838 17748 20838 17748 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23506 12240 23506 12240 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23322 8942 23322 8942 0 sb_0__1_.mux_right_track_50.out
rlabel metal1 21298 19482 21298 19482 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20194 16218 20194 16218 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20746 19448 20746 19448 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23414 4590 23414 4590 0 sb_0__1_.mux_right_track_52.out
rlabel metal1 20516 15402 20516 15402 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21114 10812 21114 10812 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24058 4522 24058 4522 0 sb_0__1_.mux_right_track_54.out
rlabel metal1 18584 13430 18584 13430 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21206 8942 21206 8942 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24702 5576 24702 5576 0 sb_0__1_.mux_right_track_56.out
rlabel metal2 19918 14416 19918 14416 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21206 13226 21206 13226 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24564 26350 24564 26350 0 sb_0__1_.mux_right_track_6.out
rlabel metal1 23506 43078 23506 43078 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24702 38080 24702 38080 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20930 33320 20930 33320 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23782 37196 23782 37196 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23460 34714 23460 34714 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23874 36278 23874 36278 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24564 34714 24564 34714 0 sb_0__1_.mux_right_track_8.out
rlabel metal1 22172 42738 22172 42738 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21712 42602 21712 42602 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21850 41514 21850 41514 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21988 42534 21988 42534 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 21666 40970 21666 40970 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23966 34578 23966 34578 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12282 51986 12282 51986 0 sb_0__1_.mux_top_track_0.out
rlabel metal1 10442 43146 10442 43146 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17158 42568 17158 42568 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14950 39168 14950 39168 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10304 37978 10304 37978 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11546 44506 11546 44506 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 11730 41321 11730 41321 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 10718 47668 10718 47668 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7958 44506 7958 44506 0 sb_0__1_.mux_top_track_10.out
rlabel metal1 9430 38386 9430 38386 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13110 36992 13110 36992 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12742 30906 12742 30906 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8602 33898 8602 33898 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8234 36890 8234 36890 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8510 34170 8510 34170 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7866 44370 7866 44370 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 7774 46614 7774 46614 0 sb_0__1_.mux_top_track_12.out
rlabel metal2 10902 35088 10902 35088 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11914 32742 11914 32742 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7866 32810 7866 32810 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 10442 34850 10442 34850 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 7498 34544 7498 34544 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7820 43282 7820 43282 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12788 48858 12788 48858 0 sb_0__1_.mux_top_track_2.out
rlabel metal1 16376 42330 16376 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16836 42262 16836 42262 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13432 42058 13432 42058 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15318 42330 15318 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13248 42330 13248 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12788 45050 12788 45050 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8924 43962 8924 43962 0 sb_0__1_.mux_top_track_20.out
rlabel metal1 14030 35054 14030 35054 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15364 34578 15364 34578 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9706 32742 9706 32742 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 9430 35938 9430 35938 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9384 33082 9384 33082 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8786 40902 8786 40902 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 5842 47396 5842 47396 0 sb_0__1_.mux_top_track_28.out
rlabel metal1 10994 36142 10994 36142 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11362 34816 11362 34816 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9154 37162 9154 37162 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 5014 35190 5014 35190 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 5658 44370 5658 44370 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7360 46682 7360 46682 0 sb_0__1_.mux_top_track_36.out
rlabel metal1 12282 38386 12282 38386 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11040 38454 11040 38454 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7820 38522 7820 38522 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 9706 42466 9706 42466 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11408 51986 11408 51986 0 sb_0__1_.mux_top_track_4.out
rlabel metal1 14996 38318 14996 38318 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19366 36346 19366 36346 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11132 33082 11132 33082 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13340 38522 13340 38522 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10764 38522 10764 38522 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10902 41786 10902 41786 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8050 52054 8050 52054 0 sb_0__1_.mux_top_track_44.out
rlabel metal2 15594 41208 15594 41208 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10810 38794 10810 38794 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11638 42330 11638 42330 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8878 46070 8878 46070 0 sb_0__1_.mux_top_track_52.out
rlabel metal1 20240 38998 20240 38998 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17618 39066 17618 39066 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14858 36346 14858 36346 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14168 45866 14168 45866 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9844 51374 9844 51374 0 sb_0__1_.mux_top_track_6.out
rlabel metal1 9752 39474 9752 39474 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17710 38454 17710 38454 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14260 31926 14260 31926 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9200 34986 9200 34986 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9154 39610 9154 39610 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9062 35258 9062 35258 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7268 40154 7268 40154 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 1380 45594 1380 45594 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 1518 48042 1518 48042 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 1334 50439 1334 50439 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 4002 52564 4002 52564 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
